C0000737|ICD9CM|HT|789.0|Abdominal pain
C0000737|ICD9CM|PT|789.00|Abdominal pain, unspecified site
C0000768|ICD9CM|HT|740-759.99|CONGENITAL ANOMALIES
C0000768|ICD9CM|PT|759.9|Congenital anomaly, unspecified
C0000770|ICD9CM|PT|520.2|Abnormalities of size and form of teeth
C0000774|ICD9CM|PT|251.5|Abnormality of secretion of gastrin
C0000786|ICD9CM|HT|634|Spontaneous abortion
C0000804|ICD9CM|HT|636|Illegally induced abortion
C0000814|ICD9CM|PT|632|Missed abortion
C0000821|ICD9CM|HT|640.0|Threatened abortion

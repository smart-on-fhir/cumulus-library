C0000727|ICD10CM|PT|R10.0|Acute abdomen
C0000737|ICD10CM|PT|R10.9|Unspecified abdominal pain
C0000744|ICD10CM|ET|E78.6|Abetalipoproteinemia
C0000768|ICD10CM|ET|Q89.9|Congenital anomaly NOS
C0000768|ICD10CM|PT|Q89.9|Congenital malformation, unspecified
C0000768|ICD10CM|ET|Q89.9|Congenital deformity NOS
C0000770|ICD10CM|PT|K00.2|Abnormalities of size and form of teeth
C0000772|ICD10CM|ET|Q89.7|Multiple congenital anomalies NOS
C0000772|ICD10CM|ET|Q89.7|Multiple congenital deformities NOS
C0000786|ICD10CM|HT|O03|Spontaneous abortion

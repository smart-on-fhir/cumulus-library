C0000727|ICD10CM|PT|R10.0|Acute abdomen
C0000737|ICD10CM|PT|R10.9|Unspecified abdominal pain
C0000744|ICD10CM|ET|E78.6|Abetalipoproteinemia

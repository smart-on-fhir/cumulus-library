C0005491|ICD10PCS|PT|GZC9ZZZ|Biofeedback
C0005491|ICD10PCS|PX|GZC9ZZZ|Mental Health @ None @ Biofeedback @ Other Biofeedback @ None @ None @ None
C0010332|ICD10PCS|PT|GZ2ZZZZ|Crisis Intervention
C0010332|ICD10PCS|PX|GZ2ZZZZ|Mental Health @ None @ Crisis Intervention @ None @ None @ None @ None
C0011931|ICD10PCS|PT|BH4CZZZ|Ultrasonography of Head and Neck
C0011931|ICD10PCS|PX|BH4CZZZ|Imaging @ Skin, Subcutaneous Tissue and Breast @ Ultrasonography @ Head and Neck @ None @ None @ None
C0015400|ICD10PCS|HT|08P|Eye, Removal
C0015400|ICD10PCS|HX|08P|Medical and Surgical @ Eye @ Removal
C0015618|ICD10PCS|PT|GZ72ZZZ|Family Psychotherapy
C0015618|ICD10PCS|PX|GZ72ZZZ|Mental Health @ None @ Family Psychotherapy @ Other Family Psychotherapy @ None @ None @ None

C0005491|ICD10PCS|PT|GZC9ZZZ|Biofeedback
C0005491|ICD10PCS|PX|GZC9ZZZ|Mental Health @ None @ Biofeedback @ Other Biofeedback @ None @ None @ None
C0010332|ICD10PCS|PT|GZ2ZZZZ|Crisis Intervention

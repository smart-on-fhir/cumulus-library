C0008354|T047|HT|001|ICD9CM|Cholera|Cholera
C0178238|T047|HT|001-009.99|ICD9CM|INTESTINAL INFECTIOUS DISEASES|INTESTINAL INFECTIOUS DISEASES
C0041849|T047|HT|001-139.99|ICD9CM|INFECTIOUS AND PARASITIC DISEASES|INFECTIOUS AND PARASITIC DISEASES
C0178237|T047|HT|001-999.99|ICD9CM|DISEASES AND INJURIES|DISEASES AND INJURIES
C0008354|T047|AB|001.0|ICD9CM|Cholera d/t vib cholerae|Cholera d/t vib cholerae
C0008354|T047|PT|001.0|ICD9CM|Cholera due to vibrio cholerae|Cholera due to vibrio cholerae
C0343372|T047|AB|001.1|ICD9CM|Cholera d/t vib el tor|Cholera d/t vib el tor
C0343372|T047|PT|001.1|ICD9CM|Cholera due to vibrio cholerae el tor|Cholera due to vibrio cholerae el tor
C0008354|T047|AB|001.9|ICD9CM|Cholera NOS|Cholera NOS
C0008354|T047|PT|001.9|ICD9CM|Cholera, unspecified|Cholera, unspecified
C0275976|T047|HT|002|ICD9CM|Typhoid and paratyphoid fevers|Typhoid and paratyphoid fevers
C0041466|T047|AB|002.0|ICD9CM|Typhoid fever|Typhoid fever
C0041466|T047|PT|002.0|ICD9CM|Typhoid fever|Typhoid fever
C0343375|T047|AB|002.1|ICD9CM|Paratyphoid fever a|Paratyphoid fever a
C0343375|T047|PT|002.1|ICD9CM|Paratyphoid fever A|Paratyphoid fever A
C0343376|T047|AB|002.2|ICD9CM|Paratyphoid fever b|Paratyphoid fever b
C0343376|T047|PT|002.2|ICD9CM|Paratyphoid fever B|Paratyphoid fever B
C0343377|T047|AB|002.3|ICD9CM|Paratyphoid fever c|Paratyphoid fever c
C0343377|T047|PT|002.3|ICD9CM|Paratyphoid fever C|Paratyphoid fever C
C0030528|T047|AB|002.9|ICD9CM|Paratyphoid fever NOS|Paratyphoid fever NOS
C0030528|T047|PT|002.9|ICD9CM|Paratyphoid fever, unspecified|Paratyphoid fever, unspecified
C0152485|T047|HT|003|ICD9CM|Other salmonella infections|Other salmonella infections
C0036114|T037|AB|003.0|ICD9CM|Salmonella enteritis|Salmonella enteritis
C0036114|T037|PT|003.0|ICD9CM|Salmonella gastroenteritis|Salmonella gastroenteritis
C0152486|T047|AB|003.1|ICD9CM|Salmonella septicemia|Salmonella septicemia
C0152486|T047|PT|003.1|ICD9CM|Salmonella septicemia|Salmonella septicemia
C0152487|T047|HT|003.2|ICD9CM|Localized salmonella infections|Localized salmonella infections
C0152487|T047|AB|003.20|ICD9CM|Local salmonella inf NOS|Local salmonella inf NOS
C0152487|T047|PT|003.20|ICD9CM|Localized salmonella infection, unspecified|Localized salmonella infection, unspecified
C0152488|T047|AB|003.21|ICD9CM|Salmonella meningitis|Salmonella meningitis
C0152488|T047|PT|003.21|ICD9CM|Salmonella meningitis|Salmonella meningitis
C0152489|T047|AB|003.22|ICD9CM|Salmonella pneumonia|Salmonella pneumonia
C0152489|T047|PT|003.22|ICD9CM|Salmonella pneumonia|Salmonella pneumonia
C0152490|T047|AB|003.23|ICD9CM|Salmonella arthritis|Salmonella arthritis
C0152490|T047|PT|003.23|ICD9CM|Salmonella arthritis|Salmonella arthritis
C0152491|T047|AB|003.24|ICD9CM|Salmonella osteomyelitis|Salmonella osteomyelitis
C0152491|T047|PT|003.24|ICD9CM|Salmonella osteomyelitis|Salmonella osteomyelitis
C0152492|T047|AB|003.29|ICD9CM|Local salmonella inf NEC|Local salmonella inf NEC
C0152492|T047|PT|003.29|ICD9CM|Other localized salmonella infections|Other localized salmonella infections
C0029826|T047|PT|003.8|ICD9CM|Other specified salmonella infections|Other specified salmonella infections
C0029826|T047|AB|003.8|ICD9CM|Salmonella infection NEC|Salmonella infection NEC
C0036117|T047|AB|003.9|ICD9CM|Salmonella infection NOS|Salmonella infection NOS
C0036117|T047|PT|003.9|ICD9CM|Salmonella infection, unspecified|Salmonella infection, unspecified
C0013371|T047|HT|004|ICD9CM|Shigellosis|Shigellosis
C0302358|T047|AB|004.0|ICD9CM|Shigella dysenteriae|Shigella dysenteriae
C0302358|T047|PT|004.0|ICD9CM|Shigella dysenteriae|Shigella dysenteriae
C0302359|T047|AB|004.1|ICD9CM|Shigella flexneri|Shigella flexneri
C0302359|T047|PT|004.1|ICD9CM|Shigella flexneri|Shigella flexneri
C0302360|T047|AB|004.2|ICD9CM|Shigella boydii|Shigella boydii
C0302360|T047|PT|004.2|ICD9CM|Shigella boydii|Shigella boydii
C0302361|T047|AB|004.3|ICD9CM|Shigella sonnei|Shigella sonnei
C0302361|T047|PT|004.3|ICD9CM|Shigella sonnei|Shigella sonnei
C0152493|T047|PT|004.8|ICD9CM|Other specified shigella infections|Other specified shigella infections
C0152493|T047|AB|004.8|ICD9CM|Shigella infection NEC|Shigella infection NEC
C0013371|T047|AB|004.9|ICD9CM|Shigellosis NOS|Shigellosis NOS
C0013371|T047|PT|004.9|ICD9CM|Shigellosis, unspecified|Shigellosis, unspecified
C0152498|T037|HT|005|ICD9CM|Other food poisoning (bacterial)|Other food poisoning (bacterial)
C0038159|T047|AB|005.0|ICD9CM|Staph food poisoning|Staph food poisoning
C0038159|T047|PT|005.0|ICD9CM|Staphylococcal food poisoning|Staphylococcal food poisoning
C1739094|T047|PT|005.1|ICD9CM|Botulism food poisoning|Botulism food poisoning
C1739094|T047|AB|005.1|ICD9CM|Botulism food poisoning|Botulism food poisoning
C0275590|T037|AB|005.2|ICD9CM|Food pois d/t c. perfrin|Food pois d/t c. perfrin
C0275590|T037|PT|005.2|ICD9CM|Food poisoning due to Clostridium perfringens (C. welchii)|Food poisoning due to Clostridium perfringens (C. welchii)
C0152496|T037|AB|005.3|ICD9CM|Food pois: clostrid NEC|Food pois: clostrid NEC
C0152496|T037|PT|005.3|ICD9CM|Food poisoning due to other Clostridia|Food poisoning due to other Clostridia
C0152497|T047|AB|005.4|ICD9CM|Food pois: v. parahaem|Food pois: v. parahaem
C0152497|T047|PT|005.4|ICD9CM|Food poisoning due to Vibrio parahaemolyticus|Food poisoning due to Vibrio parahaemolyticus
C0152498|T037|HT|005.8|ICD9CM|Other bacterial food poisoning|Other bacterial food poisoning
C0374921|T037|AB|005.81|ICD9CM|Food poisn d/t v. vulnif|Food poisn d/t v. vulnif
C0374921|T037|PT|005.81|ICD9CM|Food poisoning due to Vibrio vulnificus|Food poisoning due to Vibrio vulnificus
C0152498|T037|AB|005.89|ICD9CM|Bact food poisoning NEC|Bact food poisoning NEC
C0152498|T037|PT|005.89|ICD9CM|Other bacterial food poisoning|Other bacterial food poisoning
C0016479|T037|AB|005.9|ICD9CM|Food poisoning NOS|Food poisoning NOS
C0016479|T037|PT|005.9|ICD9CM|Food poisoning, unspecified|Food poisoning, unspecified
C0002438|T047|HT|006|ICD9CM|Amebiasis|Amebiasis
C1363999|T047|AB|006.0|ICD9CM|Ac amebiasis w/o abscess|Ac amebiasis w/o abscess
C1363999|T047|PT|006.0|ICD9CM|Acute amebic dysentery without mention of abscess|Acute amebic dysentery without mention of abscess
C0152500|T047|AB|006.1|ICD9CM|Chr amebiasis w/o absces|Chr amebiasis w/o absces
C0152500|T047|PT|006.1|ICD9CM|Chronic intestinal amebiasis without mention of abscess|Chronic intestinal amebiasis without mention of abscess
C0152501|T047|AB|006.2|ICD9CM|Amebic nondysent colitis|Amebic nondysent colitis
C0152501|T047|PT|006.2|ICD9CM|Amebic nondysenteric colitis|Amebic nondysenteric colitis
C0023886|T047|AB|006.3|ICD9CM|Amebic liver abscess|Amebic liver abscess
C0023886|T047|PT|006.3|ICD9CM|Amebic liver abscess|Amebic liver abscess
C0152502|T047|AB|006.4|ICD9CM|Amebic lung abscess|Amebic lung abscess
C0152502|T047|PT|006.4|ICD9CM|Amebic lung abscess|Amebic lung abscess
C0152503|T047|AB|006.5|ICD9CM|Amebic brain abscess|Amebic brain abscess
C0152503|T047|PT|006.5|ICD9CM|Amebic brain abscess|Amebic brain abscess
C1318565|T047|AB|006.6|ICD9CM|Amebic skin ulceration|Amebic skin ulceration
C1318565|T047|PT|006.6|ICD9CM|Amebic skin ulceration|Amebic skin ulceration
C0152505|T047|AB|006.8|ICD9CM|Amebic infection NEC|Amebic infection NEC
C0152505|T047|PT|006.8|ICD9CM|Amebic infection of other sites|Amebic infection of other sites
C0002438|T047|AB|006.9|ICD9CM|Amebiasis NOS|Amebiasis NOS
C0002438|T047|PT|006.9|ICD9CM|Amebiasis, unspecified|Amebiasis, unspecified
C0152506|T047|HT|007|ICD9CM|Other protozoal intestinal diseases|Other protozoal intestinal diseases
C0004692|T047|AB|007.0|ICD9CM|Balantidiasis|Balantidiasis
C0004692|T047|PT|007.0|ICD9CM|Balantidiasis|Balantidiasis
C0017536|T047|AB|007.1|ICD9CM|Giardiasis|Giardiasis
C0017536|T047|PT|007.1|ICD9CM|Giardiasis|Giardiasis
C1299919|T047|AB|007.2|ICD9CM|Coccidiosis|Coccidiosis
C1299919|T047|PT|007.2|ICD9CM|Coccidiosis|Coccidiosis
C0411268|T047|AB|007.3|ICD9CM|Intest trichomoniasis|Intest trichomoniasis
C0411268|T047|PT|007.3|ICD9CM|Intestinal trichomoniasis|Intestinal trichomoniasis
C0010418|T047|AB|007.4|ICD9CM|Cryptosporidiosis|Cryptosporidiosis
C0010418|T047|PT|007.4|ICD9CM|Cryptosporidiosis|Cryptosporidiosis
C0343398|T047|AB|007.5|ICD9CM|Cyclosporiasis|Cyclosporiasis
C0343398|T047|PT|007.5|ICD9CM|Cyclosporiasis|Cyclosporiasis
C0152507|T047|PT|007.8|ICD9CM|Other specified protozoal intestinal diseases|Other specified protozoal intestinal diseases
C0152507|T047|AB|007.8|ICD9CM|Protozoal intest dis NEC|Protozoal intest dis NEC
C0276774|T047|AB|007.9|ICD9CM|Protozoal intest dis NOS|Protozoal intest dis NOS
C0276774|T047|PT|007.9|ICD9CM|Unspecified protozoal intestinal disease|Unspecified protozoal intestinal disease
C0152518|T047|HT|008|ICD9CM|Intestinal infections due to other organisms|Intestinal infections due to other organisms
C0341558|T047|HT|008.0|ICD9CM|Intestinal infection due to escherichia coli [E. coli]|Intestinal infection due to escherichia coli [E. coli]
C0341558|T047|AB|008.00|ICD9CM|Intest infec e coli NOS|Intest infec e coli NOS
C0341558|T047|PT|008.00|ICD9CM|Intestinal infection due to E. coli, unspecified|Intestinal infection due to E. coli, unspecified
C0343380|T047|AB|008.01|ICD9CM|Int inf e coli entrpath|Int inf e coli entrpath
C0343380|T047|PT|008.01|ICD9CM|Intestinal infection due to enteropathogenic E. coli|Intestinal infection due to enteropathogenic E. coli
C0343379|T047|AB|008.02|ICD9CM|Int inf e coli entrtoxgn|Int inf e coli entrtoxgn
C0343379|T047|PT|008.02|ICD9CM|Intestinal infection due to enterotoxigenic E. coli|Intestinal infection due to enterotoxigenic E. coli
C0343382|T047|AB|008.03|ICD9CM|Int inf e coli entrnvsv|Int inf e coli entrnvsv
C0343382|T047|PT|008.03|ICD9CM|Intestinal infection due to enteroinvasive E. coli|Intestinal infection due to enteroinvasive E. coli
C0343381|T047|AB|008.04|ICD9CM|Int inf e coli entrhmrg|Int inf e coli entrhmrg
C0343381|T047|PT|008.04|ICD9CM|Intestinal infection due to enterohemorrhagic E. coli|Intestinal infection due to enterohemorrhagic E. coli
C0494024|T047|AB|008.09|ICD9CM|Int inf e coli spcf NEC|Int inf e coli spcf NEC
C0494024|T047|PT|008.09|ICD9CM|Intestinal infection due to other intestinal E. coli infections|Intestinal infection due to other intestinal E. coli infections
C0152511|T047|AB|008.1|ICD9CM|Arizona enteritis|Arizona enteritis
C0152511|T047|PT|008.1|ICD9CM|Intestinal infection due to arizona group of paracolon bacilli|Intestinal infection due to arizona group of paracolon bacilli
C0276058|T047|AB|008.2|ICD9CM|Aerobacter enteritis|Aerobacter enteritis
C0276058|T047|PT|008.2|ICD9CM|Intestinal infection due to aerobacter aerogenes|Intestinal infection due to aerobacter aerogenes
C0152513|T047|PT|008.3|ICD9CM|Intestinal infection due to proteus (mirabilis) (morganii)|Intestinal infection due to proteus (mirabilis) (morganii)
C0152513|T047|AB|008.3|ICD9CM|Proteus enteritis|Proteus enteritis
C0489951|T047|HT|008.4|ICD9CM|Intestinal infection due to other specified bacteria|Intestinal infection due to other specified bacteria
C0038157|T047|PT|008.41|ICD9CM|Intestinal infection due to staphylococcus|Intestinal infection due to staphylococcus
C0038157|T047|AB|008.41|ICD9CM|Staphylococc enteritis|Staphylococc enteritis
C0152515|T047|PT|008.42|ICD9CM|Intestinal infection due to pseudomonas|Intestinal infection due to pseudomonas
C0152515|T047|AB|008.42|ICD9CM|Pseudomonas enteritis|Pseudomonas enteritis
C0275982|T047|AB|008.43|ICD9CM|Int infec campylobacter|Int infec campylobacter
C0275982|T047|PT|008.43|ICD9CM|Intestinal infection due to campylobacter|Intestinal infection due to campylobacter
C0238528|T047|AB|008.44|ICD9CM|Int inf yrsnia entrcltca|Int inf yrsnia entrcltca
C0238528|T047|PT|008.44|ICD9CM|Intestinal infection due to yersinia enterocolitica|Intestinal infection due to yersinia enterocolitica
C0494025|T047|AB|008.45|ICD9CM|Int inf clstrdium dfcile|Int inf clstrdium dfcile
C0494025|T047|PT|008.45|ICD9CM|Intestinal infection due to Clostridium difficile|Intestinal infection due to Clostridium difficile
C0374931|T047|AB|008.46|ICD9CM|Intes infec oth anerobes|Intes infec oth anerobes
C0374931|T047|PT|008.46|ICD9CM|Intestinal infection due to other anaerobes|Intestinal infection due to other anaerobes
C0374932|T047|AB|008.47|ICD9CM|Int inf oth grm neg bctr|Int inf oth grm neg bctr
C0374932|T047|PT|008.47|ICD9CM|Intestinal infection due to other gram-negative bacteria|Intestinal infection due to other gram-negative bacteria
C0489951|T047|AB|008.49|ICD9CM|Bacterial enteritis NEC|Bacterial enteritis NEC
C0489951|T047|PT|008.49|ICD9CM|Intestinal infection due to other organisms|Intestinal infection due to other organisms
C0152516|T047|AB|008.5|ICD9CM|Bacterial enteritis NOS|Bacterial enteritis NOS
C0152516|T047|PT|008.5|ICD9CM|Bacterial enteritis, unspecified|Bacterial enteritis, unspecified
C0152517|T047|HT|008.6|ICD9CM|Enteritis due to specified virus|Enteritis due to specified virus
C0347854|T047|PT|008.61|ICD9CM|Enteritis due to rotavirus|Enteritis due to rotavirus
C0347854|T047|AB|008.61|ICD9CM|Intes infec rotavirus|Intes infec rotavirus
C0276162|T047|PT|008.62|ICD9CM|Enteritis due to adenovirus|Enteritis due to adenovirus
C0276162|T047|AB|008.62|ICD9CM|Intes infec adenovirus|Intes infec adenovirus
C0374933|T047|PT|008.63|ICD9CM|Enteritis due to norwalk virus|Enteritis due to norwalk virus
C0374933|T047|AB|008.63|ICD9CM|Int inf norwalk virus|Int inf norwalk virus
C0374934|T047|PT|008.64|ICD9CM|Enteritis due to other small round viruses [SRV's]|Enteritis due to other small round viruses [SRV's]
C0374934|T047|AB|008.64|ICD9CM|Int inf oth sml rnd vrus|Int inf oth sml rnd vrus
C1611187|T047|AB|008.65|ICD9CM|Enteritis d/t calicivirs|Enteritis d/t calicivirs
C1611187|T047|PT|008.65|ICD9CM|Enteritis due to calicivirus|Enteritis due to calicivirus
C0374936|T047|PT|008.66|ICD9CM|Enteritis due to astrovirus|Enteritis due to astrovirus
C0374936|T047|AB|008.66|ICD9CM|Intes infec astrovirus|Intes infec astrovirus
C0374937|T047|PT|008.67|ICD9CM|Enteritis due to enterovirus nec|Enteritis due to enterovirus nec
C0374937|T047|AB|008.67|ICD9CM|Int inf enterovirus NEC|Int inf enterovirus NEC
C0348098|T047|PT|008.69|ICD9CM|Enteritis due to other viral enteritis|Enteritis due to other viral enteritis
C0348098|T047|AB|008.69|ICD9CM|Other viral intes infec|Other viral intes infec
C0489952|T047|PT|008.8|ICD9CM|Intestinal infection due to other organism, not elsewhere classified|Intestinal infection due to other organism, not elsewhere classified
C0489952|T047|AB|008.8|ICD9CM|Viral enteritis NOS|Viral enteritis NOS
C0152519|T047|HT|009|ICD9CM|Ill-defined intestinal infections|Ill-defined intestinal infections
C1279224|T047|PT|009.0|ICD9CM|Infectious colitis, enteritis, and gastroenteritis|Infectious colitis, enteritis, and gastroenteritis
C1279224|T047|AB|009.0|ICD9CM|Infectious enteritis NOS|Infectious enteritis NOS
C0595979|T047|PT|009.1|ICD9CM|Colitis, enteritis, and gastroenteritis of presumed infectious origin|Colitis, enteritis, and gastroenteritis of presumed infectious origin
C0595979|T047|AB|009.1|ICD9CM|Enteritis of infect orig|Enteritis of infect orig
C0013369|T047|PT|009.2|ICD9CM|Infectious diarrhea|Infectious diarrhea
C0013369|T047|AB|009.2|ICD9CM|Infectious diarrhea NOS|Infectious diarrhea NOS
C0152522|T047|AB|009.3|ICD9CM|Diarrhea of infect orig|Diarrhea of infect orig
C0152522|T047|PT|009.3|ICD9CM|Diarrhea of presumed infectious origin|Diarrhea of presumed infectious origin
C0152545|T047|HT|010|ICD9CM|Primary tuberculous infection|Primary tuberculous infection
C0041296|T047|HT|010-018.99|ICD9CM|TUBERCULOSIS|TUBERCULOSIS
C0152545|T047|HT|010.0|ICD9CM|Primary tuberculous infection|Primary tuberculous infection
C1812612|T047|AB|010.00|ICD9CM|Prim TB complex-unspec|Prim TB complex-unspec
C1812612|T047|PT|010.00|ICD9CM|Primary tuberculous infection, unspecified|Primary tuberculous infection, unspecified
C0374939|T047|AB|010.01|ICD9CM|Prim TB complex-no exam|Prim TB complex-no exam
C0374939|T047|PT|010.01|ICD9CM|Primary tuberculous infection, bacteriological or histological examination not done|Primary tuberculous infection, bacteriological or histological examination not done
C0374940|T047|AB|010.02|ICD9CM|Prim TB complex-exm unkn|Prim TB complex-exm unkn
C0374940|T047|PT|010.02|ICD9CM|Primary tuberculous infection, bacteriological or histological examination unknown (at present)|Primary tuberculous infection, bacteriological or histological examination unknown (at present)
C0374941|T047|AB|010.03|ICD9CM|Prim TB complex-micro dx|Prim TB complex-micro dx
C0374941|T047|PT|010.03|ICD9CM|Primary tuberculous infection, tubercle bacilli found (in sputum) by microscopy|Primary tuberculous infection, tubercle bacilli found (in sputum) by microscopy
C0374942|T047|AB|010.04|ICD9CM|Prim TB complex-cult dx|Prim TB complex-cult dx
C0374943|T047|AB|010.05|ICD9CM|Prim TB complex-histo dx|Prim TB complex-histo dx
C0374944|T047|AB|010.06|ICD9CM|Prim TB complex-oth test|Prim TB complex-oth test
C0152531|T047|HT|010.1|ICD9CM|Tuberculous pleurisy in primary progressive tuberculosis|Tuberculous pleurisy in primary progressive tuberculosis
C0374945|T047|AB|010.10|ICD9CM|Prim TB pleurisy-unspec|Prim TB pleurisy-unspec
C0374945|T047|PT|010.10|ICD9CM|Tuberculous pleurisy in primary progressive tuberculosis, unspecified|Tuberculous pleurisy in primary progressive tuberculosis, unspecified
C0152532|T047|AB|010.11|ICD9CM|Prim TB pleurisy-no exam|Prim TB pleurisy-no exam
C0152533|T047|AB|010.12|ICD9CM|Prim TB pleur-exam unkn|Prim TB pleur-exam unkn
C0152534|T047|AB|010.13|ICD9CM|Prim TB pleuris-micro dx|Prim TB pleuris-micro dx
C0152535|T047|AB|010.14|ICD9CM|Prim TB pleurisy-cult dx|Prim TB pleurisy-cult dx
C0152536|T047|AB|010.15|ICD9CM|Prim TB pleuris-histo dx|Prim TB pleuris-histo dx
C0152537|T047|AB|010.16|ICD9CM|Prim TB pleuris-oth test|Prim TB pleuris-oth test
C0152538|T047|HT|010.8|ICD9CM|Other primary progressive tuberculosis|Other primary progressive tuberculosis
C0374946|T047|PT|010.80|ICD9CM|Other primary progressive tuberculosis, unspecified|Other primary progressive tuberculosis, unspecified
C0374946|T047|AB|010.80|ICD9CM|Prim prog TB NEC-unspec|Prim prog TB NEC-unspec
C0152539|T047|PT|010.81|ICD9CM|Other primary progressive tuberculosis, bacteriological or histological examination not done|Other primary progressive tuberculosis, bacteriological or histological examination not done
C0152539|T047|AB|010.81|ICD9CM|Prim prog TB NEC-no exam|Prim prog TB NEC-no exam
C0152540|T047|AB|010.82|ICD9CM|Prim pr TB NEC-exam unkn|Prim pr TB NEC-exam unkn
C0152541|T047|PT|010.83|ICD9CM|Other primary progressive tuberculosis, tubercle bacilli found (in sputum) by microscopy|Other primary progressive tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152541|T047|AB|010.83|ICD9CM|Prim prg TB NEC-micro dx|Prim prg TB NEC-micro dx
C0152542|T047|AB|010.84|ICD9CM|Prim prog TB NEC-cult dx|Prim prog TB NEC-cult dx
C0152543|T047|AB|010.85|ICD9CM|Prim prg TB NEC-histo dx|Prim prg TB NEC-histo dx
C0152544|T047|AB|010.86|ICD9CM|Prim prg TB NEC-oth test|Prim prg TB NEC-oth test
C1812610|T047|HT|010.9|ICD9CM|Primary tuberculous infection, unspecified type|Primary tuberculous infection, unspecified type
C1812611|T047|AB|010.90|ICD9CM|Primary TB NOS-unspec|Primary TB NOS-unspec
C1812611|T047|PT|010.90|ICD9CM|Primary tuberculous infection, unspecified, unspecified|Primary tuberculous infection, unspecified, unspecified
C0152546|T047|AB|010.91|ICD9CM|Primary TB NOS-no exam|Primary TB NOS-no exam
C0152546|T047|PT|010.91|ICD9CM|Primary tuberculous infection, unspecified, bacteriological or histological examination not done|Primary tuberculous infection, unspecified, bacteriological or histological examination not done
C0152547|T047|AB|010.92|ICD9CM|Primary TB NOS-exam unkn|Primary TB NOS-exam unkn
C0152548|T033|AB|010.93|ICD9CM|Primary TB NOS-micro dx|Primary TB NOS-micro dx
C0152548|T033|PT|010.93|ICD9CM|Primary tuberculous infection, unspecified, tubercle bacilli found (in sputum) by microscopy|Primary tuberculous infection, unspecified, tubercle bacilli found (in sputum) by microscopy
C0152549|T047|AB|010.94|ICD9CM|Primary TB NOS-cult dx|Primary TB NOS-cult dx
C0152550|T047|AB|010.95|ICD9CM|Primary TB NOS-histo dx|Primary TB NOS-histo dx
C0152551|T047|AB|010.96|ICD9CM|Primary TB NOS-oth test|Primary TB NOS-oth test
C0041327|T047|HT|011|ICD9CM|Pulmonary tuberculosis|Pulmonary tuberculosis
C0152552|T047|HT|011.0|ICD9CM|Tuberculosis of lung, infiltrative|Tuberculosis of lung, infiltrative
C0152552|T047|AB|011.00|ICD9CM|TB lung infiltr-unspec|TB lung infiltr-unspec
C0152552|T047|PT|011.00|ICD9CM|Tuberculosis of lung, infiltrative, unspecified|Tuberculosis of lung, infiltrative, unspecified
C0152553|T047|AB|011.01|ICD9CM|TB lung infiltr-no exam|TB lung infiltr-no exam
C0152553|T047|PT|011.01|ICD9CM|Tuberculosis of lung, infiltrative, bacteriological or histological examination not done|Tuberculosis of lung, infiltrative, bacteriological or histological examination not done
C0152554|T047|AB|011.02|ICD9CM|TB lung infiltr-exm unkn|TB lung infiltr-exm unkn
C0152554|T047|PT|011.02|ICD9CM|Tuberculosis of lung, infiltrative, bacteriological or histological examination unknown (at present)|Tuberculosis of lung, infiltrative, bacteriological or histological examination unknown (at present)
C0152555|T047|AB|011.03|ICD9CM|TB lung infiltr-micro dx|TB lung infiltr-micro dx
C0152555|T047|PT|011.03|ICD9CM|Tuberculosis of lung, infiltrative, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of lung, infiltrative, tubercle bacilli found (in sputum) by microscopy
C0152556|T047|AB|011.04|ICD9CM|TB lung infiltr-cult dx|TB lung infiltr-cult dx
C0152557|T047|AB|011.05|ICD9CM|TB lung infiltr-histo dx|TB lung infiltr-histo dx
C0152558|T047|AB|011.06|ICD9CM|TB lung infiltr-oth test|TB lung infiltr-oth test
C0152559|T047|HT|011.1|ICD9CM|Tuberculosis of lung, nodular|Tuberculosis of lung, nodular
C0152559|T047|AB|011.10|ICD9CM|TB lung nodular-unspec|TB lung nodular-unspec
C0152559|T047|PT|011.10|ICD9CM|Tuberculosis of lung, nodular, unspecified|Tuberculosis of lung, nodular, unspecified
C0152560|T047|AB|011.11|ICD9CM|TB lung nodular-no exam|TB lung nodular-no exam
C0152560|T047|PT|011.11|ICD9CM|Tuberculosis of lung, nodular, bacteriological or histological examination not done|Tuberculosis of lung, nodular, bacteriological or histological examination not done
C0152561|T047|AB|011.12|ICD9CM|TB lung nodul-exam unkn|TB lung nodul-exam unkn
C0152561|T047|PT|011.12|ICD9CM|Tuberculosis of lung, nodular, bacteriological or histological examination unknown (at present)|Tuberculosis of lung, nodular, bacteriological or histological examination unknown (at present)
C0152562|T047|AB|011.13|ICD9CM|TB lung nodular-micro dx|TB lung nodular-micro dx
C0152562|T047|PT|011.13|ICD9CM|Tuberculosis of lung, nodular, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of lung, nodular, tubercle bacilli found (in sputum) by microscopy
C0152563|T047|AB|011.14|ICD9CM|TB lung nodular-cult dx|TB lung nodular-cult dx
C0152564|T047|AB|011.15|ICD9CM|TB lung nodular-histo dx|TB lung nodular-histo dx
C0152565|T047|AB|011.16|ICD9CM|TB lung nodular-oth test|TB lung nodular-oth test
C0152566|T047|HT|011.2|ICD9CM|Tuberculosis of lung with cavitation|Tuberculosis of lung with cavitation
C0152566|T047|AB|011.20|ICD9CM|TB lung w cavity-unspec|TB lung w cavity-unspec
C0152566|T047|PT|011.20|ICD9CM|Tuberculosis of lung with cavitation, unspecified|Tuberculosis of lung with cavitation, unspecified
C0152567|T047|AB|011.21|ICD9CM|TB lung w cavity-no exam|TB lung w cavity-no exam
C0152567|T047|PT|011.21|ICD9CM|Tuberculosis of lung with cavitation, bacteriological or histological examination not done|Tuberculosis of lung with cavitation, bacteriological or histological examination not done
C0152568|T047|AB|011.22|ICD9CM|TB lung cavity-exam unkn|TB lung cavity-exam unkn
C0152569|T047|AB|011.23|ICD9CM|TB lung w cavit-micro dx|TB lung w cavit-micro dx
C0152569|T047|PT|011.23|ICD9CM|Tuberculosis of lung with cavitation, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of lung with cavitation, tubercle bacilli found (in sputum) by microscopy
C0152570|T047|AB|011.24|ICD9CM|TB lung w cavity-cult dx|TB lung w cavity-cult dx
C0152571|T047|AB|011.25|ICD9CM|TB lung w cavit-histo dx|TB lung w cavit-histo dx
C0152572|T047|AB|011.26|ICD9CM|TB lung w cavit-oth test|TB lung w cavit-oth test
C0152573|T047|HT|011.3|ICD9CM|Tuberculosis of bronchus|Tuberculosis of bronchus
C0152573|T047|AB|011.30|ICD9CM|TB of bronchus-unspec|TB of bronchus-unspec
C0152573|T047|PT|011.30|ICD9CM|Tuberculosis of bronchus, unspecified|Tuberculosis of bronchus, unspecified
C0152574|T047|AB|011.31|ICD9CM|TB of bronchus-no exam|TB of bronchus-no exam
C0152574|T047|PT|011.31|ICD9CM|Tuberculosis of bronchus, bacteriological or histological examination not done|Tuberculosis of bronchus, bacteriological or histological examination not done
C0152575|T047|AB|011.32|ICD9CM|TB of bronchus-exam unkn|TB of bronchus-exam unkn
C0152575|T047|PT|011.32|ICD9CM|Tuberculosis of bronchus, bacteriological or histological examination unknown (at present)|Tuberculosis of bronchus, bacteriological or histological examination unknown (at present)
C0152576|T047|AB|011.33|ICD9CM|TB of bronchus-micro dx|TB of bronchus-micro dx
C0152576|T047|PT|011.33|ICD9CM|Tuberculosis of bronchus, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of bronchus, tubercle bacilli found (in sputum) by microscopy
C0152577|T047|AB|011.34|ICD9CM|TB of bronchus-cult dx|TB of bronchus-cult dx
C0152578|T047|AB|011.35|ICD9CM|TB of bronchus-histo dx|TB of bronchus-histo dx
C0152579|T047|AB|011.36|ICD9CM|TB of bronchus-oth test|TB of bronchus-oth test
C0041336|T047|HT|011.4|ICD9CM|Tuberculous fibrosis of lung|Tuberculous fibrosis of lung
C0041336|T047|AB|011.40|ICD9CM|TB lung fibrosis-unspec|TB lung fibrosis-unspec
C0041336|T047|PT|011.40|ICD9CM|Tuberculous fibrosis of lung, unspecified|Tuberculous fibrosis of lung, unspecified
C0152580|T047|AB|011.41|ICD9CM|TB lung fibrosis-no exam|TB lung fibrosis-no exam
C0152580|T047|PT|011.41|ICD9CM|Tuberculous fibrosis of lung, bacteriological or histological examination not done|Tuberculous fibrosis of lung, bacteriological or histological examination not done
C0152581|T047|AB|011.42|ICD9CM|TB lung fibros-exam unkn|TB lung fibros-exam unkn
C0152581|T047|PT|011.42|ICD9CM|Tuberculous fibrosis of lung, bacteriological or histological examination unknown (at present)|Tuberculous fibrosis of lung, bacteriological or histological examination unknown (at present)
C0152582|T047|AB|011.43|ICD9CM|TB lung fibros-micro dx|TB lung fibros-micro dx
C0152582|T047|PT|011.43|ICD9CM|Tuberculous fibrosis of lung, tubercle bacilli found (in sputum) by microscopy|Tuberculous fibrosis of lung, tubercle bacilli found (in sputum) by microscopy
C0152583|T047|AB|011.44|ICD9CM|TB lung fibrosis-cult dx|TB lung fibrosis-cult dx
C0152584|T047|AB|011.45|ICD9CM|TB lung fibros-histo dx|TB lung fibros-histo dx
C0152585|T047|AB|011.46|ICD9CM|TB lung fibros-oth test|TB lung fibros-oth test
C0152586|T047|HT|011.5|ICD9CM|Tuberculous bronchiectasis|Tuberculous bronchiectasis
C0152586|T047|AB|011.50|ICD9CM|TB bronchiectasis-unspec|TB bronchiectasis-unspec
C0152586|T047|PT|011.50|ICD9CM|Tuberculous bronchiectasis, unspecified|Tuberculous bronchiectasis, unspecified
C0152587|T047|AB|011.51|ICD9CM|TB bronchiect-no exam|TB bronchiect-no exam
C0152587|T047|PT|011.51|ICD9CM|Tuberculous bronchiectasis, bacteriological or histological examination not done|Tuberculous bronchiectasis, bacteriological or histological examination not done
C0152588|T047|AB|011.52|ICD9CM|TB bronchiect-exam unkn|TB bronchiect-exam unkn
C0152588|T047|PT|011.52|ICD9CM|Tuberculous bronchiectasis, bacteriological or histological examination unknown (at present)|Tuberculous bronchiectasis, bacteriological or histological examination unknown (at present)
C0152589|T047|AB|011.53|ICD9CM|TB bronchiect-micro dx|TB bronchiect-micro dx
C0152589|T047|PT|011.53|ICD9CM|Tuberculous bronchiectasis, tubercle bacilli found (in sputum) by microscopy|Tuberculous bronchiectasis, tubercle bacilli found (in sputum) by microscopy
C0152590|T047|AB|011.54|ICD9CM|TB bronchiect-cult dx|TB bronchiect-cult dx
C0152591|T047|AB|011.55|ICD9CM|TB bronchiect-histo dx|TB bronchiect-histo dx
C0152592|T047|AB|011.56|ICD9CM|TB bronchiect-oth test|TB bronchiect-oth test
C0275891|T047|HT|011.6|ICD9CM|Tuberculous pneumonia [any form]|Tuberculous pneumonia [any form]
C0374952|T047|AB|011.60|ICD9CM|TB pneumonia-unspec|TB pneumonia-unspec
C0374952|T047|PT|011.60|ICD9CM|Tuberculous pneumonia [any form], unspecified|Tuberculous pneumonia [any form], unspecified
C0152594|T047|AB|011.61|ICD9CM|TB pneumonia-no exam|TB pneumonia-no exam
C0152594|T047|PT|011.61|ICD9CM|Tuberculous pneumonia [any form], bacteriological or histological examination not done|Tuberculous pneumonia [any form], bacteriological or histological examination not done
C0152595|T047|AB|011.62|ICD9CM|TB pneumonia-exam unkn|TB pneumonia-exam unkn
C0152595|T047|PT|011.62|ICD9CM|Tuberculous pneumonia [any form], bacteriological or histological examination unknown (at present)|Tuberculous pneumonia [any form], bacteriological or histological examination unknown (at present)
C0152596|T047|AB|011.63|ICD9CM|TB pneumonia-micro dx|TB pneumonia-micro dx
C0152596|T047|PT|011.63|ICD9CM|Tuberculous pneumonia [any form], tubercle bacilli found (in sputum) by microscopy|Tuberculous pneumonia [any form], tubercle bacilli found (in sputum) by microscopy
C0152597|T047|AB|011.64|ICD9CM|TB pneumonia-cult dx|TB pneumonia-cult dx
C0152598|T047|AB|011.65|ICD9CM|TB pneumonia-histo dx|TB pneumonia-histo dx
C0152599|T047|AB|011.66|ICD9CM|TB pneumonia-oth test|TB pneumonia-oth test
C0152600|T047|HT|011.7|ICD9CM|Tuberculous pneumothorax|Tuberculous pneumothorax
C0152600|T047|AB|011.70|ICD9CM|TB pneumothorax-unspec|TB pneumothorax-unspec
C0152600|T047|PT|011.70|ICD9CM|Tuberculous pneumothorax, unspecified|Tuberculous pneumothorax, unspecified
C0152601|T047|AB|011.71|ICD9CM|TB pneumothorax-no exam|TB pneumothorax-no exam
C0152601|T047|PT|011.71|ICD9CM|Tuberculous pneumothorax, bacteriological or histological examination not done|Tuberculous pneumothorax, bacteriological or histological examination not done
C0152602|T047|AB|011.72|ICD9CM|TB pneumothorx-exam unkn|TB pneumothorx-exam unkn
C0152602|T047|PT|011.72|ICD9CM|Tuberculous pneumothorax, bacteriological or histological examination unknown (at present)|Tuberculous pneumothorax, bacteriological or histological examination unknown (at present)
C0152603|T047|AB|011.73|ICD9CM|TB pneumothorax-micro dx|TB pneumothorax-micro dx
C0152603|T047|PT|011.73|ICD9CM|Tuberculous pneumothorax, tubercle bacilli found (in sputum) by microscopy|Tuberculous pneumothorax, tubercle bacilli found (in sputum) by microscopy
C0152604|T047|AB|011.74|ICD9CM|TB pneumothorax-cult dx|TB pneumothorax-cult dx
C0152605|T047|AB|011.75|ICD9CM|TB pneumothorax-histo dx|TB pneumothorax-histo dx
C0152606|T047|AB|011.76|ICD9CM|TB pneumothorax-oth test|TB pneumothorax-oth test
C0152607|T047|HT|011.8|ICD9CM|Other specified pulmonary tuberculosis|Other specified pulmonary tuberculosis
C0374954|T047|PT|011.80|ICD9CM|Other specified pulmonary tuberculosis, unspecified|Other specified pulmonary tuberculosis, unspecified
C0374954|T047|AB|011.80|ICD9CM|Pulmonary TB NEC-unspec|Pulmonary TB NEC-unspec
C0152608|T047|PT|011.81|ICD9CM|Other specified pulmonary tuberculosis, bacteriological or histological examination not done|Other specified pulmonary tuberculosis, bacteriological or histological examination not done
C0152608|T047|AB|011.81|ICD9CM|Pulmonary TB NEC-no exam|Pulmonary TB NEC-no exam
C0152609|T047|AB|011.82|ICD9CM|Pulmon TB NEC-exam unkn|Pulmon TB NEC-exam unkn
C0152610|T047|PT|011.83|ICD9CM|Other specified pulmonary tuberculosis, tubercle bacilli found (in sputum) by microscopy|Other specified pulmonary tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152610|T047|AB|011.83|ICD9CM|Pulmon TB NEC-micro dx|Pulmon TB NEC-micro dx
C0152611|T047|AB|011.84|ICD9CM|Pulmon TB NEC-cult dx|Pulmon TB NEC-cult dx
C0152612|T047|AB|011.85|ICD9CM|Pulmon TB NEC-histo dx|Pulmon TB NEC-histo dx
C0152613|T047|AB|011.86|ICD9CM|Pulmon TB NEC-oth test|Pulmon TB NEC-oth test
C0041327|T047|HT|011.9|ICD9CM|Unspecified pulmonary tuberculosis|Unspecified pulmonary tuberculosis
C0041327|T047|AB|011.90|ICD9CM|Pulmonary TB NOS-unspec|Pulmonary TB NOS-unspec
C0041327|T047|PT|011.90|ICD9CM|Pulmonary tuberculosis, unspecified, unspecified|Pulmonary tuberculosis, unspecified, unspecified
C0152614|T047|AB|011.91|ICD9CM|Pulmonary TB NOS-no exam|Pulmonary TB NOS-no exam
C0152614|T047|PT|011.91|ICD9CM|Pulmonary tuberculosis, unspecified, bacteriological or histological examination not done|Pulmonary tuberculosis, unspecified, bacteriological or histological examination not done
C0152615|T047|AB|011.92|ICD9CM|Pulmon TB NOS-exam unkn|Pulmon TB NOS-exam unkn
C0152616|T047|AB|011.93|ICD9CM|Pulmon TB NOS-micro dx|Pulmon TB NOS-micro dx
C0152616|T047|PT|011.93|ICD9CM|Pulmonary tuberculosis, unspecified, tubercle bacilli found (in sputum) by microscopy|Pulmonary tuberculosis, unspecified, tubercle bacilli found (in sputum) by microscopy
C0152617|T047|AB|011.94|ICD9CM|Pulmon TB NOS-cult dx|Pulmon TB NOS-cult dx
C0152618|T047|AB|011.95|ICD9CM|Pulmon TB NOS-histo dx|Pulmon TB NOS-histo dx
C0152619|T047|AB|011.96|ICD9CM|Pulmon TB NOS-oth test|Pulmon TB NOS-oth test
C0152620|T047|HT|012|ICD9CM|Other respiratory tuberculosis|Other respiratory tuberculosis
C0041326|T047|HT|012.0|ICD9CM|Tuberculous pleurisy|Tuberculous pleurisy
C0041326|T047|AB|012.00|ICD9CM|TB pleurisy-unspec|TB pleurisy-unspec
C0041326|T047|PT|012.00|ICD9CM|Tuberculous pleurisy, unspecified|Tuberculous pleurisy, unspecified
C0152621|T047|AB|012.01|ICD9CM|TB pleurisy-no exam|TB pleurisy-no exam
C0152621|T047|PT|012.01|ICD9CM|Tuberculous pleurisy, bacteriological or histological examination not done|Tuberculous pleurisy, bacteriological or histological examination not done
C0152622|T047|AB|012.02|ICD9CM|TB pleurisy-exam unkn|TB pleurisy-exam unkn
C0152622|T047|PT|012.02|ICD9CM|Tuberculous pleurisy, bacteriological or histological examination unknown (at present)|Tuberculous pleurisy, bacteriological or histological examination unknown (at present)
C0152623|T047|AB|012.03|ICD9CM|TB pleurisy-micro dx|TB pleurisy-micro dx
C0152623|T047|PT|012.03|ICD9CM|Tuberculous pleurisy, tubercle bacilli found (in sputum) by microscopy|Tuberculous pleurisy, tubercle bacilli found (in sputum) by microscopy
C0152624|T047|AB|012.04|ICD9CM|TB pleurisy-cult dx|TB pleurisy-cult dx
C0152625|T047|AB|012.05|ICD9CM|TB pleurisy-histolog dx|TB pleurisy-histolog dx
C0152626|T047|AB|012.06|ICD9CM|TB pleurisy-oth test|TB pleurisy-oth test
C0152627|T047|HT|012.1|ICD9CM|Tuberculosis of intrathoracic lymph nodes|Tuberculosis of intrathoracic lymph nodes
C0152627|T047|AB|012.10|ICD9CM|TB thoracic nodes-unspec|TB thoracic nodes-unspec
C0152627|T047|PT|012.10|ICD9CM|Tuberculosis of intrathoracic lymph nodes, unspecified|Tuberculosis of intrathoracic lymph nodes, unspecified
C0152628|T047|AB|012.11|ICD9CM|TB thorax node-no exam|TB thorax node-no exam
C0152628|T047|PT|012.11|ICD9CM|Tuberculosis of intrathoracic lymph nodes, bacteriological or histological examination not done|Tuberculosis of intrathoracic lymph nodes, bacteriological or histological examination not done
C0152629|T047|AB|012.12|ICD9CM|TB thorax node-exam unkn|TB thorax node-exam unkn
C0152630|T047|AB|012.13|ICD9CM|TB thorax node-micro dx|TB thorax node-micro dx
C0152630|T047|PT|012.13|ICD9CM|Tuberculosis of intrathoracic lymph nodes, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of intrathoracic lymph nodes, tubercle bacilli found (in sputum) by microscopy
C0152631|T047|AB|012.14|ICD9CM|TB thorax node-cult dx|TB thorax node-cult dx
C0152632|T047|AB|012.15|ICD9CM|TB thorax node-histo dx|TB thorax node-histo dx
C0152633|T047|AB|012.16|ICD9CM|TB thorax node-oth test|TB thorax node-oth test
C0152634|T047|HT|012.2|ICD9CM|Isolated tracheal or bronchial tuberculosis|Isolated tracheal or bronchial tuberculosis
C0152634|T047|AB|012.20|ICD9CM|Isol tracheal tb-unspec|Isol tracheal tb-unspec
C0152634|T047|PT|012.20|ICD9CM|Isolated tracheal or bronchial tuberculosis, unspecified|Isolated tracheal or bronchial tuberculosis, unspecified
C0152635|T047|AB|012.21|ICD9CM|Isol tracheal tb-no exam|Isol tracheal tb-no exam
C0152635|T047|PT|012.21|ICD9CM|Isolated tracheal or bronchial tuberculosis, bacteriological or histological examination not done|Isolated tracheal or bronchial tuberculosis, bacteriological or histological examination not done
C0152636|T047|AB|012.22|ICD9CM|Isol trach tb-exam unkn|Isol trach tb-exam unkn
C0152637|T047|AB|012.23|ICD9CM|Isolat trach tb-micro dx|Isolat trach tb-micro dx
C0152637|T047|PT|012.23|ICD9CM|Isolated tracheal or bronchial tuberculosis, tubercle bacilli found (in sputum) by microscopy|Isolated tracheal or bronchial tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152638|T047|AB|012.24|ICD9CM|Isol tracheal tb-cult dx|Isol tracheal tb-cult dx
C0152639|T047|AB|012.25|ICD9CM|Isolat trach tb-histo dx|Isolat trach tb-histo dx
C0152640|T047|AB|012.26|ICD9CM|Isolat trach tb-oth test|Isolat trach tb-oth test
C0041315|T047|HT|012.3|ICD9CM|Tuberculous laryngitis|Tuberculous laryngitis
C0374955|T047|AB|012.30|ICD9CM|TB laryngitis-unspec|TB laryngitis-unspec
C0374955|T047|PT|012.30|ICD9CM|Tuberculous laryngitis, unspecified|Tuberculous laryngitis, unspecified
C0152641|T047|AB|012.31|ICD9CM|TB laryngitis-no exam|TB laryngitis-no exam
C0152641|T047|PT|012.31|ICD9CM|Tuberculous laryngitis, bacteriological or histological examination not done|Tuberculous laryngitis, bacteriological or histological examination not done
C0152642|T047|AB|012.32|ICD9CM|TB laryngitis-exam unkn|TB laryngitis-exam unkn
C0152642|T047|PT|012.32|ICD9CM|Tuberculous laryngitis, bacteriological or histological examination unknown (at present)|Tuberculous laryngitis, bacteriological or histological examination unknown (at present)
C0152643|T047|AB|012.33|ICD9CM|TB laryngitis-micro dx|TB laryngitis-micro dx
C0152643|T047|PT|012.33|ICD9CM|Tuberculous laryngitis, tubercle bacilli found (in sputum) by microscopy|Tuberculous laryngitis, tubercle bacilli found (in sputum) by microscopy
C0152644|T047|AB|012.34|ICD9CM|TB laryngitis-cult dx|TB laryngitis-cult dx
C0152645|T047|AB|012.35|ICD9CM|TB laryngitis-histo dx|TB laryngitis-histo dx
C0152646|T047|AB|012.36|ICD9CM|TB laryngitis-oth test|TB laryngitis-oth test
C0152647|T047|HT|012.8|ICD9CM|Other specified respiratory tuberculosis|Other specified respiratory tuberculosis
C0152647|T047|PT|012.80|ICD9CM|Other specified respiratory tuberculosis, unspecified|Other specified respiratory tuberculosis, unspecified
C0152647|T047|AB|012.80|ICD9CM|Resp TB NEC-unspec|Resp TB NEC-unspec
C0152648|T047|PT|012.81|ICD9CM|Other specified respiratory tuberculosis, bacteriological or histological examination not done|Other specified respiratory tuberculosis, bacteriological or histological examination not done
C0152648|T047|AB|012.81|ICD9CM|Resp TB NEC-no exam|Resp TB NEC-no exam
C0152649|T047|AB|012.82|ICD9CM|Resp TB NEC-exam unkn|Resp TB NEC-exam unkn
C0152650|T047|PT|012.83|ICD9CM|Other specified respiratory tuberculosis, tubercle bacilli found (in sputum) by microscopy|Other specified respiratory tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152650|T047|AB|012.83|ICD9CM|Resp TB NEC-micro dx|Resp TB NEC-micro dx
C0152651|T047|AB|012.84|ICD9CM|Resp TB NEC-cult dx|Resp TB NEC-cult dx
C0152652|T047|AB|012.85|ICD9CM|Resp TB NEC-histo dx|Resp TB NEC-histo dx
C0152653|T047|AB|012.86|ICD9CM|Resp TB NEC-oth test|Resp TB NEC-oth test
C0152654|T047|HT|013|ICD9CM|Tuberculosis of meninges and central nervous system|Tuberculosis of meninges and central nervous system
C0041318|T047|HT|013.0|ICD9CM|Tuberculous meningitis|Tuberculous meningitis
C0041318|T047|AB|013.00|ICD9CM|TB meningitis-unspec|TB meningitis-unspec
C0041318|T047|PT|013.00|ICD9CM|Tuberculous meningitis, unspecified|Tuberculous meningitis, unspecified
C0152655|T047|AB|013.01|ICD9CM|TB meningitis-no exam|TB meningitis-no exam
C0152655|T047|PT|013.01|ICD9CM|Tuberculous meningitis, bacteriological or histological examination not done|Tuberculous meningitis, bacteriological or histological examination not done
C0152656|T047|AB|013.02|ICD9CM|TB meningitis-exam unkn|TB meningitis-exam unkn
C0152656|T047|PT|013.02|ICD9CM|Tuberculous meningitis, bacteriological or histological examination unknown (at present)|Tuberculous meningitis, bacteriological or histological examination unknown (at present)
C0152657|T047|AB|013.03|ICD9CM|TB meningitis-micro dx|TB meningitis-micro dx
C0152657|T047|PT|013.03|ICD9CM|Tuberculous meningitis, tubercle bacilli found (in sputum) by microscopy|Tuberculous meningitis, tubercle bacilli found (in sputum) by microscopy
C0152658|T047|AB|013.04|ICD9CM|TB meningitis-cult dx|TB meningitis-cult dx
C0152659|T047|AB|013.05|ICD9CM|TB meningitis-histo dx|TB meningitis-histo dx
C0152660|T047|AB|013.06|ICD9CM|TB meningitis-oth test|TB meningitis-oth test
C0152661|T047|HT|013.1|ICD9CM|Tuberculoma of meninges|Tuberculoma of meninges
C0152661|T047|PT|013.10|ICD9CM|Tuberculoma of meninges, unspecified|Tuberculoma of meninges, unspecified
C0152661|T047|AB|013.10|ICD9CM|Tubrclma meninges-unspec|Tubrclma meninges-unspec
C0152662|T047|PT|013.11|ICD9CM|Tuberculoma of meninges, bacteriological or histological examination not done|Tuberculoma of meninges, bacteriological or histological examination not done
C0152662|T047|AB|013.11|ICD9CM|Tubrclma mening-no exam|Tubrclma mening-no exam
C0152663|T047|PT|013.12|ICD9CM|Tuberculoma of meninges, bacteriological or histological examination unknown (at present)|Tuberculoma of meninges, bacteriological or histological examination unknown (at present)
C0152663|T047|AB|013.12|ICD9CM|Tubrclma menin-exam unkn|Tubrclma menin-exam unkn
C0152664|T047|PT|013.13|ICD9CM|Tuberculoma of meninges, tubercle bacilli found (in sputum) by microscopy|Tuberculoma of meninges, tubercle bacilli found (in sputum) by microscopy
C0152664|T047|AB|013.13|ICD9CM|Tubrclma mening-micro dx|Tubrclma mening-micro dx
C0152665|T047|AB|013.14|ICD9CM|Tubrclma mening-cult dx|Tubrclma mening-cult dx
C0152666|T047|AB|013.15|ICD9CM|Tubrclma mening-histo dx|Tubrclma mening-histo dx
C0152667|T047|AB|013.16|ICD9CM|Tubrclma mening-oth test|Tubrclma mening-oth test
C0085388|T047|HT|013.2|ICD9CM|Tuberculoma of brain|Tuberculoma of brain
C0085388|T047|AB|013.20|ICD9CM|Tuberculoma brain-unspec|Tuberculoma brain-unspec
C0085388|T047|PT|013.20|ICD9CM|Tuberculoma of brain, unspecified|Tuberculoma of brain, unspecified
C0152669|T047|PT|013.21|ICD9CM|Tuberculoma of brain, bacteriological or histological examination not done|Tuberculoma of brain, bacteriological or histological examination not done
C0152669|T047|AB|013.21|ICD9CM|Tubrcloma brain-no exam|Tubrcloma brain-no exam
C0152670|T047|PT|013.22|ICD9CM|Tuberculoma of brain, bacteriological or histological examination unknown (at present)|Tuberculoma of brain, bacteriological or histological examination unknown (at present)
C0152670|T047|AB|013.22|ICD9CM|Tubrclma brain-exam unkn|Tubrclma brain-exam unkn
C0152671|T047|PT|013.23|ICD9CM|Tuberculoma of brain, tubercle bacilli found (in sputum) by microscopy|Tuberculoma of brain, tubercle bacilli found (in sputum) by microscopy
C0152671|T047|AB|013.23|ICD9CM|Tubrcloma brain-micro dx|Tubrcloma brain-micro dx
C0152672|T047|AB|013.24|ICD9CM|Tubrcloma brain-cult dx|Tubrcloma brain-cult dx
C0152673|T047|AB|013.25|ICD9CM|Tubrcloma brain-histo dx|Tubrcloma brain-histo dx
C0152674|T047|AB|013.26|ICD9CM|Tubrcloma brain-oth test|Tubrcloma brain-oth test
C2607948|T047|HT|013.3|ICD9CM|Tuberculous abscess of brain|Tuberculous abscess of brain
C0374958|T047|AB|013.30|ICD9CM|TB brain abscess-unspec|TB brain abscess-unspec
C0374958|T047|PT|013.30|ICD9CM|Tuberculous abscess of brain, unspecified|Tuberculous abscess of brain, unspecified
C0152676|T047|AB|013.31|ICD9CM|TB brain abscess-no exam|TB brain abscess-no exam
C0152676|T047|PT|013.31|ICD9CM|Tuberculous abscess of brain, bacteriological or histological examination not done|Tuberculous abscess of brain, bacteriological or histological examination not done
C0152677|T047|AB|013.32|ICD9CM|TB brain absc-exam unkn|TB brain absc-exam unkn
C0152677|T047|PT|013.32|ICD9CM|Tuberculous abscess of brain, bacteriological or histological examination unknown (at present)|Tuberculous abscess of brain, bacteriological or histological examination unknown (at present)
C0152678|T047|AB|013.33|ICD9CM|TB brain absc-micro dx|TB brain absc-micro dx
C0152678|T047|PT|013.33|ICD9CM|Tuberculous abscess of brain, tubercle bacilli found (in sputum) by microscopy|Tuberculous abscess of brain, tubercle bacilli found (in sputum) by microscopy
C0152679|T047|AB|013.34|ICD9CM|TB brain abscess-cult dx|TB brain abscess-cult dx
C0152680|T047|AB|013.35|ICD9CM|TB brain absc-histo dx|TB brain absc-histo dx
C0152681|T047|AB|013.36|ICD9CM|TB brain absc-oth test|TB brain absc-oth test
C0338439|T047|HT|013.4|ICD9CM|Tuberculoma of spinal cord|Tuberculoma of spinal cord
C0338439|T047|PT|013.40|ICD9CM|Tuberculoma of spinal cord, unspecified|Tuberculoma of spinal cord, unspecified
C0338439|T047|AB|013.40|ICD9CM|Tubrclma sp cord-unspec|Tubrclma sp cord-unspec
C0152683|T047|PT|013.41|ICD9CM|Tuberculoma of spinal cord, bacteriological or histological examination not done|Tuberculoma of spinal cord, bacteriological or histological examination not done
C0152683|T047|AB|013.41|ICD9CM|Tubrclma sp cord-no exam|Tubrclma sp cord-no exam
C0152684|T047|PT|013.42|ICD9CM|Tuberculoma of spinal cord, bacteriological or histological examination unknown (at present)|Tuberculoma of spinal cord, bacteriological or histological examination unknown (at present)
C0152684|T047|AB|013.42|ICD9CM|Tubrclma sp cd-exam unkn|Tubrclma sp cd-exam unkn
C0152685|T047|PT|013.43|ICD9CM|Tuberculoma of spinal cord, tubercle bacilli found (in sputum) by microscopy|Tuberculoma of spinal cord, tubercle bacilli found (in sputum) by microscopy
C0152685|T047|AB|013.43|ICD9CM|Tubrclma sp crd-micro dx|Tubrclma sp crd-micro dx
C0152686|T047|AB|013.44|ICD9CM|Tubrclma sp cord-cult dx|Tubrclma sp cord-cult dx
C0152687|T047|AB|013.45|ICD9CM|Tubrclma sp crd-histo dx|Tubrclma sp crd-histo dx
C0152688|T047|AB|013.46|ICD9CM|Tubrclma sp crd-oth test|Tubrclma sp crd-oth test
C0338439|T047|HT|013.5|ICD9CM|Tuberculous abscess of spinal cord|Tuberculous abscess of spinal cord
C0338439|T047|AB|013.50|ICD9CM|TB sp crd abscess-unspec|TB sp crd abscess-unspec
C0338439|T047|PT|013.50|ICD9CM|Tuberculous abscess of spinal cord, unspecified|Tuberculous abscess of spinal cord, unspecified
C0152690|T047|AB|013.51|ICD9CM|TB sp crd absc-no exam|TB sp crd absc-no exam
C0152690|T047|PT|013.51|ICD9CM|Tuberculous abscess of spinal cord, bacteriological or histological examination not done|Tuberculous abscess of spinal cord, bacteriological or histological examination not done
C0152691|T047|AB|013.52|ICD9CM|TB sp crd absc-exam unkn|TB sp crd absc-exam unkn
C0152691|T047|PT|013.52|ICD9CM|Tuberculous abscess of spinal cord, bacteriological or histological examination unknown (at present)|Tuberculous abscess of spinal cord, bacteriological or histological examination unknown (at present)
C0152692|T047|AB|013.53|ICD9CM|TB sp crd absc-micro dx|TB sp crd absc-micro dx
C0152692|T047|PT|013.53|ICD9CM|Tuberculous abscess of spinal cord, tubercle bacilli found (in sputum) by microscopy|Tuberculous abscess of spinal cord, tubercle bacilli found (in sputum) by microscopy
C0152693|T047|AB|013.54|ICD9CM|TB sp crd absc-cult dx|TB sp crd absc-cult dx
C0152694|T047|AB|013.55|ICD9CM|TB sp crd absc-histo dx|TB sp crd absc-histo dx
C0152695|T047|AB|013.56|ICD9CM|TB sp crd absc-oth test|TB sp crd absc-oth test
C0152696|T047|HT|013.6|ICD9CM|Tuberculous encephalitis or myelitis|Tuberculous encephalitis or myelitis
C0152696|T047|AB|013.60|ICD9CM|TB encephalitis-unspec|TB encephalitis-unspec
C0152696|T047|PT|013.60|ICD9CM|Tuberculous encephalitis or myelitis, unspecified|Tuberculous encephalitis or myelitis, unspecified
C0152697|T047|AB|013.61|ICD9CM|TB encephalitis-no exam|TB encephalitis-no exam
C0152697|T047|PT|013.61|ICD9CM|Tuberculous encephalitis or myelitis, bacteriological or histological examination not done|Tuberculous encephalitis or myelitis, bacteriological or histological examination not done
C0152698|T047|AB|013.62|ICD9CM|TB encephalit-exam unkn|TB encephalit-exam unkn
C0152699|T047|AB|013.63|ICD9CM|TB encephalitis-micro dx|TB encephalitis-micro dx
C0152699|T047|PT|013.63|ICD9CM|Tuberculous encephalitis or myelitis, tubercle bacilli found (in sputum) by microscopy|Tuberculous encephalitis or myelitis, tubercle bacilli found (in sputum) by microscopy
C0152700|T047|AB|013.64|ICD9CM|TB encephalitis-cult dx|TB encephalitis-cult dx
C0152701|T047|AB|013.65|ICD9CM|TB encephalitis-histo dx|TB encephalitis-histo dx
C0152702|T047|AB|013.66|ICD9CM|TB encephalitis-oth test|TB encephalitis-oth test
C0152703|T047|HT|013.8|ICD9CM|Other specified tuberculosis of central nervous system|Other specified tuberculosis of central nervous system
C0374959|T047|AB|013.80|ICD9CM|Cns TB NEC-unspec|Cns TB NEC-unspec
C0374959|T047|PT|013.80|ICD9CM|Other specified tuberculosis of central nervous system, unspecified|Other specified tuberculosis of central nervous system, unspecified
C0152704|T047|AB|013.81|ICD9CM|Cns TB NEC-no exam|Cns TB NEC-no exam
C0152705|T047|AB|013.82|ICD9CM|Cns TB NEC-exam unkn|Cns TB NEC-exam unkn
C0152706|T047|AB|013.83|ICD9CM|Cns TB NEC-micro dx|Cns TB NEC-micro dx
C0152707|T047|AB|013.84|ICD9CM|Cns TB NEC-cult dx|Cns TB NEC-cult dx
C0152708|T047|AB|013.85|ICD9CM|Cns TB NEC-histo dx|Cns TB NEC-histo dx
C0152709|T047|AB|013.86|ICD9CM|Cns TB NEC-oth test|Cns TB NEC-oth test
C0275904|T047|HT|013.9|ICD9CM|Unspecified tuberculosis of central nervous system|Unspecified tuberculosis of central nervous system
C0275904|T047|AB|013.90|ICD9CM|Cns TB NOS-unspec|Cns TB NOS-unspec
C0275904|T047|PT|013.90|ICD9CM|Unspecified tuberculosis of central nervous system, unspecified|Unspecified tuberculosis of central nervous system, unspecified
C0152711|T047|AB|013.91|ICD9CM|Cns TB NOS-no exam|Cns TB NOS-no exam
C0152712|T047|AB|013.92|ICD9CM|Cns TB NOS-exam unkn|Cns TB NOS-exam unkn
C0152713|T047|AB|013.93|ICD9CM|Cns TB NOS-micro dx|Cns TB NOS-micro dx
C0152713|T047|PT|013.93|ICD9CM|Unspecified tuberculosis of central nervous system, tubercle bacilli found (in sputum) by microscopy|Unspecified tuberculosis of central nervous system, tubercle bacilli found (in sputum) by microscopy
C0152714|T047|AB|013.94|ICD9CM|Cns TB NOS-cult dx|Cns TB NOS-cult dx
C0152715|T047|AB|013.95|ICD9CM|Cns TB NOS-histo dx|Cns TB NOS-histo dx
C0152716|T047|AB|013.96|ICD9CM|Cns TB NOS-oth test|Cns TB NOS-oth test
C0152717|T047|HT|014|ICD9CM|Tuberculosis of intestines, peritoneum, and mesenteric glands|Tuberculosis of intestines, peritoneum, and mesenteric glands
C0041325|T047|HT|014.0|ICD9CM|Tuberculous peritonitis|Tuberculous peritonitis
C0374961|T047|AB|014.00|ICD9CM|TB peritonitis-unspec|TB peritonitis-unspec
C0374961|T047|PT|014.00|ICD9CM|Tuberculous peritonitis, unspecified|Tuberculous peritonitis, unspecified
C0152718|T047|AB|014.01|ICD9CM|TB peritonitis-no exam|TB peritonitis-no exam
C0152718|T047|PT|014.01|ICD9CM|Tuberculous peritonitis, bacteriological or histological examination not done|Tuberculous peritonitis, bacteriological or histological examination not done
C0152719|T047|AB|014.02|ICD9CM|TB peritonitis-exam unkn|TB peritonitis-exam unkn
C0152719|T047|PT|014.02|ICD9CM|Tuberculous peritonitis, bacteriological or histological examination unknown (at present)|Tuberculous peritonitis, bacteriological or histological examination unknown (at present)
C0152720|T047|AB|014.03|ICD9CM|TB peritonitis-micro dx|TB peritonitis-micro dx
C0152720|T047|PT|014.03|ICD9CM|Tuberculous peritonitis, tubercle bacilli found (in sputum) by microscopy|Tuberculous peritonitis, tubercle bacilli found (in sputum) by microscopy
C0152721|T047|AB|014.04|ICD9CM|TB peritonitis-cult dx|TB peritonitis-cult dx
C0152722|T047|AB|014.05|ICD9CM|TB peritonitis-histo dx|TB peritonitis-histo dx
C0152723|T047|AB|014.06|ICD9CM|TB peritonitis-oth test|TB peritonitis-oth test
C0152724|T047|HT|014.8|ICD9CM|Tuberculosis of intestines and mesenteric glands|Tuberculosis of intestines and mesenteric glands
C0374962|T047|AB|014.80|ICD9CM|Intestinal TB NEC-unspec|Intestinal TB NEC-unspec
C0374962|T047|PT|014.80|ICD9CM|Other tuberculosis of intestines, peritoneum, and mesenteric glands, unspecified|Other tuberculosis of intestines, peritoneum, and mesenteric glands, unspecified
C0152725|T047|AB|014.81|ICD9CM|Intestin TB NEC-no exam|Intestin TB NEC-no exam
C0152726|T047|AB|014.82|ICD9CM|Intest TB NEC-exam unkn|Intest TB NEC-exam unkn
C0152727|T047|AB|014.83|ICD9CM|Intestin TB NEC-micro dx|Intestin TB NEC-micro dx
C0152728|T047|AB|014.84|ICD9CM|Intestin TB NEC-cult dx|Intestin TB NEC-cult dx
C0152729|T047|AB|014.85|ICD9CM|Intestin TB NEC-histo dx|Intestin TB NEC-histo dx
C0152730|T047|AB|014.86|ICD9CM|Intestin TB NEC-oth test|Intestin TB NEC-oth test
C0041324|T047|HT|015|ICD9CM|Tuberculosis of bones and joints|Tuberculosis of bones and joints
C0041330|T047|HT|015.0|ICD9CM|Tuberculosis of vertebral column|Tuberculosis of vertebral column
C0041330|T047|AB|015.00|ICD9CM|TB of vertebra-unspec|TB of vertebra-unspec
C0041330|T047|PT|015.00|ICD9CM|Tuberculosis of vertebral column, unspecified|Tuberculosis of vertebral column, unspecified
C0152731|T047|AB|015.01|ICD9CM|TB of vertebra-no exam|TB of vertebra-no exam
C0152731|T047|PT|015.01|ICD9CM|Tuberculosis of vertebral column, bacteriological or histological examination not done|Tuberculosis of vertebral column, bacteriological or histological examination not done
C0152732|T047|AB|015.02|ICD9CM|TB of vertebra-exam unkn|TB of vertebra-exam unkn
C0152732|T047|PT|015.02|ICD9CM|Tuberculosis of vertebral column, bacteriological or histological examination unknown (at present)|Tuberculosis of vertebral column, bacteriological or histological examination unknown (at present)
C0152733|T047|AB|015.03|ICD9CM|TB of vertebra-micro dx|TB of vertebra-micro dx
C0152733|T047|PT|015.03|ICD9CM|Tuberculosis of vertebral column, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of vertebral column, tubercle bacilli found (in sputum) by microscopy
C0152734|T047|AB|015.04|ICD9CM|TB of vertebra-cult dx|TB of vertebra-cult dx
C0152735|T047|AB|015.05|ICD9CM|TB of vertebra-histo dx|TB of vertebra-histo dx
C0152736|T047|AB|015.06|ICD9CM|TB of vertebra-oth test|TB of vertebra-oth test
C0152737|T047|HT|015.1|ICD9CM|Tuberculosis of hip|Tuberculosis of hip
C0374963|T047|AB|015.10|ICD9CM|TB of hip-unspec|TB of hip-unspec
C0374963|T047|PT|015.10|ICD9CM|Tuberculosis of hip, unspecified|Tuberculosis of hip, unspecified
C0152738|T047|AB|015.11|ICD9CM|TB of hip-no exam|TB of hip-no exam
C0152738|T047|PT|015.11|ICD9CM|Tuberculosis of hip, bacteriological or histological examination not done|Tuberculosis of hip, bacteriological or histological examination not done
C0152739|T047|AB|015.12|ICD9CM|TB of hip-exam unkn|TB of hip-exam unkn
C0152739|T047|PT|015.12|ICD9CM|Tuberculosis of hip, bacteriological or histological examination unknown (at present)|Tuberculosis of hip, bacteriological or histological examination unknown (at present)
C0152740|T047|AB|015.13|ICD9CM|TB of hip-micro dx|TB of hip-micro dx
C0152740|T047|PT|015.13|ICD9CM|Tuberculosis of hip, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of hip, tubercle bacilli found (in sputum) by microscopy
C0152741|T047|AB|015.14|ICD9CM|TB of hip-cult dx|TB of hip-cult dx
C0152742|T047|AB|015.15|ICD9CM|TB of hip-histo dx|TB of hip-histo dx
C0152743|T047|AB|015.16|ICD9CM|TB of hip-oth test|TB of hip-oth test
C0152744|T047|HT|015.2|ICD9CM|Tuberculosis of knee|Tuberculosis of knee
C0374964|T047|AB|015.20|ICD9CM|TB of knee-unspec|TB of knee-unspec
C0374964|T047|PT|015.20|ICD9CM|Tuberculosis of knee, unspecified|Tuberculosis of knee, unspecified
C0152745|T047|AB|015.21|ICD9CM|TB of knee-no exam|TB of knee-no exam
C0152745|T047|PT|015.21|ICD9CM|Tuberculosis of knee, bacteriological or histological examination not done|Tuberculosis of knee, bacteriological or histological examination not done
C0152746|T047|AB|015.22|ICD9CM|TB of knee-exam unkn|TB of knee-exam unkn
C0152746|T047|PT|015.22|ICD9CM|Tuberculosis of knee, bacteriological or histological examination unknown (at present)|Tuberculosis of knee, bacteriological or histological examination unknown (at present)
C0152747|T047|AB|015.23|ICD9CM|TB of knee-micro dx|TB of knee-micro dx
C0152747|T047|PT|015.23|ICD9CM|Tuberculosis of knee, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of knee, tubercle bacilli found (in sputum) by microscopy
C0152748|T047|AB|015.24|ICD9CM|TB of knee-cult dx|TB of knee-cult dx
C0152749|T047|AB|015.25|ICD9CM|TB of knee-histo dx|TB of knee-histo dx
C0152750|T047|AB|015.26|ICD9CM|TB of knee-oth test|TB of knee-oth test
C0347900|T047|HT|015.5|ICD9CM|Tuberculosis of limb bones|Tuberculosis of limb bones
C0347900|T047|AB|015.50|ICD9CM|TB of limb bones-unspec|TB of limb bones-unspec
C0347900|T047|PT|015.50|ICD9CM|Tuberculosis of limb bones, unspecified|Tuberculosis of limb bones, unspecified
C0152752|T047|AB|015.51|ICD9CM|TB limb bones-no exam|TB limb bones-no exam
C0152752|T047|PT|015.51|ICD9CM|Tuberculosis of limb bones, bacteriological or histological examination not done|Tuberculosis of limb bones, bacteriological or histological examination not done
C0152753|T047|AB|015.52|ICD9CM|TB limb bones-exam unkn|TB limb bones-exam unkn
C0152753|T047|PT|015.52|ICD9CM|Tuberculosis of limb bones, bacteriological or histological examination unknown (at present)|Tuberculosis of limb bones, bacteriological or histological examination unknown (at present)
C0152754|T047|AB|015.53|ICD9CM|TB limb bones-micro dx|TB limb bones-micro dx
C0152754|T047|PT|015.53|ICD9CM|Tuberculosis of limb bones, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of limb bones, tubercle bacilli found (in sputum) by microscopy
C0152755|T047|AB|015.54|ICD9CM|TB limb bones-cult dx|TB limb bones-cult dx
C0152756|T047|AB|015.55|ICD9CM|TB limb bones-histo dx|TB limb bones-histo dx
C0152757|T047|AB|015.56|ICD9CM|TB limb bones-oth test|TB limb bones-oth test
C0275956|T047|HT|015.6|ICD9CM|Tuberculosis of mastoid|Tuberculosis of mastoid
C0374965|T047|AB|015.60|ICD9CM|TB of mastoid-unspec|TB of mastoid-unspec
C0374965|T047|PT|015.60|ICD9CM|Tuberculosis of mastoid, unspecified|Tuberculosis of mastoid, unspecified
C0152759|T047|AB|015.61|ICD9CM|TB of mastoid-no exam|TB of mastoid-no exam
C0152759|T047|PT|015.61|ICD9CM|Tuberculosis of mastoid, bacteriological or histological examination not done|Tuberculosis of mastoid, bacteriological or histological examination not done
C0152760|T047|AB|015.62|ICD9CM|TB of mastoid-exam unkn|TB of mastoid-exam unkn
C0152760|T047|PT|015.62|ICD9CM|Tuberculosis of mastoid, bacteriological or histological examination unknown (at present)|Tuberculosis of mastoid, bacteriological or histological examination unknown (at present)
C0152761|T047|AB|015.63|ICD9CM|TB of mastoid-micro dx|TB of mastoid-micro dx
C0152761|T047|PT|015.63|ICD9CM|Tuberculosis of mastoid, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of mastoid, tubercle bacilli found (in sputum) by microscopy
C0152762|T047|AB|015.64|ICD9CM|TB of mastoid-cult dx|TB of mastoid-cult dx
C0152763|T047|AB|015.65|ICD9CM|TB of mastoid-histo dx|TB of mastoid-histo dx
C0152764|T047|AB|015.66|ICD9CM|TB of mastoid-oth test|TB of mastoid-oth test
C0152765|T047|HT|015.7|ICD9CM|Tuberculosis of other specified bone|Tuberculosis of other specified bone
C0374966|T047|AB|015.70|ICD9CM|TB of bone NEC-unspec|TB of bone NEC-unspec
C0374966|T047|PT|015.70|ICD9CM|Tuberculosis of other specified bone, unspecified|Tuberculosis of other specified bone, unspecified
C0152766|T047|AB|015.71|ICD9CM|TB of bone NEC-no exam|TB of bone NEC-no exam
C0152766|T047|PT|015.71|ICD9CM|Tuberculosis of other specified bone, bacteriological or histological examination not done|Tuberculosis of other specified bone, bacteriological or histological examination not done
C0152767|T047|AB|015.72|ICD9CM|TB of bone NEC-exam unkn|TB of bone NEC-exam unkn
C0152768|T047|AB|015.73|ICD9CM|TB of bone NEC-micro dx|TB of bone NEC-micro dx
C0152768|T047|PT|015.73|ICD9CM|Tuberculosis of other specified bone, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of other specified bone, tubercle bacilli found (in sputum) by microscopy
C0152769|T047|AB|015.74|ICD9CM|TB of bone NEC-cult dx|TB of bone NEC-cult dx
C0152770|T047|AB|015.75|ICD9CM|TB of bone NEC-histo dx|TB of bone NEC-histo dx
C0152771|T047|AB|015.76|ICD9CM|TB of bone NEC-oth test|TB of bone NEC-oth test
C0152772|T047|HT|015.8|ICD9CM|Tuberculosis of other specified joint|Tuberculosis of other specified joint
C0374967|T047|AB|015.80|ICD9CM|TB of joint NEC-unspec|TB of joint NEC-unspec
C0374967|T047|PT|015.80|ICD9CM|Tuberculosis of other specified joint, unspecified|Tuberculosis of other specified joint, unspecified
C0152773|T047|AB|015.81|ICD9CM|TB of joint NEC-no exam|TB of joint NEC-no exam
C0152773|T047|PT|015.81|ICD9CM|Tuberculosis of other specified joint, bacteriological or histological examination not done|Tuberculosis of other specified joint, bacteriological or histological examination not done
C0152774|T047|AB|015.82|ICD9CM|TB joint NEC-exam unkn|TB joint NEC-exam unkn
C0152775|T047|AB|015.83|ICD9CM|TB of joint NEC-micro dx|TB of joint NEC-micro dx
C0152775|T047|PT|015.83|ICD9CM|Tuberculosis of other specified joint, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of other specified joint, tubercle bacilli found (in sputum) by microscopy
C0152776|T047|AB|015.84|ICD9CM|TB of joint NEC-cult dx|TB of joint NEC-cult dx
C0152777|T047|AB|015.85|ICD9CM|TB of joint NEC-histo dx|TB of joint NEC-histo dx
C0152778|T047|AB|015.86|ICD9CM|TB of joint NEC-oth test|TB of joint NEC-oth test
C0041324|T047|HT|015.9|ICD9CM|Tuberculosis of unspecified bones and joints|Tuberculosis of unspecified bones and joints
C0374968|T047|AB|015.90|ICD9CM|TB bone/joint NOS-unspec|TB bone/joint NOS-unspec
C0374968|T047|PT|015.90|ICD9CM|Tuberculosis of unspecified bones and joints, unspecified|Tuberculosis of unspecified bones and joints, unspecified
C0152780|T047|AB|015.91|ICD9CM|TB bone/jt NOS-no exam|TB bone/jt NOS-no exam
C0152780|T047|PT|015.91|ICD9CM|Tuberculosis of unspecified bones and joints, bacteriological or histological examination not done|Tuberculosis of unspecified bones and joints, bacteriological or histological examination not done
C0152781|T047|AB|015.92|ICD9CM|TB bone/jt NOS-exam unkn|TB bone/jt NOS-exam unkn
C0152782|T047|AB|015.93|ICD9CM|TB bone/jt NOS-micro dx|TB bone/jt NOS-micro dx
C0152782|T047|PT|015.93|ICD9CM|Tuberculosis of unspecified bones and joints, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of unspecified bones and joints, tubercle bacilli found (in sputum) by microscopy
C0152783|T047|AB|015.94|ICD9CM|TB bone/jt NOS-cult dx|TB bone/jt NOS-cult dx
C0152784|T047|AB|015.95|ICD9CM|TB bone/jt NOS-histo dx|TB bone/jt NOS-histo dx
C0152785|T047|AB|015.96|ICD9CM|TB bone/jt NOS-oth test|TB bone/jt NOS-oth test
C0041333|T047|HT|016|ICD9CM|Tuberculosis of genitourinary system|Tuberculosis of genitourinary system
C0041328|T047|HT|016.0|ICD9CM|Tuberculosis of kidney|Tuberculosis of kidney
C0041328|T047|AB|016.00|ICD9CM|TB of kidney-unspec|TB of kidney-unspec
C0041328|T047|PT|016.00|ICD9CM|Tuberculosis of kidney, unspecified|Tuberculosis of kidney, unspecified
C0152787|T047|AB|016.01|ICD9CM|TB of kidney-no exam|TB of kidney-no exam
C0152787|T047|PT|016.01|ICD9CM|Tuberculosis of kidney, bacteriological or histological examination not done|Tuberculosis of kidney, bacteriological or histological examination not done
C0152788|T047|AB|016.02|ICD9CM|TB of kidney-exam unkn|TB of kidney-exam unkn
C0152788|T047|PT|016.02|ICD9CM|Tuberculosis of kidney, bacteriological or histological examination unknown (at present)|Tuberculosis of kidney, bacteriological or histological examination unknown (at present)
C0152789|T047|AB|016.03|ICD9CM|TB of kidney-micro dx|TB of kidney-micro dx
C0152789|T047|PT|016.03|ICD9CM|Tuberculosis of kidney, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of kidney, tubercle bacilli found (in sputum) by microscopy
C0152790|T047|AB|016.04|ICD9CM|TB of kidney-cult dx|TB of kidney-cult dx
C0152791|T047|AB|016.05|ICD9CM|TB of kidney-histo dx|TB of kidney-histo dx
C0152792|T047|AB|016.06|ICD9CM|TB of kidney-oth test|TB of kidney-oth test
C0152793|T047|HT|016.1|ICD9CM|Tuberculosis of bladder|Tuberculosis of bladder
C0152793|T047|AB|016.10|ICD9CM|TB of bladder-unspec|TB of bladder-unspec
C0152793|T047|PT|016.10|ICD9CM|Tuberculosis of bladder, unspecified|Tuberculosis of bladder, unspecified
C0152794|T047|AB|016.11|ICD9CM|TB of bladder-no exam|TB of bladder-no exam
C0152794|T047|PT|016.11|ICD9CM|Tuberculosis of bladder, bacteriological or histological examination not done|Tuberculosis of bladder, bacteriological or histological examination not done
C0152795|T047|AB|016.12|ICD9CM|TB of bladder-exam unkn|TB of bladder-exam unkn
C0152795|T047|PT|016.12|ICD9CM|Tuberculosis of bladder, bacteriological or histological examination unknown (at present)|Tuberculosis of bladder, bacteriological or histological examination unknown (at present)
C0152796|T047|AB|016.13|ICD9CM|TB of bladder-micro dx|TB of bladder-micro dx
C0152796|T047|PT|016.13|ICD9CM|Tuberculosis of bladder, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of bladder, tubercle bacilli found (in sputum) by microscopy
C0152797|T047|AB|016.14|ICD9CM|TB of bladder-cult dx|TB of bladder-cult dx
C0152798|T047|AB|016.15|ICD9CM|TB of bladder-histo dx|TB of bladder-histo dx
C0152799|T047|AB|016.16|ICD9CM|TB of bladder-oth test|TB of bladder-oth test
C0152800|T047|HT|016.2|ICD9CM|Tuberculosis of ureter|Tuberculosis of ureter
C0374969|T047|AB|016.20|ICD9CM|TB of ureter-unspec|TB of ureter-unspec
C0374969|T047|PT|016.20|ICD9CM|Tuberculosis of ureter, unspecified|Tuberculosis of ureter, unspecified
C0152801|T047|AB|016.21|ICD9CM|TB of ureter-no exam|TB of ureter-no exam
C0152801|T047|PT|016.21|ICD9CM|Tuberculosis of ureter, bacteriological or histological examination not done|Tuberculosis of ureter, bacteriological or histological examination not done
C0152802|T047|AB|016.22|ICD9CM|TB of ureter-exam unkn|TB of ureter-exam unkn
C0152802|T047|PT|016.22|ICD9CM|Tuberculosis of ureter, bacteriological or histological examination unknown (at present)|Tuberculosis of ureter, bacteriological or histological examination unknown (at present)
C0152803|T047|AB|016.23|ICD9CM|TB of ureter-micro dx|TB of ureter-micro dx
C0152803|T047|PT|016.23|ICD9CM|Tuberculosis of ureter, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of ureter, tubercle bacilli found (in sputum) by microscopy
C0152804|T047|AB|016.24|ICD9CM|TB of ureter-cult dx|TB of ureter-cult dx
C0152805|T047|AB|016.25|ICD9CM|TB of ureter-histo dx|TB of ureter-histo dx
C0152806|T047|AB|016.26|ICD9CM|TB of ureter-oth test|TB of ureter-oth test
C0041332|T047|HT|016.3|ICD9CM|Tuberculosis of other urinary organs|Tuberculosis of other urinary organs
C0374970|T047|AB|016.30|ICD9CM|TB urinary NEC-unspec|TB urinary NEC-unspec
C0374970|T047|PT|016.30|ICD9CM|Tuberculosis of other urinary organs, unspecified|Tuberculosis of other urinary organs, unspecified
C0152808|T047|AB|016.31|ICD9CM|TB urinary NEC-no exam|TB urinary NEC-no exam
C0152808|T047|PT|016.31|ICD9CM|Tuberculosis of other urinary organs, bacteriological or histological examination not done|Tuberculosis of other urinary organs, bacteriological or histological examination not done
C0152809|T047|AB|016.32|ICD9CM|TB urinary NEC-exam unkn|TB urinary NEC-exam unkn
C0152810|T047|AB|016.33|ICD9CM|TB urinary NEC-micro dx|TB urinary NEC-micro dx
C0152810|T047|PT|016.33|ICD9CM|Tuberculosis of other urinary organs, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of other urinary organs, tubercle bacilli found (in sputum) by microscopy
C0152811|T047|AB|016.34|ICD9CM|TB urinary NEC-cult dx|TB urinary NEC-cult dx
C0152812|T047|AB|016.35|ICD9CM|TB urinary NEC-histo dx|TB urinary NEC-histo dx
C0152813|T047|AB|016.36|ICD9CM|TB urinary NEC-oth test|TB urinary NEC-oth test
C0152814|T047|HT|016.4|ICD9CM|Tuberculosis of epididymis|Tuberculosis of epididymis
C0374971|T047|AB|016.40|ICD9CM|TB epididymis-unspec|TB epididymis-unspec
C0374971|T047|PT|016.40|ICD9CM|Tuberculosis of epididymis, unspecified|Tuberculosis of epididymis, unspecified
C0152815|T047|AB|016.41|ICD9CM|TB epididymis-no exam|TB epididymis-no exam
C0152815|T047|PT|016.41|ICD9CM|Tuberculosis of epididymis, bacteriological or histological examination not done|Tuberculosis of epididymis, bacteriological or histological examination not done
C0152816|T047|AB|016.42|ICD9CM|TB epididymis-exam unkn|TB epididymis-exam unkn
C0152816|T047|PT|016.42|ICD9CM|Tuberculosis of epididymis, bacteriological or histological examination unknown (at present)|Tuberculosis of epididymis, bacteriological or histological examination unknown (at present)
C0152817|T047|AB|016.43|ICD9CM|TB epididymis-micro dx|TB epididymis-micro dx
C0152817|T047|PT|016.43|ICD9CM|Tuberculosis of epididymis, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of epididymis, tubercle bacilli found (in sputum) by microscopy
C0152818|T047|AB|016.44|ICD9CM|TB epididymis-cult dx|TB epididymis-cult dx
C0152819|T047|AB|016.45|ICD9CM|TB epididymis-histo dx|TB epididymis-histo dx
C0152820|T047|AB|016.46|ICD9CM|TB epididymis-oth test|TB epididymis-oth test
C0152821|T047|HT|016.5|ICD9CM|Tuberculosis of other male genital organs|Tuberculosis of other male genital organs
C0152821|T047|AB|016.50|ICD9CM|TB male genit NEC-unspec|TB male genit NEC-unspec
C0152821|T047|PT|016.50|ICD9CM|Tuberculosis of other male genital organs, unspecified|Tuberculosis of other male genital organs, unspecified
C0152822|T047|AB|016.51|ICD9CM|TB male gen NEC-no exam|TB male gen NEC-no exam
C0152822|T047|PT|016.51|ICD9CM|Tuberculosis of other male genital organs, bacteriological or histological examination not done|Tuberculosis of other male genital organs, bacteriological or histological examination not done
C0152823|T047|AB|016.52|ICD9CM|TB male gen NEC-ex unkn|TB male gen NEC-ex unkn
C0152824|T047|AB|016.53|ICD9CM|TB male gen NEC-micro dx|TB male gen NEC-micro dx
C0152824|T047|PT|016.53|ICD9CM|Tuberculosis of other male genital organs, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of other male genital organs, tubercle bacilli found (in sputum) by microscopy
C0152825|T047|AB|016.54|ICD9CM|TB male gen NEC-cult dx|TB male gen NEC-cult dx
C0152826|T047|AB|016.55|ICD9CM|TB male gen NEC-histo dx|TB male gen NEC-histo dx
C0152827|T047|AB|016.56|ICD9CM|TB male gen NEC-oth test|TB male gen NEC-oth test
C0152828|T047|HT|016.6|ICD9CM|Tuberculous oophoritis and salpingitis|Tuberculous oophoritis and salpingitis
C0374972|T047|AB|016.60|ICD9CM|TB ovary & tube-unspec|TB ovary & tube-unspec
C0374972|T047|PT|016.60|ICD9CM|Tuberculous oophoritis and salpingitis, unspecified|Tuberculous oophoritis and salpingitis, unspecified
C0152829|T047|AB|016.61|ICD9CM|TB ovary & tube-no exam|TB ovary & tube-no exam
C0152829|T047|PT|016.61|ICD9CM|Tuberculous oophoritis and salpingitis, bacteriological or histological examination not done|Tuberculous oophoritis and salpingitis, bacteriological or histological examination not done
C0152830|T047|AB|016.62|ICD9CM|TB ovary/tube-exam unkn|TB ovary/tube-exam unkn
C0152831|T047|AB|016.63|ICD9CM|TB ovary & tube-micro dx|TB ovary & tube-micro dx
C0152831|T047|PT|016.63|ICD9CM|Tuberculous oophoritis and salpingitis, tubercle bacilli found (in sputum) by microscopy|Tuberculous oophoritis and salpingitis, tubercle bacilli found (in sputum) by microscopy
C0152832|T047|AB|016.64|ICD9CM|TB ovary & tube-cult dx|TB ovary & tube-cult dx
C0152833|T047|AB|016.65|ICD9CM|TB ovary & tube-histo dx|TB ovary & tube-histo dx
C0152834|T047|AB|016.66|ICD9CM|TB ovary & tube-oth test|TB ovary & tube-oth test
C0152835|T047|HT|016.7|ICD9CM|Tuberculosis of other female genital organs|Tuberculosis of other female genital organs
C0152835|T047|AB|016.70|ICD9CM|TB female gen NEC-unspec|TB female gen NEC-unspec
C0152835|T047|PT|016.70|ICD9CM|Tuberculosis of other female genital organs, unspecified|Tuberculosis of other female genital organs, unspecified
C0152836|T047|AB|016.71|ICD9CM|TB fem gen NEC-no exam|TB fem gen NEC-no exam
C0152836|T047|PT|016.71|ICD9CM|Tuberculosis of other female genital organs, bacteriological or histological examination not done|Tuberculosis of other female genital organs, bacteriological or histological examination not done
C0152837|T047|AB|016.72|ICD9CM|TB fem gen NEC-exam unkn|TB fem gen NEC-exam unkn
C0152838|T047|AB|016.73|ICD9CM|TB fem gen NEC-micro dx|TB fem gen NEC-micro dx
C0152838|T047|PT|016.73|ICD9CM|Tuberculosis of other female genital organs, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of other female genital organs, tubercle bacilli found (in sputum) by microscopy
C0152839|T047|AB|016.74|ICD9CM|TB fem gen NEC-cult dx|TB fem gen NEC-cult dx
C0152840|T047|AB|016.75|ICD9CM|TB fem gen NEC-histo dx|TB fem gen NEC-histo dx
C0152841|T047|AB|016.76|ICD9CM|TB fem gen NEC-oth test|TB fem gen NEC-oth test
C0041333|T047|HT|016.9|ICD9CM|Genitourinary tuberculosis, unspecified|Genitourinary tuberculosis, unspecified
C0374973|T047|PT|016.90|ICD9CM|Genitourinary tuberculosis, unspecified, unspecified|Genitourinary tuberculosis, unspecified, unspecified
C0374973|T047|AB|016.90|ICD9CM|Gu TB NOS-unspec|Gu TB NOS-unspec
C0152843|T047|PT|016.91|ICD9CM|Genitourinary tuberculosis, unspecified, bacteriological or histological examination not done|Genitourinary tuberculosis, unspecified, bacteriological or histological examination not done
C0152843|T047|AB|016.91|ICD9CM|Gu TB NOS-no exam|Gu TB NOS-no exam
C0152844|T047|AB|016.92|ICD9CM|Gu TB NOS-exam unkn|Gu TB NOS-exam unkn
C0152845|T047|PT|016.93|ICD9CM|Genitourinary tuberculosis, unspecified, tubercle bacilli found (in sputum) by microscopy|Genitourinary tuberculosis, unspecified, tubercle bacilli found (in sputum) by microscopy
C0152845|T047|AB|016.93|ICD9CM|Gu TB NOS-micro dx|Gu TB NOS-micro dx
C0152846|T047|AB|016.94|ICD9CM|Gu TB NOS-cult dx|Gu TB NOS-cult dx
C0152847|T047|AB|016.95|ICD9CM|Gu TB NOS-histo dx|Gu TB NOS-histo dx
C0152848|T047|AB|016.96|ICD9CM|Gu TB NOS-oth test|Gu TB NOS-oth test
C0041300|T047|HT|017|ICD9CM|Tuberculosis of other organs|Tuberculosis of other organs
C0374974|T047|HT|017.0|ICD9CM|Tuberculosis of skin and subcutaneous cellular tissue|Tuberculosis of skin and subcutaneous cellular tissue
C0374974|T047|AB|017.00|ICD9CM|TB skin/subcutan-unspec|TB skin/subcutan-unspec
C0374974|T047|PT|017.00|ICD9CM|Tuberculosis of skin and subcutaneous cellular tissue, unspecified|Tuberculosis of skin and subcutaneous cellular tissue, unspecified
C0152849|T047|AB|017.01|ICD9CM|TB skin/subcut-no exam|TB skin/subcut-no exam
C0152850|T047|AB|017.02|ICD9CM|TB skin/subcut-exam unkn|TB skin/subcut-exam unkn
C0152851|T047|AB|017.03|ICD9CM|TB skin/subcut-micro dx|TB skin/subcut-micro dx
C0152852|T047|AB|017.04|ICD9CM|TB skin/subcut-cult dx|TB skin/subcut-cult dx
C0152853|T047|AB|017.05|ICD9CM|TB skin/subcut-histo dx|TB skin/subcut-histo dx
C0152854|T047|AB|017.06|ICD9CM|TB skin/subcut-oth test|TB skin/subcut-oth test
C0014744|T047|HT|017.1|ICD9CM|Erythema nodosum with hypersensitivity reaction in tuberculosis|Erythema nodosum with hypersensitivity reaction in tuberculosis
C0014744|T047|AB|017.10|ICD9CM|Erythema nodos tb-unspec|Erythema nodos tb-unspec
C0014744|T047|PT|017.10|ICD9CM|Erythema nodosum with hypersensitivity reaction in tuberculosis, unspecified|Erythema nodosum with hypersensitivity reaction in tuberculosis, unspecified
C0152855|T047|AB|017.11|ICD9CM|Erythem nodos tb-no exam|Erythem nodos tb-no exam
C0152856|T047|AB|017.12|ICD9CM|Erythem nod tb-exam unkn|Erythem nod tb-exam unkn
C0152857|T047|AB|017.13|ICD9CM|Erythem nod tb-micro dx|Erythem nod tb-micro dx
C0152858|T047|AB|017.14|ICD9CM|Erythem nodos tb-cult dx|Erythem nodos tb-cult dx
C0152859|T047|AB|017.15|ICD9CM|Erythem nod tb-histo dx|Erythem nod tb-histo dx
C0152860|T047|AB|017.16|ICD9CM|Erythem nod tb-oth test|Erythem nod tb-oth test
C0152861|T047|HT|017.2|ICD9CM|Tuberculosis of peripheral lymph nodes|Tuberculosis of peripheral lymph nodes
C0152861|T047|AB|017.20|ICD9CM|TB periph lymph-unspec|TB periph lymph-unspec
C0152861|T047|PT|017.20|ICD9CM|Tuberculosis of peripheral lymph nodes, unspecified|Tuberculosis of peripheral lymph nodes, unspecified
C0152862|T047|AB|017.21|ICD9CM|TB periph lymph-no exam|TB periph lymph-no exam
C0152862|T047|PT|017.21|ICD9CM|Tuberculosis of peripheral lymph nodes, bacteriological or histological examination not done|Tuberculosis of peripheral lymph nodes, bacteriological or histological examination not done
C0152863|T047|AB|017.22|ICD9CM|TB periph lymph-exam unk|TB periph lymph-exam unk
C0152864|T047|AB|017.23|ICD9CM|TB periph lymph-micro dx|TB periph lymph-micro dx
C0152864|T047|PT|017.23|ICD9CM|Tuberculosis of peripheral lymph nodes, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of peripheral lymph nodes, tubercle bacilli found (in sputum) by microscopy
C0152865|T047|AB|017.24|ICD9CM|TB periph lymph-cult dx|TB periph lymph-cult dx
C0152866|T047|AB|017.25|ICD9CM|TB periph lymph-histo dx|TB periph lymph-histo dx
C0152867|T047|AB|017.26|ICD9CM|TB periph lymph-oth test|TB periph lymph-oth test
C0041322|T047|HT|017.3|ICD9CM|Tuberculosis of eye|Tuberculosis of eye
C0041322|T047|AB|017.30|ICD9CM|TB of eye-unspec|TB of eye-unspec
C0041322|T047|PT|017.30|ICD9CM|Tuberculosis of eye, unspecified|Tuberculosis of eye, unspecified
C0152868|T047|AB|017.31|ICD9CM|TB of eye-no exam|TB of eye-no exam
C0152868|T047|PT|017.31|ICD9CM|Tuberculosis of eye, bacteriological or histological examination not done|Tuberculosis of eye, bacteriological or histological examination not done
C0152869|T047|AB|017.32|ICD9CM|TB of eye-exam unkn|TB of eye-exam unkn
C0152869|T047|PT|017.32|ICD9CM|Tuberculosis of eye, bacteriological or histological examination unknown (at present)|Tuberculosis of eye, bacteriological or histological examination unknown (at present)
C0152870|T047|AB|017.33|ICD9CM|TB of eye-micro dx|TB of eye-micro dx
C0152870|T047|PT|017.33|ICD9CM|Tuberculosis of eye, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of eye, tubercle bacilli found (in sputum) by microscopy
C0152871|T047|AB|017.34|ICD9CM|TB of eye-cult dx|TB of eye-cult dx
C0152872|T047|AB|017.35|ICD9CM|TB of eye-histo dx|TB of eye-histo dx
C0152873|T047|AB|017.36|ICD9CM|TB of eye-oth test|TB of eye-oth test
C0152874|T047|HT|017.4|ICD9CM|Tuberculosis of ear|Tuberculosis of ear
C0374976|T047|AB|017.40|ICD9CM|TB of ear-unspec|TB of ear-unspec
C0374976|T047|PT|017.40|ICD9CM|Tuberculosis of ear, unspecified|Tuberculosis of ear, unspecified
C0152875|T047|AB|017.41|ICD9CM|TB of ear-no exam|TB of ear-no exam
C0152875|T047|PT|017.41|ICD9CM|Tuberculosis of ear, bacteriological or histological examination not done|Tuberculosis of ear, bacteriological or histological examination not done
C0152876|T047|AB|017.42|ICD9CM|TB of ear-exam unkn|TB of ear-exam unkn
C0152876|T047|PT|017.42|ICD9CM|Tuberculosis of ear, bacteriological or histological examination unknown (at present)|Tuberculosis of ear, bacteriological or histological examination unknown (at present)
C0152877|T047|AB|017.43|ICD9CM|TB of ear-micro dx|TB of ear-micro dx
C0152877|T047|PT|017.43|ICD9CM|Tuberculosis of ear, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of ear, tubercle bacilli found (in sputum) by microscopy
C0152878|T047|AB|017.44|ICD9CM|TB of ear-cult dx|TB of ear-cult dx
C0152879|T047|AB|017.45|ICD9CM|TB of ear-histo dx|TB of ear-histo dx
C0152880|T047|AB|017.46|ICD9CM|TB of ear-oth test|TB of ear-oth test
C0152881|T047|HT|017.5|ICD9CM|Tuberculosis of thyroid gland|Tuberculosis of thyroid gland
C0152882|T047|AB|017.50|ICD9CM|TB of thyroid-unspec|TB of thyroid-unspec
C0152882|T047|PT|017.50|ICD9CM|Tuberculosis of thyroid gland, unspecified|Tuberculosis of thyroid gland, unspecified
C0152883|T047|AB|017.51|ICD9CM|TB of thyroid-no exam|TB of thyroid-no exam
C0152883|T047|PT|017.51|ICD9CM|Tuberculosis of thyroid gland, bacteriological or histological examination not done|Tuberculosis of thyroid gland, bacteriological or histological examination not done
C0152884|T047|AB|017.52|ICD9CM|TB of thyroid-exam unkn|TB of thyroid-exam unkn
C0152884|T047|PT|017.52|ICD9CM|Tuberculosis of thyroid gland, bacteriological or histological examination unknown (at present)|Tuberculosis of thyroid gland, bacteriological or histological examination unknown (at present)
C0152885|T047|AB|017.53|ICD9CM|TB of thyroid-micro dx|TB of thyroid-micro dx
C0152885|T047|PT|017.53|ICD9CM|Tuberculosis of thyroid gland, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of thyroid gland, tubercle bacilli found (in sputum) by microscopy
C0152886|T047|AB|017.54|ICD9CM|TB of thyroid-cult dx|TB of thyroid-cult dx
C0152887|T047|AB|017.55|ICD9CM|TB of thyroid-histo dx|TB of thyroid-histo dx
C0152888|T047|AB|017.56|ICD9CM|TB of thyroid-oth test|TB of thyroid-oth test
C0152889|T047|HT|017.6|ICD9CM|Tuberculosis of adrenal glands|Tuberculosis of adrenal glands
C0152889|T047|AB|017.60|ICD9CM|TB of adrenal-unspec|TB of adrenal-unspec
C0152889|T047|PT|017.60|ICD9CM|Tuberculosis of adrenal glands, unspecified|Tuberculosis of adrenal glands, unspecified
C0152890|T047|AB|017.61|ICD9CM|TB of adrenal-no exam|TB of adrenal-no exam
C0152890|T047|PT|017.61|ICD9CM|Tuberculosis of adrenal glands, bacteriological or histological examination not done|Tuberculosis of adrenal glands, bacteriological or histological examination not done
C0152891|T047|AB|017.62|ICD9CM|TB of adrenal-exam unkn|TB of adrenal-exam unkn
C0152891|T047|PT|017.62|ICD9CM|Tuberculosis of adrenal glands, bacteriological or histological examination unknown (at present)|Tuberculosis of adrenal glands, bacteriological or histological examination unknown (at present)
C0152892|T047|AB|017.63|ICD9CM|TB of adrenal-micro dx|TB of adrenal-micro dx
C0152892|T047|PT|017.63|ICD9CM|Tuberculosis of adrenal glands, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of adrenal glands, tubercle bacilli found (in sputum) by microscopy
C0152893|T047|AB|017.64|ICD9CM|TB of adrenal-cult dx|TB of adrenal-cult dx
C0152894|T047|AB|017.65|ICD9CM|TB of adrenal-histo dx|TB of adrenal-histo dx
C0152895|T047|AB|017.66|ICD9CM|TB of adrenal-oth test|TB of adrenal-oth test
C0041331|T047|HT|017.7|ICD9CM|Tuberculosis of spleen|Tuberculosis of spleen
C0374977|T047|AB|017.70|ICD9CM|TB of spleen-unspec|TB of spleen-unspec
C0374977|T047|PT|017.70|ICD9CM|Tuberculosis of spleen, unspecified|Tuberculosis of spleen, unspecified
C0152896|T047|AB|017.71|ICD9CM|TB of spleen-no exam|TB of spleen-no exam
C0152896|T047|PT|017.71|ICD9CM|Tuberculosis of spleen, bacteriological or histological examination not done|Tuberculosis of spleen, bacteriological or histological examination not done
C0152897|T047|AB|017.72|ICD9CM|TB of spleen-exam unkn|TB of spleen-exam unkn
C0152897|T047|PT|017.72|ICD9CM|Tuberculosis of spleen, bacteriological or histological examination unknown (at present)|Tuberculosis of spleen, bacteriological or histological examination unknown (at present)
C0152898|T047|AB|017.73|ICD9CM|TB of spleen-micro dx|TB of spleen-micro dx
C0152898|T047|PT|017.73|ICD9CM|Tuberculosis of spleen, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of spleen, tubercle bacilli found (in sputum) by microscopy
C0152899|T047|AB|017.74|ICD9CM|TB of spleen-cult dx|TB of spleen-cult dx
C0152900|T047|AB|017.75|ICD9CM|TB of spleen-histo dx|TB of spleen-histo dx
C0152901|T047|AB|017.76|ICD9CM|TB of spleen-oth test|TB of spleen-oth test
C0152902|T047|HT|017.8|ICD9CM|Tuberculosis of esophagus|Tuberculosis of esophagus
C0374978|T047|AB|017.80|ICD9CM|TB esophagus-unspec|TB esophagus-unspec
C0374978|T047|PT|017.80|ICD9CM|Tuberculosis of esophagus, unspecified|Tuberculosis of esophagus, unspecified
C0152903|T047|AB|017.81|ICD9CM|TB esophagus-no exam|TB esophagus-no exam
C0152903|T047|PT|017.81|ICD9CM|Tuberculosis of esophagus, bacteriological or histological examination not done|Tuberculosis of esophagus, bacteriological or histological examination not done
C0152904|T047|AB|017.82|ICD9CM|TB esophagus-exam unkn|TB esophagus-exam unkn
C0152904|T047|PT|017.82|ICD9CM|Tuberculosis of esophagus, bacteriological or histological examination unknown (at present)|Tuberculosis of esophagus, bacteriological or histological examination unknown (at present)
C0152905|T047|AB|017.83|ICD9CM|TB esophagus-micro dx|TB esophagus-micro dx
C0152905|T047|PT|017.83|ICD9CM|Tuberculosis of esophagus, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of esophagus, tubercle bacilli found (in sputum) by microscopy
C0152906|T047|AB|017.84|ICD9CM|TB esophagus-cult dx|TB esophagus-cult dx
C0152907|T047|AB|017.85|ICD9CM|TB esophagus-histo dx|TB esophagus-histo dx
C0152908|T047|AB|017.86|ICD9CM|TB esophagus-oth test|TB esophagus-oth test
C0041301|T047|HT|017.9|ICD9CM|Tuberculosis of other specified organs|Tuberculosis of other specified organs
C0041301|T047|AB|017.90|ICD9CM|TB of organ NEC-unspec|TB of organ NEC-unspec
C0041301|T047|PT|017.90|ICD9CM|Tuberculosis of other specified organs, unspecified|Tuberculosis of other specified organs, unspecified
C0152909|T047|AB|017.91|ICD9CM|TB of organ NEC-no exam|TB of organ NEC-no exam
C0152909|T047|PT|017.91|ICD9CM|Tuberculosis of other specified organs, bacteriological or histological examination not done|Tuberculosis of other specified organs, bacteriological or histological examination not done
C0152910|T047|AB|017.92|ICD9CM|TB organ NEC-exam unkn|TB organ NEC-exam unkn
C0152911|T047|AB|017.93|ICD9CM|TB of organ NEC-micro dx|TB of organ NEC-micro dx
C0152911|T047|PT|017.93|ICD9CM|Tuberculosis of other specified organs, tubercle bacilli found (in sputum) by microscopy|Tuberculosis of other specified organs, tubercle bacilli found (in sputum) by microscopy
C0152912|T047|AB|017.94|ICD9CM|TB of organ NEC-cult dx|TB of organ NEC-cult dx
C0152913|T047|AB|017.95|ICD9CM|TB of organ NEC-histo dx|TB of organ NEC-histo dx
C0152914|T047|AB|017.96|ICD9CM|TB of organ NEC-oth test|TB of organ NEC-oth test
C0041321|T047|HT|018|ICD9CM|Miliary tuberculosis|Miliary tuberculosis
C0152915|T047|HT|018.0|ICD9CM|Acute miliary tuberculosis|Acute miliary tuberculosis
C0152915|T047|AB|018.00|ICD9CM|Acute miliary tb-unspec|Acute miliary tb-unspec
C0152915|T047|PT|018.00|ICD9CM|Acute miliary tuberculosis, unspecified|Acute miliary tuberculosis, unspecified
C0152916|T047|AB|018.01|ICD9CM|Acute miliary tb-no exam|Acute miliary tb-no exam
C0152916|T047|PT|018.01|ICD9CM|Acute miliary tuberculosis, bacteriological or histological examination not done|Acute miliary tuberculosis, bacteriological or histological examination not done
C0152917|T047|AB|018.02|ICD9CM|Ac miliary tb-exam unkn|Ac miliary tb-exam unkn
C0152917|T047|PT|018.02|ICD9CM|Acute miliary tuberculosis, bacteriological or histological examination unknown (at present)|Acute miliary tuberculosis, bacteriological or histological examination unknown (at present)
C0152918|T047|AB|018.03|ICD9CM|Ac miliary tb-micro dx|Ac miliary tb-micro dx
C0152918|T047|PT|018.03|ICD9CM|Acute miliary tuberculosis, tubercle bacilli found (in sputum) by microscopy|Acute miliary tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152919|T047|AB|018.04|ICD9CM|Acute miliary tb-cult dx|Acute miliary tb-cult dx
C0152920|T047|AB|018.05|ICD9CM|Ac miliary tb-histo dx|Ac miliary tb-histo dx
C0152921|T047|AB|018.06|ICD9CM|Ac miliary tb-oth test|Ac miliary tb-oth test
C0152922|T047|HT|018.8|ICD9CM|Other specified miliary tuberculosis|Other specified miliary tuberculosis
C0152922|T047|AB|018.80|ICD9CM|Miliary TB NEC-unspec|Miliary TB NEC-unspec
C0152922|T047|PT|018.80|ICD9CM|Other specified miliary tuberculosis, unspecified|Other specified miliary tuberculosis, unspecified
C0152923|T047|AB|018.81|ICD9CM|Miliary TB NEC-no exam|Miliary TB NEC-no exam
C0152923|T047|PT|018.81|ICD9CM|Other specified miliary tuberculosis, bacteriological or histological examination not done|Other specified miliary tuberculosis, bacteriological or histological examination not done
C0152924|T047|AB|018.82|ICD9CM|Miliary TB NEC-exam unkn|Miliary TB NEC-exam unkn
C0152925|T047|AB|018.83|ICD9CM|Miliary TB NEC-micro dx|Miliary TB NEC-micro dx
C0152925|T047|PT|018.83|ICD9CM|Other specified miliary tuberculosis, tubercle bacilli found (in sputum) by microscopy|Other specified miliary tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152926|T047|AB|018.84|ICD9CM|Miliary TB NEC-cult dx|Miliary TB NEC-cult dx
C0152927|T047|AB|018.85|ICD9CM|Miliary TB NEC-histo dx|Miliary TB NEC-histo dx
C0152928|T047|AB|018.86|ICD9CM|Miliary TB NEC-oth test|Miliary TB NEC-oth test
C0041321|T047|HT|018.9|ICD9CM|Unspecified miliary tuberculosis|Unspecified miliary tuberculosis
C0041321|T047|AB|018.90|ICD9CM|Miliary TB NOS-unspec|Miliary TB NOS-unspec
C0041321|T047|PT|018.90|ICD9CM|Miliary tuberculosis, unspecified, unspecified|Miliary tuberculosis, unspecified, unspecified
C0152929|T047|AB|018.91|ICD9CM|Miliary TB NOS-no exam|Miliary TB NOS-no exam
C0152929|T047|PT|018.91|ICD9CM|Miliary tuberculosis, unspecified, bacteriological or histological examination not done|Miliary tuberculosis, unspecified, bacteriological or histological examination not done
C0152930|T047|AB|018.92|ICD9CM|Miliary TB NOS-exam unkn|Miliary TB NOS-exam unkn
C0152930|T047|PT|018.92|ICD9CM|Miliary tuberculosis, unspecified, bacteriological or histological examination unknown (at present)|Miliary tuberculosis, unspecified, bacteriological or histological examination unknown (at present)
C0152931|T047|AB|018.93|ICD9CM|Miliary TB NOS-micro dx|Miliary TB NOS-micro dx
C0152931|T047|PT|018.93|ICD9CM|Miliary tuberculosis, unspecified, tubercle bacilli found (in sputum) by microscopy|Miliary tuberculosis, unspecified, tubercle bacilli found (in sputum) by microscopy
C0152932|T047|AB|018.94|ICD9CM|Miliary TB NOS-cult dx|Miliary TB NOS-cult dx
C0152933|T047|AB|018.95|ICD9CM|Miliary TB NOS-histo dx|Miliary TB NOS-histo dx
C0152934|T047|AB|018.96|ICD9CM|Miliary TB NOS-oth test|Miliary TB NOS-oth test
C0032064|T047|HT|020|ICD9CM|Plague|Plague
C0311376|T047|HT|020-027.99|ICD9CM|ZOONOTIC BACTERIAL DISEASES|ZOONOTIC BACTERIAL DISEASES
C0282312|T047|AB|020.0|ICD9CM|Bubonic plague|Bubonic plague
C0282312|T047|PT|020.0|ICD9CM|Bubonic plague|Bubonic plague
C0152935|T047|AB|020.1|ICD9CM|Cellulocutaneous plague|Cellulocutaneous plague
C0152935|T047|PT|020.1|ICD9CM|Cellulocutaneous plague|Cellulocutaneous plague
C0152936|T047|AB|020.2|ICD9CM|Septicemic plague|Septicemic plague
C0152936|T047|PT|020.2|ICD9CM|Septicemic plague|Septicemic plague
C0152937|T047|AB|020.3|ICD9CM|Primary pneumonic plague|Primary pneumonic plague
C0152937|T047|PT|020.3|ICD9CM|Primary pneumonic plague|Primary pneumonic plague
C0152938|T047|AB|020.4|ICD9CM|Secondary pneumon plague|Secondary pneumon plague
C0152938|T047|PT|020.4|ICD9CM|Secondary pneumonic plague|Secondary pneumonic plague
C0524688|T047|AB|020.5|ICD9CM|Pneumonic plague NOS|Pneumonic plague NOS
C0524688|T047|PT|020.5|ICD9CM|Pneumonic plague, unspecified|Pneumonic plague, unspecified
C0152940|T047|PT|020.8|ICD9CM|Other specified types of plague|Other specified types of plague
C0152940|T047|AB|020.8|ICD9CM|Other types of plague|Other types of plague
C0032064|T047|AB|020.9|ICD9CM|Plague NOS|Plague NOS
C0032064|T047|PT|020.9|ICD9CM|Plague, unspecified|Plague, unspecified
C0041351|T047|HT|021|ICD9CM|Tularemia|Tularemia
C0152941|T047|AB|021.0|ICD9CM|Ulceroglandul tularemia|Ulceroglandul tularemia
C0152941|T047|PT|021.0|ICD9CM|Ulceroglandular tularemia|Ulceroglandular tularemia
C0152942|T047|AB|021.1|ICD9CM|Enteric tularemia|Enteric tularemia
C0152942|T047|PT|021.1|ICD9CM|Enteric tularemia|Enteric tularemia
C0339946|T047|AB|021.2|ICD9CM|Pulmonary tularemia|Pulmonary tularemia
C0339946|T047|PT|021.2|ICD9CM|Pulmonary tularemia|Pulmonary tularemia
C0152944|T047|AB|021.3|ICD9CM|Oculoglandular tularemia|Oculoglandular tularemia
C0152944|T047|PT|021.3|ICD9CM|Oculoglandular tularemia|Oculoglandular tularemia
C0029835|T047|PT|021.8|ICD9CM|Other specified tularemia|Other specified tularemia
C0029835|T047|AB|021.8|ICD9CM|Tularemia NEC|Tularemia NEC
C0041351|T047|AB|021.9|ICD9CM|Tularemia NOS|Tularemia NOS
C0041351|T047|PT|021.9|ICD9CM|Unspecified tularemia|Unspecified tularemia
C0003175|T047|HT|022|ICD9CM|Anthrax|Anthrax
C0003177|T047|AB|022.0|ICD9CM|Cutaneous anthrax|Cutaneous anthrax
C0003177|T047|PT|022.0|ICD9CM|Cutaneous anthrax|Cutaneous anthrax
C0155866|T047|AB|022.1|ICD9CM|Pulmonary anthrax|Pulmonary anthrax
C0155866|T047|PT|022.1|ICD9CM|Pulmonary anthrax|Pulmonary anthrax
C0152945|T047|AB|022.2|ICD9CM|Gastrointestinal anthrax|Gastrointestinal anthrax
C0152945|T047|PT|022.2|ICD9CM|Gastrointestinal anthrax|Gastrointestinal anthrax
C0152946|T047|AB|022.3|ICD9CM|Anthrax septicemia|Anthrax septicemia
C0152946|T047|PT|022.3|ICD9CM|Anthrax septicemia|Anthrax septicemia
C0152947|T047|AB|022.8|ICD9CM|Other anthrax manifest|Other anthrax manifest
C0152947|T047|PT|022.8|ICD9CM|Other specified manifestations of anthrax|Other specified manifestations of anthrax
C0003175|T047|AB|022.9|ICD9CM|Anthrax NOS|Anthrax NOS
C0003175|T047|PT|022.9|ICD9CM|Anthrax, unspecified|Anthrax, unspecified
C0006309|T047|HT|023|ICD9CM|Brucellosis|Brucellosis
C0302362|T047|AB|023.0|ICD9CM|Brucella melitensis|Brucella melitensis
C0302362|T047|PT|023.0|ICD9CM|Brucella melitensis|Brucella melitensis
C0302363|T047|AB|023.1|ICD9CM|Brucella abortus|Brucella abortus
C0302363|T047|PT|023.1|ICD9CM|Brucella abortus|Brucella abortus
C0275594|T047|AB|023.2|ICD9CM|Brucella suis|Brucella suis
C0275594|T047|PT|023.2|ICD9CM|Brucella suis|Brucella suis
C0494040|T047|AB|023.3|ICD9CM|Brucella canis|Brucella canis
C0494040|T047|PT|023.3|ICD9CM|Brucella canis|Brucella canis
C0029527|T047|AB|023.8|ICD9CM|Brucellosis NEC|Brucellosis NEC
C0029527|T047|PT|023.8|ICD9CM|Other brucellosis|Other brucellosis
C0006309|T047|AB|023.9|ICD9CM|Brucellosis NOS|Brucellosis NOS
C0006309|T047|PT|023.9|ICD9CM|Brucellosis, unspecified|Brucellosis, unspecified
C0017589|T047|AB|024|ICD9CM|Glanders|Glanders
C0017589|T047|PT|024|ICD9CM|Glanders|Glanders
C0025229|T047|AB|025|ICD9CM|Melioidosis|Melioidosis
C0025229|T047|PT|025|ICD9CM|Melioidosis|Melioidosis
C0034686|T047|HT|026|ICD9CM|Rat-bite fever|Rat-bite fever
C0152062|T047|AB|026.0|ICD9CM|Spirillary fever|Spirillary fever
C0152062|T047|PT|026.0|ICD9CM|Spirillary fever|Spirillary fever
C0152063|T047|AB|026.1|ICD9CM|Streptobacillary fever|Streptobacillary fever
C0152063|T047|PT|026.1|ICD9CM|Streptobacillary fever|Streptobacillary fever
C0034686|T047|AB|026.9|ICD9CM|Rat-bite fever NOS|Rat-bite fever NOS
C0034686|T047|PT|026.9|ICD9CM|Unspecified rat-bite fever|Unspecified rat-bite fever
C0152948|T047|HT|027|ICD9CM|Other zoonotic bacterial diseases|Other zoonotic bacterial diseases
C0023860|T047|AB|027.0|ICD9CM|Listeriosis|Listeriosis
C0023860|T047|PT|027.0|ICD9CM|Listeriosis|Listeriosis
C0014736|T047|AB|027.1|ICD9CM|Erysipelothrix infection|Erysipelothrix infection
C0014736|T047|PT|027.1|ICD9CM|Erysipelothrix infection|Erysipelothrix infection
C0030636|T047|AB|027.2|ICD9CM|Pasteurellosis|Pasteurellosis
C0030636|T047|PT|027.2|ICD9CM|Pasteurellosis|Pasteurellosis
C0152949|T047|PT|027.8|ICD9CM|Other specified zoonotic bacterial diseases|Other specified zoonotic bacterial diseases
C0152949|T047|AB|027.8|ICD9CM|Zoonotic bact dis NEC|Zoonotic bact dis NEC
C0311376|T047|PT|027.9|ICD9CM|Unspecified zoonotic bacterial disease|Unspecified zoonotic bacterial disease
C0311376|T047|AB|027.9|ICD9CM|Zoonotic bact dis NOS|Zoonotic bact dis NOS
C0023343|T047|HT|030|ICD9CM|Leprosy|Leprosy
C2939130|T047|HT|030-041.99|ICD9CM|OTHER BACTERIAL DISEASES|OTHER BACTERIAL DISEASES
C0023348|T047|AB|030.0|ICD9CM|Lepromatous leprosy|Lepromatous leprosy
C0023348|T047|PT|030.0|ICD9CM|Lepromatous leprosy [type L]|Lepromatous leprosy [type L]
C0023351|T047|AB|030.1|ICD9CM|Tuberculoid leprosy|Tuberculoid leprosy
C0023351|T047|PT|030.1|ICD9CM|Tuberculoid leprosy [type T]|Tuberculoid leprosy [type T]
C0021192|T047|AB|030.2|ICD9CM|Indeterminate leprosy|Indeterminate leprosy
C0021192|T047|PT|030.2|ICD9CM|Indeterminate leprosy [group I]|Indeterminate leprosy [group I]
C0023346|T047|AB|030.3|ICD9CM|Borderline leprosy|Borderline leprosy
C0023346|T047|PT|030.3|ICD9CM|Borderline leprosy [group B]|Borderline leprosy [group B]
C0029811|T047|AB|030.8|ICD9CM|Leprosy NEC|Leprosy NEC
C0029811|T047|PT|030.8|ICD9CM|Other specified leprosy|Other specified leprosy
C0023343|T047|AB|030.9|ICD9CM|Leprosy NOS|Leprosy NOS
C0023343|T047|PT|030.9|ICD9CM|Leprosy, unspecified|Leprosy, unspecified
C0152950|T047|HT|031|ICD9CM|Diseases due to other mycobacteria|Diseases due to other mycobacteria
C0392054|T047|PT|031.0|ICD9CM|Pulmonary diseases due to other mycobacteria|Pulmonary diseases due to other mycobacteria
C0392054|T047|AB|031.0|ICD9CM|Pulmonary mycobacteria|Pulmonary mycobacteria
C0010487|T047|PT|031.1|ICD9CM|Cutaneous diseases due to other mycobacteria|Cutaneous diseases due to other mycobacteria
C0010487|T047|AB|031.1|ICD9CM|Cutaneous mycobacteria|Cutaneous mycobacteria
C0489980|T047|PT|031.2|ICD9CM|Disseminated due to other mycobacteria|Disseminated due to other mycobacteria
C0489980|T047|AB|031.2|ICD9CM|DMAC bacteremia|DMAC bacteremia
C0152951|T047|AB|031.8|ICD9CM|Mycobacterial dis NEC|Mycobacterial dis NEC
C0152951|T047|PT|031.8|ICD9CM|Other specified mycobacterial diseases|Other specified mycobacterial diseases
C0026918|T047|AB|031.9|ICD9CM|Mycobacterial dis NOS|Mycobacterial dis NOS
C0026918|T047|PT|031.9|ICD9CM|Unspecified diseases due to mycobacteria|Unspecified diseases due to mycobacteria
C0012546|T047|HT|032|ICD9CM|Diphtheria|Diphtheria
C0012556|T047|AB|032.0|ICD9CM|Faucial diphtheria|Faucial diphtheria
C0012556|T047|PT|032.0|ICD9CM|Faucial diphtheria|Faucial diphtheria
C0012558|T047|PT|032.1|ICD9CM|Nasopharyngeal diphtheria|Nasopharyngeal diphtheria
C0012558|T047|AB|032.1|ICD9CM|Nasopharynx diphtheria|Nasopharynx diphtheria
C0012553|T047|AB|032.2|ICD9CM|Ant nasal diphtheria|Ant nasal diphtheria
C0012553|T047|PT|032.2|ICD9CM|Anterior nasal diphtheria|Anterior nasal diphtheria
C0012557|T047|AB|032.3|ICD9CM|Laryngeal diphtheria|Laryngeal diphtheria
C0012557|T047|PT|032.3|ICD9CM|Laryngeal diphtheria|Laryngeal diphtheria
C0029764|T047|HT|032.8|ICD9CM|Other specified diphtheria|Other specified diphtheria
C0012554|T047|AB|032.81|ICD9CM|Conjunctival diphtheria|Conjunctival diphtheria
C0012554|T047|PT|032.81|ICD9CM|Conjunctival diphtheria|Conjunctival diphtheria
C0152952|T047|AB|032.82|ICD9CM|Diphtheritic myocarditis|Diphtheritic myocarditis
C0152952|T047|PT|032.82|ICD9CM|Diphtheritic myocarditis|Diphtheritic myocarditis
C0152953|T047|AB|032.83|ICD9CM|Diphtheritic peritonitis|Diphtheritic peritonitis
C0152953|T047|PT|032.83|ICD9CM|Diphtheritic peritonitis|Diphtheritic peritonitis
C0152954|T047|AB|032.84|ICD9CM|Diphtheritic cystitis|Diphtheritic cystitis
C0152954|T047|PT|032.84|ICD9CM|Diphtheritic cystitis|Diphtheritic cystitis
C0012555|T047|AB|032.85|ICD9CM|Cutaneous diphtheria|Cutaneous diphtheria
C0012555|T047|PT|032.85|ICD9CM|Cutaneous diphtheria|Cutaneous diphtheria
C0029764|T047|AB|032.89|ICD9CM|Diphtheria NEC|Diphtheria NEC
C0029764|T047|PT|032.89|ICD9CM|Other specified diphtheria|Other specified diphtheria
C0012546|T047|AB|032.9|ICD9CM|Diphtheria NOS|Diphtheria NOS
C0012546|T047|PT|032.9|ICD9CM|Diphtheria, unspecified|Diphtheria, unspecified
C0043168|T047|HT|033|ICD9CM|Whooping cough|Whooping cough
C0043167|T047|AB|033.0|ICD9CM|Bordetella pertussis|Bordetella pertussis
C0043167|T047|PT|033.0|ICD9CM|Whooping cough due to bordetella pertussis [B. pertussis]|Whooping cough due to bordetella pertussis [B. pertussis]
C0275742|T047|AB|033.1|ICD9CM|Bordetella parapertussis|Bordetella parapertussis
C0275742|T047|PT|033.1|ICD9CM|Whooping cough due to bordetella parapertussis [B. parapertussis]|Whooping cough due to bordetella parapertussis [B. parapertussis]
C0043170|T047|PT|033.8|ICD9CM|Whooping cough due to other specified organism|Whooping cough due to other specified organism
C0043170|T047|AB|033.8|ICD9CM|Whooping cough NEC|Whooping cough NEC
C0043168|T047|AB|033.9|ICD9CM|Whooping cough NOS|Whooping cough NOS
C0043168|T047|PT|033.9|ICD9CM|Whooping cough, unspecified organism|Whooping cough, unspecified organism
C0343487|T047|HT|034|ICD9CM|Streptococcal sore throat and scarlet fever|Streptococcal sore throat and scarlet fever
C0036689|T047|AB|034.0|ICD9CM|Strep sore throat|Strep sore throat
C0036689|T047|PT|034.0|ICD9CM|Streptococcal sore throat|Streptococcal sore throat
C0036285|T047|AB|034.1|ICD9CM|Scarlet fever|Scarlet fever
C0036285|T047|PT|034.1|ICD9CM|Scarlet fever|Scarlet fever
C0014733|T047|AB|035|ICD9CM|Erysipelas|Erysipelas
C0014733|T047|PT|035|ICD9CM|Erysipelas|Erysipelas
C0025303|T047|HT|036|ICD9CM|Meningococcal infection|Meningococcal infection
C0025294|T047|AB|036.0|ICD9CM|Meningococcal meningitis|Meningococcal meningitis
C0025294|T047|PT|036.0|ICD9CM|Meningococcal meningitis|Meningococcal meningitis
C0152957|T047|AB|036.1|ICD9CM|Meningococc encephalitis|Meningococc encephalitis
C0152957|T047|PT|036.1|ICD9CM|Meningococcal encephalitis|Meningococcal encephalitis
C0025306|T047|AB|036.2|ICD9CM|Meningococcemia|Meningococcemia
C0025306|T047|PT|036.2|ICD9CM|Meningococcemia|Meningococcemia
C1403891|T047|AB|036.3|ICD9CM|Meningococc adrenal synd|Meningococc adrenal synd
C1403891|T047|PT|036.3|ICD9CM|Waterhouse-Friderichsen syndrome, meningococcal|Waterhouse-Friderichsen syndrome, meningococcal
C0152958|T047|HT|036.4|ICD9CM|Meningococcal carditis|Meningococcal carditis
C0152958|T047|AB|036.40|ICD9CM|Meningococc carditis NOS|Meningococc carditis NOS
C0152958|T047|PT|036.40|ICD9CM|Meningococcal carditis, unspecified|Meningococcal carditis, unspecified
C0152959|T047|AB|036.41|ICD9CM|Meningococc pericarditis|Meningococc pericarditis
C0152959|T047|PT|036.41|ICD9CM|Meningococcal pericarditis|Meningococcal pericarditis
C0152960|T047|AB|036.42|ICD9CM|Meningococc endocarditis|Meningococc endocarditis
C0152960|T047|PT|036.42|ICD9CM|Meningococcal endocarditis|Meningococcal endocarditis
C0152961|T047|AB|036.43|ICD9CM|Meningococc myocarditis|Meningococc myocarditis
C0152961|T047|PT|036.43|ICD9CM|Meningococcal myocarditis|Meningococcal myocarditis
C0029815|T047|HT|036.8|ICD9CM|Other specified meningococcal infections|Other specified meningococcal infections
C0152962|T047|AB|036.81|ICD9CM|Meningococc optic neurit|Meningococc optic neurit
C0152962|T047|PT|036.81|ICD9CM|Meningococcal optic neuritis|Meningococcal optic neuritis
C0238009|T047|AB|036.82|ICD9CM|Meningococc arthropathy|Meningococc arthropathy
C0238009|T047|PT|036.82|ICD9CM|Meningococcal arthropathy|Meningococcal arthropathy
C0029815|T047|AB|036.89|ICD9CM|Meningococcal infect NEC|Meningococcal infect NEC
C0029815|T047|PT|036.89|ICD9CM|Other specified meningococcal infections|Other specified meningococcal infections
C0025303|T047|AB|036.9|ICD9CM|Meningococcal infect NOS|Meningococcal infect NOS
C0025303|T047|PT|036.9|ICD9CM|Meningococcal infection, unspecified|Meningococcal infection, unspecified
C0039614|T047|AB|037|ICD9CM|Tetanus|Tetanus
C0039614|T047|PT|037|ICD9CM|Tetanus|Tetanus
C0036690|T047|HT|038|ICD9CM|Septicemia|Septicemia
C0152964|T047|AB|038.0|ICD9CM|Streptococcal septicemia|Streptococcal septicemia
C0152964|T047|PT|038.0|ICD9CM|Streptococcal septicemia|Streptococcal septicemia
C0152965|T047|HT|038.1|ICD9CM|Staphylococcal septicemia|Staphylococcal septicemia
C0152965|T047|AB|038.10|ICD9CM|Staphylcocc septicem NOS|Staphylcocc septicem NOS
C0152965|T047|PT|038.10|ICD9CM|Staphylococcal septicemia, unspecified|Staphylococcal septicemia, unspecified
C2349736|T047|AB|038.11|ICD9CM|Meth susc Staph aur sept|Meth susc Staph aur sept
C2349736|T047|PT|038.11|ICD9CM|Methicillin susceptible Staphylococcus aureus septicemia|Methicillin susceptible Staphylococcus aureus septicemia
C0877176|T047|PT|038.12|ICD9CM|Methicillin resistant Staphylococcus aureus septicemia|Methicillin resistant Staphylococcus aureus septicemia
C0877176|T047|AB|038.12|ICD9CM|MRSA septicemia|MRSA septicemia
C0489981|T047|PT|038.19|ICD9CM|Other staphylococcal septicemia|Other staphylococcal septicemia
C0489981|T047|AB|038.19|ICD9CM|Staphylcocc septicem NEC|Staphylcocc septicem NEC
C0152966|T047|AB|038.2|ICD9CM|Pneumococcal septicemia|Pneumococcal septicemia
C0152966|T047|PT|038.2|ICD9CM|Pneumococcal septicemia [Streptococcus pneumoniae septicemia]|Pneumococcal septicemia [Streptococcus pneumoniae septicemia]
C0152967|T047|AB|038.3|ICD9CM|Anaerobic septicemia|Anaerobic septicemia
C0152967|T047|PT|038.3|ICD9CM|Septicemia due to anaerobes|Septicemia due to anaerobes
C0276063|T047|HT|038.4|ICD9CM|Septicemia due to other gram-negative organisms|Septicemia due to other gram-negative organisms
C0036685|T047|AB|038.40|ICD9CM|Gram-neg septicemia NOS|Gram-neg septicemia NOS
C0036685|T047|PT|038.40|ICD9CM|Septicemia due to gram-negative organism, unspecified|Septicemia due to gram-negative organism, unspecified
C0276029|T047|AB|038.41|ICD9CM|H. influenae septicemia|H. influenae septicemia
C0276029|T047|PT|038.41|ICD9CM|Septicemia due to hemophilus influenzae [H. influenzae]|Septicemia due to hemophilus influenzae [H. influenzae]
C0276088|T047|AB|038.42|ICD9CM|E coli septicemia|E coli septicemia
C0276088|T047|PT|038.42|ICD9CM|Septicemia due to escherichia coli [E. coli]|Septicemia due to escherichia coli [E. coli]
C0152972|T047|AB|038.43|ICD9CM|Pseudomonas septicemia|Pseudomonas septicemia
C0152972|T047|PT|038.43|ICD9CM|Septicemia due to pseudomonas|Septicemia due to pseudomonas
C0152973|T047|PT|038.44|ICD9CM|Septicemia due to serratia|Septicemia due to serratia
C0152973|T047|AB|038.44|ICD9CM|Serratia septicemia|Serratia septicemia
C0276063|T047|AB|038.49|ICD9CM|Gram-neg septicemia NEC|Gram-neg septicemia NEC
C0276063|T047|PT|038.49|ICD9CM|Other septicemia due to gram-negative organisms|Other septicemia due to gram-negative organisms
C0348133|T047|PT|038.8|ICD9CM|Other specified septicemias|Other specified septicemias
C0348133|T047|AB|038.8|ICD9CM|Septicemia NEC|Septicemia NEC
C0036690|T047|AB|038.9|ICD9CM|Septicemia NOS|Septicemia NOS
C0036690|T047|PT|038.9|ICD9CM|Unspecified septicemia|Unspecified septicemia
C0001261|T047|HT|039|ICD9CM|Actinomycotic infections|Actinomycotic infections
C0275567|T047|AB|039.0|ICD9CM|Cutaneous actinomycosis|Cutaneous actinomycosis
C0275567|T047|PT|039.0|ICD9CM|Cutaneous actinomycotic infection|Cutaneous actinomycotic infection
C0275566|T047|AB|039.1|ICD9CM|Pulmonary actinomycosis|Pulmonary actinomycosis
C0275566|T047|PT|039.1|ICD9CM|Pulmonary actinomycotic infection|Pulmonary actinomycotic infection
C0001263|T047|AB|039.2|ICD9CM|Abdominal actinomycosis|Abdominal actinomycosis
C0001263|T047|PT|039.2|ICD9CM|Abdominal actinomycotic infection|Abdominal actinomycotic infection
C0001264|T047|AB|039.3|ICD9CM|Cervicofac actinomycosis|Cervicofac actinomycosis
C0001264|T047|PT|039.3|ICD9CM|Cervicofacial actinomycotic infection|Cervicofacial actinomycotic infection
C2355609|T047|AB|039.4|ICD9CM|Madura foot|Madura foot
C2355609|T047|PT|039.4|ICD9CM|Madura foot|Madura foot
C0001265|T047|AB|039.8|ICD9CM|Actinomycosis NEC|Actinomycosis NEC
C0001265|T047|PT|039.8|ICD9CM|Actinomycotic infection of other specified sites|Actinomycotic infection of other specified sites
C0001261|T047|AB|039.9|ICD9CM|Actinomycosis NOS|Actinomycosis NOS
C0001261|T047|PT|039.9|ICD9CM|Actinomycotic infection of unspecified site|Actinomycotic infection of unspecified site
C2939130|T047|HT|040|ICD9CM|Other bacterial diseases|Other bacterial diseases
C0017105|T047|AB|040.0|ICD9CM|Gas gangrene|Gas gangrene
C0017105|T047|PT|040.0|ICD9CM|Gas gangrene|Gas gangrene
C0035468|T047|AB|040.1|ICD9CM|Rhinoscleroma|Rhinoscleroma
C0035468|T047|PT|040.1|ICD9CM|Rhinoscleroma|Rhinoscleroma
C0023788|T047|AB|040.2|ICD9CM|Whipple's disease|Whipple's disease
C0023788|T047|PT|040.2|ICD9CM|Whipple's disease|Whipple's disease
C0027537|T047|AB|040.3|ICD9CM|Necrobacillosis|Necrobacillosis
C0027537|T047|PT|040.3|ICD9CM|Necrobacillosis|Necrobacillosis
C1955553|T047|HT|040.4|ICD9CM|Other specified botulism|Other specified botulism
C0238027|T047|PT|040.41|ICD9CM|Infant botulism|Infant botulism
C0238027|T047|AB|040.41|ICD9CM|Infant botulism|Infant botulism
C1306794|T047|PT|040.42|ICD9CM|Wound botulism|Wound botulism
C1306794|T047|AB|040.42|ICD9CM|Wound botulism|Wound botulism
C0152977|T047|HT|040.8|ICD9CM|Other specified bacterial disease|Other specified bacterial disease
C0041188|T047|AB|040.81|ICD9CM|Tropical pyomyositis|Tropical pyomyositis
C0041188|T047|PT|040.81|ICD9CM|Tropical pyomyositis|Tropical pyomyositis
C0600327|T047|AB|040.82|ICD9CM|Toxic shock syndrome|Toxic shock syndrome
C0600327|T047|PT|040.82|ICD9CM|Toxic shock syndrome|Toxic shock syndrome
C0152977|T047|AB|040.89|ICD9CM|Bacterial diseases NEC|Bacterial diseases NEC
C0152977|T047|PT|040.89|ICD9CM|Other specified bacterial diseases|Other specified bacterial diseases
C0004622|T047|HT|041|ICD9CM|Bacterial infection in conditions classified elsewhere and of unspecified site|Bacterial infection in conditions classified elsewhere and of unspecified site
C0374982|T047|HT|041.0|ICD9CM|Streptococcus infection in conditions classified elsewhere and of unspecified site|Streptococcus infection in conditions classified elsewhere and of unspecified site
C0374982|T047|AB|041.00|ICD9CM|Streptococcus unspecf|Streptococcus unspecf
C0374983|T047|AB|041.01|ICD9CM|Streptococcus group a|Streptococcus group a
C0374984|T047|AB|041.02|ICD9CM|Streptococcus group b|Streptococcus group b
C0374985|T047|AB|041.03|ICD9CM|Streptococcus group c|Streptococcus group c
C0490039|T047|AB|041.04|ICD9CM|Enterococcus group d|Enterococcus group d
C0374987|T047|AB|041.05|ICD9CM|Streptococcus group g|Streptococcus group g
C0374988|T047|AB|041.09|ICD9CM|Other streptococcus|Other streptococcus
C0374989|T047|HT|041.1|ICD9CM|Staphylococcus infection in conditions classified elsewhere and of unspecified site|Staphylococcus infection in conditions classified elsewhere and of unspecified site
C0374989|T047|AB|041.10|ICD9CM|Staphylococcus unspcfied|Staphylococcus unspcfied
C0374990|T047|AB|041.11|ICD9CM|Mth sus Stph aur els/NOS|Mth sus Stph aur els/NOS
C2349738|T047|AB|041.12|ICD9CM|MRSA elsewhere/NOS|MRSA elsewhere/NOS
C0374991|T047|AB|041.19|ICD9CM|Other staphylococcus|Other staphylococcus
C0032272|T047|AB|041.2|ICD9CM|Pneumococcus infect NOS|Pneumococcus infect NOS
C0032272|T047|PT|041.2|ICD9CM|Pneumococcus infection in conditions classified elsewhere and of unspecified site|Pneumococcus infection in conditions classified elsewhere and of unspecified site
C2712605|T047|PT|041.3|ICD9CM|Friedländer's bacillus infection in conditions classified elsewhere and of unspecified site|Friedländer's bacillus infection in conditions classified elsewhere and of unspecified site
C2712605|T047|AB|041.3|ICD9CM|Klebsiella pneumoniae|Klebsiella pneumoniae
C0014835|T047|HT|041.4|ICD9CM|Escherichia coli [E. coli] infection in conditions classified elsewhere and of unspecified site|Escherichia coli [E. coli] infection in conditions classified elsewhere and of unspecified site
C3161036|T047|PT|041.41|ICD9CM|Shiga toxin-producing Escherichia coli [E. coli] (STEC) O157|Shiga toxin-producing Escherichia coli [E. coli] (STEC) O157
C3161036|T047|AB|041.41|ICD9CM|Shiga txn-produce E.coli|Shiga txn-produce E.coli
C3161167|T047|PT|041.42|ICD9CM|Other specified Shiga toxin-producing Escherichia coli [E. coli] (STEC)|Other specified Shiga toxin-producing Escherichia coli [E. coli] (STEC)
C3161167|T047|AB|041.42|ICD9CM|Shga txn prod E.coli NEC|Shga txn prod E.coli NEC
C3161170|T047|AB|041.43|ICD9CM|Shga txn prod E.coli NOS|Shga txn prod E.coli NOS
C3161170|T047|PT|041.43|ICD9CM|Shiga toxin-producing Escherichia coli [E. coli] (STEC), unspecified|Shiga toxin-producing Escherichia coli [E. coli] (STEC), unspecified
C0014836|T047|AB|041.49|ICD9CM|E.coli infection NEC/NOS|E.coli infection NEC/NOS
C0014836|T047|PT|041.49|ICD9CM|Other and unspecified Escherichia coli [E. coli]|Other and unspecified Escherichia coli [E. coli]
C0019073|T047|AB|041.5|ICD9CM|H. influenzae infect NOS|H. influenzae infect NOS
C0033698|T047|PT|041.6|ICD9CM|Proteus (mirabilis) (morganii) infection in conditions classified elsewhere and of unspecified site|Proteus (mirabilis) (morganii) infection in conditions classified elsewhere and of unspecified site
C0033698|T047|AB|041.6|ICD9CM|Proteus infection NOS|Proteus infection NOS
C0033816|T047|AB|041.7|ICD9CM|Pseudomonas infect NOS|Pseudomonas infect NOS
C0033816|T047|PT|041.7|ICD9CM|Pseudomonas infection in conditions classified elsewhere and of unspecified site|Pseudomonas infection in conditions classified elsewhere and of unspecified site
C0029748|T047|HT|041.8|ICD9CM|Other specified bacterial infections in conditions classified elsewhere and of unspecified site|Other specified bacterial infections in conditions classified elsewhere and of unspecified site
C0374992|T047|AB|041.81|ICD9CM|Mycoplasma|Mycoplasma
C1456246|T047|AB|041.82|ICD9CM|Bacteroides fragilis|Bacteroides fragilis
C1456246|T047|PT|041.82|ICD9CM|Bacteroides fragilis|Bacteroides fragilis
C0374994|T047|AB|041.83|ICD9CM|Clostridium perfringens|Clostridium perfringens
C0374995|T047|AB|041.84|ICD9CM|Other anaerobes|Other anaerobes
C0374996|T047|AB|041.85|ICD9CM|Oth gram negatv bacteria|Oth gram negatv bacteria
C0374997|T047|AB|041.86|ICD9CM|Helicobacter pylori|Helicobacter pylori
C0374997|T047|PT|041.86|ICD9CM|Helicobacter pylori [H. pylori]|Helicobacter pylori [H. pylori]
C0029748|T047|AB|041.89|ICD9CM|Oth specf bacteria|Oth specf bacteria
C0004622|T047|AB|041.9|ICD9CM|Bacterial infection NOS|Bacterial infection NOS
C0004622|T047|PT|041.9|ICD9CM|Bacterial infection, unspecified, in conditions classified elsewhere and of unspecified site|Bacterial infection, unspecified, in conditions classified elsewhere and of unspecified site
C0019693|T047|AB|042|ICD9CM|Human immuno virus dis|Human immuno virus dis
C0019693|T047|PT|042|ICD9CM|Human immunodeficiency virus [HIV] disease|Human immunodeficiency virus [HIV] disease
C0019693|T047|HT|042-042.99|ICD9CM|HUMAN IMMUNODEFICIENCY VIRUS [HIV] INFECTION|HUMAN IMMUNODEFICIENCY VIRUS [HIV] INFECTION
C0032371|T047|HT|045|ICD9CM|Acute poliomyelitis|Acute poliomyelitis
C0032372|T047|HT|045.0|ICD9CM|Acute paralytic poliomyelitis specified as bulbar|Acute paralytic poliomyelitis specified as bulbar
C0152989|T047|AB|045.00|ICD9CM|Ac bulbar polio-type NOS|Ac bulbar polio-type NOS
C0152989|T047|PT|045.00|ICD9CM|Acute paralytic poliomyelitis specified as bulbar, poliovirus, unspecified type|Acute paralytic poliomyelitis specified as bulbar, poliovirus, unspecified type
C0152990|T047|AB|045.01|ICD9CM|Ac bulbar polio-type 1|Ac bulbar polio-type 1
C0152990|T047|PT|045.01|ICD9CM|Acute paralytic poliomyelitis specified as bulbar, poliovirus type I|Acute paralytic poliomyelitis specified as bulbar, poliovirus type I
C0152991|T047|AB|045.02|ICD9CM|Ac bulbar polio-type 2|Ac bulbar polio-type 2
C0152991|T047|PT|045.02|ICD9CM|Acute paralytic poliomyelitis specified as bulbar, poliovirus type II|Acute paralytic poliomyelitis specified as bulbar, poliovirus type II
C0152992|T047|AB|045.03|ICD9CM|Ac bulbar polio-type 3|Ac bulbar polio-type 3
C0152992|T047|PT|045.03|ICD9CM|Acute paralytic poliomyelitis specified as bulbar, poliovirus type III|Acute paralytic poliomyelitis specified as bulbar, poliovirus type III
C0152993|T047|HT|045.1|ICD9CM|Acute poliomyelitis with other paralysis|Acute poliomyelitis with other paralysis
C0152994|T047|PT|045.10|ICD9CM|Acute poliomyelitis with other paralysis, poliovirus, unspecified type|Acute poliomyelitis with other paralysis, poliovirus, unspecified type
C0152994|T047|AB|045.10|ICD9CM|Paral polio NEC-type NOS|Paral polio NEC-type NOS
C0152995|T047|PT|045.11|ICD9CM|Acute poliomyelitis with other paralysis, poliovirus type I|Acute poliomyelitis with other paralysis, poliovirus type I
C0152995|T047|AB|045.11|ICD9CM|Paral polio NEC-type 1|Paral polio NEC-type 1
C0152996|T047|PT|045.12|ICD9CM|Acute poliomyelitis with other paralysis, poliovirus type II|Acute poliomyelitis with other paralysis, poliovirus type II
C0152996|T047|AB|045.12|ICD9CM|Paral polio NEC-type 2|Paral polio NEC-type 2
C0152997|T047|PT|045.13|ICD9CM|Acute poliomyelitis with other paralysis, poliovirus type III|Acute poliomyelitis with other paralysis, poliovirus type III
C0152997|T047|AB|045.13|ICD9CM|Paral polio NEC-type 3|Paral polio NEC-type 3
C0152998|T047|HT|045.2|ICD9CM|Acute nonparalytic poliomyelitis|Acute nonparalytic poliomyelitis
C0152998|T047|PT|045.20|ICD9CM|Acute nonparalytic poliomyelitis, poliovirus, unspecified type|Acute nonparalytic poliomyelitis, poliovirus, unspecified type
C0152998|T047|AB|045.20|ICD9CM|Nonparaly polio-type NOS|Nonparaly polio-type NOS
C1112685|T047|PT|045.21|ICD9CM|Acute nonparalytic poliomyelitis, poliovirus type I|Acute nonparalytic poliomyelitis, poliovirus type I
C1112685|T047|AB|045.21|ICD9CM|Nonparalyt polio-type 1|Nonparalyt polio-type 1
C1112686|T047|PT|045.22|ICD9CM|Acute nonparalytic poliomyelitis, poliovirus type II|Acute nonparalytic poliomyelitis, poliovirus type II
C1112686|T047|AB|045.22|ICD9CM|Nonparalyt polio-type 2|Nonparalyt polio-type 2
C1112687|T047|PT|045.23|ICD9CM|Acute nonparalytic poliomyelitis, poliovirus type III|Acute nonparalytic poliomyelitis, poliovirus type III
C1112687|T047|AB|045.23|ICD9CM|Nonparalyt polio-type 3|Nonparalyt polio-type 3
C0032371|T047|HT|045.9|ICD9CM|Acute poliomyelitis, unspecified|Acute poliomyelitis, unspecified
C0374998|T047|AB|045.90|ICD9CM|Ac polio NOS-type NOS|Ac polio NOS-type NOS
C0374998|T047|PT|045.90|ICD9CM|Acute poliomyelitis, unspecified, poliovirus, unspecified type|Acute poliomyelitis, unspecified, poliovirus, unspecified type
C0153004|T047|AB|045.91|ICD9CM|Ac polio NOS-type 1|Ac polio NOS-type 1
C0153004|T047|PT|045.91|ICD9CM|Acute poliomyelitis, unspecified, poliovirus type I|Acute poliomyelitis, unspecified, poliovirus type I
C0153005|T047|AB|045.92|ICD9CM|Ac polio NOS-type 2|Ac polio NOS-type 2
C0153005|T047|PT|045.92|ICD9CM|Acute poliomyelitis, unspecified, poliovirus type II|Acute poliomyelitis, unspecified, poliovirus type II
C0153006|T047|AB|045.93|ICD9CM|Ac polio NOS-type 3|Ac polio NOS-type 3
C0153006|T047|PT|045.93|ICD9CM|Acute poliomyelitis, unspecified, poliovirus type III|Acute poliomyelitis, unspecified, poliovirus type III
C2349761|T047|HT|046|ICD9CM|Slow virus infections and prion diseases of central nervous system|Slow virus infections and prion diseases of central nervous system
C0022802|T047|AB|046.0|ICD9CM|Kuru|Kuru
C0022802|T047|PT|046.0|ICD9CM|Kuru|Kuru
C0022336|T047|HT|046.1|ICD9CM|Jakob-Creutzfeldt disease|Jakob-Creutzfeldt disease
C0376329|T047|PT|046.11|ICD9CM|Variant Creutzfeldt-Jakob disease|Variant Creutzfeldt-Jakob disease
C0376329|T047|AB|046.11|ICD9CM|Varnt Creutzfeldt-Jakob|Varnt Creutzfeldt-Jakob
C2349756|T047|AB|046.19|ICD9CM|Creutzfldt-Jakob NEC/NOS|Creutzfldt-Jakob NEC/NOS
C2349756|T047|PT|046.19|ICD9CM|Other and unspecified Creutzfeldt-Jakob disease|Other and unspecified Creutzfeldt-Jakob disease
C0038522|T047|AB|046.2|ICD9CM|Subac scleros panenceph|Subac scleros panenceph
C0038522|T047|PT|046.2|ICD9CM|Subacute sclerosing panencephalitis|Subacute sclerosing panencephalitis
C0023524|T047|AB|046.3|ICD9CM|Prog multifoc leukoencep|Prog multifoc leukoencep
C0023524|T047|PT|046.3|ICD9CM|Progressive multifocal leukoencephalopathy|Progressive multifocal leukoencephalopathy
C2349760|T047|HT|046.7|ICD9CM|Other specified prion diseases of central nervous system|Other specified prion diseases of central nervous system
C0017495|T047|PT|046.71|ICD9CM|Gerstmann-Sträussler-Scheinker syndrome|Gerstmann-Sträussler-Scheinker syndrome
C0017495|T047|AB|046.71|ICD9CM|Gerstmn-Straus-Schnk syn|Gerstmn-Straus-Schnk syn
C0206042|T047|PT|046.72|ICD9CM|Fatal familial insomnia|Fatal familial insomnia
C0206042|T047|AB|046.72|ICD9CM|Fatal familial insomnia|Fatal familial insomnia
C2349759|T047|PT|046.79|ICD9CM|Other and unspecified prion disease of central nervous system|Other and unspecified prion disease of central nervous system
C2349759|T047|AB|046.79|ICD9CM|Prion dis of CNS NEC/NOS|Prion dis of CNS NEC/NOS
C0153007|T047|AB|046.8|ICD9CM|Cns slow virus infec NEC|Cns slow virus infec NEC
C0153007|T047|PT|046.8|ICD9CM|Other specified slow virus infection of central nervous system|Other specified slow virus infection of central nervous system
C0153008|T047|AB|046.9|ICD9CM|Cns slow virus infec NOS|Cns slow virus infec NOS
C0153008|T047|PT|046.9|ICD9CM|Unspecified slow virus infection of central nervous system|Unspecified slow virus infection of central nervous system
C0276430|T047|HT|047|ICD9CM|Meningitis due to enterovirus|Meningitis due to enterovirus
C0276431|T047|AB|047.0|ICD9CM|Coxsackie virus mening|Coxsackie virus mening
C0276431|T047|PT|047.0|ICD9CM|Meningitis due to coxsackie virus|Meningitis due to coxsackie virus
C0338388|T047|AB|047.1|ICD9CM|Echo virus meningitis|Echo virus meningitis
C0338388|T047|PT|047.1|ICD9CM|Meningitis due to echo virus|Meningitis due to echo virus
C0029843|T047|PT|047.8|ICD9CM|Other specified viral meningitis|Other specified viral meningitis
C0029843|T047|AB|047.8|ICD9CM|Viral meningitis NEC|Viral meningitis NEC
C0025297|T047|PT|047.9|ICD9CM|Unspecified viral meningitis|Unspecified viral meningitis
C0025297|T047|AB|047.9|ICD9CM|Viral meningitis NOS|Viral meningitis NOS
C0153012|T047|AB|048|ICD9CM|Oth enteroviral cns dis|Oth enteroviral cns dis
C0153012|T047|PT|048|ICD9CM|Other enterovirus diseases of central nervous system|Other enterovirus diseases of central nervous system
C0153013|T047|HT|049|ICD9CM|Other non-arthropod-borne viral diseases of central nervous system|Other non-arthropod-borne viral diseases of central nervous system
C0153014|T047|AB|049.0|ICD9CM|Lymphocytic choriomening|Lymphocytic choriomening
C0153014|T047|PT|049.0|ICD9CM|Lymphocytic choriomeningitis|Lymphocytic choriomeningitis
C0153015|T047|AB|049.1|ICD9CM|Adenoviral meningitis|Adenoviral meningitis
C0153015|T047|PT|049.1|ICD9CM|Meningitis due to adenovirus|Meningitis due to adenovirus
C0029818|T047|PT|049.8|ICD9CM|Other specified non-arthropod-borne viral diseases of central nervous system|Other specified non-arthropod-borne viral diseases of central nervous system
C0029818|T047|AB|049.8|ICD9CM|Viral encephalitis NEC|Viral encephalitis NEC
C0276148|T047|PT|049.9|ICD9CM|Unspecified non-arthropod-borne viral diseases of central nervous system|Unspecified non-arthropod-borne viral diseases of central nervous system
C0276148|T047|AB|049.9|ICD9CM|Viral encephalitis NOS|Viral encephalitis NOS
C0037354|T047|HT|050|ICD9CM|Smallpox|Smallpox
C2712640|T047|HT|050-059.99|ICD9CM|VIRAL DISEASES GENERALLY ACCOMPANIED BY EXANTHEM|VIRAL DISEASES GENERALLY ACCOMPANIED BY EXANTHEM
C1812609|T047|AB|050.0|ICD9CM|Variola major|Variola major
C1812609|T047|PT|050.0|ICD9CM|Variola major|Variola major
C0001906|T047|AB|050.1|ICD9CM|Alastrim|Alastrim
C0001906|T047|PT|050.1|ICD9CM|Alastrim|Alastrim
C0037358|T047|AB|050.2|ICD9CM|Modified smallpox|Modified smallpox
C0037358|T047|PT|050.2|ICD9CM|Modified smallpox|Modified smallpox
C0037354|T047|AB|050.9|ICD9CM|Smallpox NOS|Smallpox NOS
C0037354|T047|PT|050.9|ICD9CM|Smallpox, unspecified|Smallpox, unspecified
C0153016|T047|HT|051|ICD9CM|Cowpox and paravaccinia|Cowpox and paravaccinia
C2349762|T047|HT|051.0|ICD9CM|Cowpox and vaccinia not from vaccination|Cowpox and vaccinia not from vaccination
C0010232|T047|PT|051.01|ICD9CM|Cowpox|Cowpox
C0010232|T047|AB|051.01|ICD9CM|Cowpox|Cowpox
C0864706|T033|AB|051.02|ICD9CM|Vaccinia n/f vaccination|Vaccinia n/f vaccination
C0864706|T033|PT|051.02|ICD9CM|Vaccinia not from vaccination|Vaccinia not from vaccination
C0026143|T047|AB|051.1|ICD9CM|Pseudocowpox|Pseudocowpox
C0026143|T047|PT|051.1|ICD9CM|Pseudocowpox|Pseudocowpox
C0013570|T047|AB|051.2|ICD9CM|Contagious pustular derm|Contagious pustular derm
C0013570|T047|PT|051.2|ICD9CM|Contagious pustular dermatitis|Contagious pustular dermatitis
C0026143|T047|AB|051.9|ICD9CM|Paravaccinia NOS|Paravaccinia NOS
C0026143|T047|PT|051.9|ICD9CM|Paravaccinia, unspecified|Paravaccinia, unspecified
C0008049|T047|HT|052|ICD9CM|Chickenpox|Chickenpox
C0153017|T047|AB|052.0|ICD9CM|Postvaricella encephalit|Postvaricella encephalit
C0153017|T047|PT|052.0|ICD9CM|Postvaricella encephalitis|Postvaricella encephalitis
C0153018|T047|PT|052.1|ICD9CM|Varicella (hemorrhagic) pneumonitis|Varicella (hemorrhagic) pneumonitis
C0153018|T047|AB|052.1|ICD9CM|Varicella pneumonitis|Varicella pneumonitis
C1719295|T047|PT|052.2|ICD9CM|Postvaricella myelitis|Postvaricella myelitis
C1719295|T047|AB|052.2|ICD9CM|Postvaricella myelitis|Postvaricella myelitis
C0153019|T047|PT|052.7|ICD9CM|Chickenpox with other specified complications|Chickenpox with other specified complications
C0153019|T047|AB|052.7|ICD9CM|Varicella complicat NEC|Varicella complicat NEC
C0348187|T047|PT|052.8|ICD9CM|Chickenpox with unspecified complication|Chickenpox with unspecified complication
C0348187|T047|AB|052.8|ICD9CM|Varicella complicat NOS|Varicella complicat NOS
C0348188|T047|AB|052.9|ICD9CM|Varicella uncomplicated|Varicella uncomplicated
C0348188|T047|PT|052.9|ICD9CM|Varicella without mention of complication|Varicella without mention of complication
C0019360|T047|HT|053|ICD9CM|Herpes zoster|Herpes zoster
C0700503|T047|AB|053.0|ICD9CM|Herpes zoster meningitis|Herpes zoster meningitis
C0700503|T047|PT|053.0|ICD9CM|Herpes zoster with meningitis|Herpes zoster with meningitis
C0153022|T047|HT|053.1|ICD9CM|Herpes zoster with other nervous system complications|Herpes zoster with other nervous system complications
C1264623|T047|AB|053.10|ICD9CM|H zoster nerv syst NOS|H zoster nerv syst NOS
C1264623|T047|PT|053.10|ICD9CM|Herpes zoster with unspecified nervous system complication|Herpes zoster with unspecified nervous system complication
C0017409|T047|AB|053.11|ICD9CM|Geniculate herpes zoster|Geniculate herpes zoster
C0017409|T047|PT|053.11|ICD9CM|Geniculate herpes zoster|Geniculate herpes zoster
C0153024|T047|AB|053.12|ICD9CM|Postherpes trigem neural|Postherpes trigem neural
C0153024|T047|PT|053.12|ICD9CM|Postherpetic trigeminal neuralgia|Postherpetic trigeminal neuralgia
C0153025|T047|AB|053.13|ICD9CM|Postherpes polyneuropath|Postherpes polyneuropath
C0153025|T047|PT|053.13|ICD9CM|Postherpetic polyneuropathy|Postherpetic polyneuropathy
C1719297|T047|PT|053.14|ICD9CM|Herpes zoster myelitis|Herpes zoster myelitis
C1719297|T047|AB|053.14|ICD9CM|Herpes zoster myelitis|Herpes zoster myelitis
C0153022|T047|AB|053.19|ICD9CM|H zoster nerv syst NEC|H zoster nerv syst NEC
C0153022|T047|PT|053.19|ICD9CM|Herpes zoster with other nervous system complications|Herpes zoster with other nervous system complications
C0019364|T047|HT|053.2|ICD9CM|Herpes zoster with ophthalmic complications|Herpes zoster with ophthalmic complications
C0019362|T047|PT|053.20|ICD9CM|Herpes zoster dermatitis of eyelid|Herpes zoster dermatitis of eyelid
C0019362|T047|AB|053.20|ICD9CM|Herpes zoster of eyelid|Herpes zoster of eyelid
C0153027|T047|AB|053.21|ICD9CM|H zoster keratoconjunct|H zoster keratoconjunct
C0153027|T047|PT|053.21|ICD9CM|Herpes zoster keratoconjunctivitis|Herpes zoster keratoconjunctivitis
C0153028|T047|AB|053.22|ICD9CM|H zoster iridocyclitis|H zoster iridocyclitis
C0153028|T047|PT|053.22|ICD9CM|Herpes zoster iridocyclitis|Herpes zoster iridocyclitis
C0795698|T047|AB|053.29|ICD9CM|Herpes zoster of eye NEC|Herpes zoster of eye NEC
C0795698|T047|PT|053.29|ICD9CM|Herpes zoster with other ophthalmic complications|Herpes zoster with other ophthalmic complications
C0153030|T047|HT|053.7|ICD9CM|Herpes zoster with other specified complications|Herpes zoster with other specified complications
C0153031|T047|AB|053.71|ICD9CM|H zoster otitis externa|H zoster otitis externa
C0153031|T047|PT|053.71|ICD9CM|Otitis externa due to herpes zoster|Otitis externa due to herpes zoster
C0153030|T047|AB|053.79|ICD9CM|H zoster complicated NEC|H zoster complicated NEC
C0153030|T047|PT|053.79|ICD9CM|Herpes zoster with other specified complications|Herpes zoster with other specified complications
C0276249|T047|AB|053.8|ICD9CM|H zoster complicated NOS|H zoster complicated NOS
C0276249|T047|PT|053.8|ICD9CM|Herpes zoster with unspecified complication|Herpes zoster with unspecified complication
C0019366|T047|AB|053.9|ICD9CM|Herpes zoster NOS|Herpes zoster NOS
C0019366|T047|PT|053.9|ICD9CM|Herpes zoster without mention of complication|Herpes zoster without mention of complication
C0019348|T047|HT|054|ICD9CM|Herpes simplex|Herpes simplex
C0936250|T047|AB|054.0|ICD9CM|Eczema herpeticum|Eczema herpeticum
C0936250|T047|PT|054.0|ICD9CM|Eczema herpeticum|Eczema herpeticum
C0019342|T047|HT|054.1|ICD9CM|Genital herpes|Genital herpes
C0019342|T047|AB|054.10|ICD9CM|Genital herpes NOS|Genital herpes NOS
C0019342|T047|PT|054.10|ICD9CM|Genital herpes, unspecified|Genital herpes, unspecified
C0019386|T047|AB|054.11|ICD9CM|Herpetic vulvovaginitis|Herpetic vulvovaginitis
C0019386|T047|PT|054.11|ICD9CM|Herpetic vulvovaginitis|Herpetic vulvovaginitis
C0153033|T047|AB|054.12|ICD9CM|Herpetic ulcer of vulva|Herpetic ulcer of vulva
C0153033|T047|PT|054.12|ICD9CM|Herpetic ulceration of vulva|Herpetic ulceration of vulva
C0153034|T047|AB|054.13|ICD9CM|Herpetic infect of penis|Herpetic infect of penis
C0153034|T047|PT|054.13|ICD9CM|Herpetic infection of penis|Herpetic infection of penis
C0029627|T047|AB|054.19|ICD9CM|Genital herpes NEC|Genital herpes NEC
C0029627|T047|PT|054.19|ICD9CM|Other genital herpes|Other genital herpes
C0376379|T047|AB|054.2|ICD9CM|Herpetic gingivostomat|Herpetic gingivostomat
C0376379|T047|PT|054.2|ICD9CM|Herpetic gingivostomatitis|Herpetic gingivostomatitis
C0019385|T047|AB|054.3|ICD9CM|Herpetic encephalitis|Herpetic encephalitis
C0019385|T047|PT|054.3|ICD9CM|Herpetic meningoencephalitis|Herpetic meningoencephalitis
C0153036|T047|HT|054.4|ICD9CM|Herpes simplex with ophthalmic complications|Herpes simplex with ophthalmic complications
C0153036|T047|AB|054.40|ICD9CM|Herpes simplex eye NOS|Herpes simplex eye NOS
C0153036|T047|PT|054.40|ICD9CM|Herpes simplex with unspecified ophthalmic complication|Herpes simplex with unspecified ophthalmic complication
C0153037|T047|PT|054.41|ICD9CM|Herpes simplex dermatitis of eyelid|Herpes simplex dermatitis of eyelid
C0153037|T047|AB|054.41|ICD9CM|Herpes simplex of eyelid|Herpes simplex of eyelid
C0022570|T047|AB|054.42|ICD9CM|Dendritic keratitis|Dendritic keratitis
C0022570|T047|PT|054.42|ICD9CM|Dendritic keratitis|Dendritic keratitis
C0153038|T047|AB|054.43|ICD9CM|H simplex keratitis|H simplex keratitis
C0153038|T047|PT|054.43|ICD9CM|Herpes simplex disciform keratitis|Herpes simplex disciform keratitis
C0153039|T047|AB|054.44|ICD9CM|H simplex iridocyclitis|H simplex iridocyclitis
C0153039|T047|PT|054.44|ICD9CM|Herpes simplex iridocyclitis|Herpes simplex iridocyclitis
C0153040|T047|AB|054.49|ICD9CM|Herpes simplex eye NEC|Herpes simplex eye NEC
C0153040|T047|PT|054.49|ICD9CM|Herpes simplex with other ophthalmic complications|Herpes simplex with other ophthalmic complications
C0153041|T047|AB|054.5|ICD9CM|Herpetic septicemia|Herpetic septicemia
C0153041|T047|PT|054.5|ICD9CM|Herpetic septicemia|Herpetic septicemia
C0153042|T047|AB|054.6|ICD9CM|Herpetic whitlow|Herpetic whitlow
C0153042|T047|PT|054.6|ICD9CM|Herpetic whitlow|Herpetic whitlow
C0153043|T047|HT|054.7|ICD9CM|Herpes simplex with other specified complications|Herpes simplex with other specified complications
C0019359|T047|AB|054.71|ICD9CM|Visceral herpes simplex|Visceral herpes simplex
C0019359|T047|PT|054.71|ICD9CM|Visceral herpes simplex|Visceral herpes simplex
C0153045|T047|AB|054.72|ICD9CM|H simplex meningitis|H simplex meningitis
C0153045|T047|PT|054.72|ICD9CM|Herpes simplex meningitis|Herpes simplex meningitis
C0153046|T047|AB|054.73|ICD9CM|H simplex otitis externa|H simplex otitis externa
C0153046|T047|PT|054.73|ICD9CM|Herpes simplex otitis externa|Herpes simplex otitis externa
C1719298|T047|PT|054.74|ICD9CM|Herpes simplex myelitis|Herpes simplex myelitis
C1719298|T047|AB|054.74|ICD9CM|Herpes simplex myelitis|Herpes simplex myelitis
C0153043|T047|AB|054.79|ICD9CM|H simplex complicat NEC|H simplex complicat NEC
C0153043|T047|PT|054.79|ICD9CM|Herpes simplex with other specified complications|Herpes simplex with other specified complications
C0153047|T047|AB|054.8|ICD9CM|H simplex complicat NOS|H simplex complicat NOS
C0153047|T047|PT|054.8|ICD9CM|Herpes simplex with unspecified complication|Herpes simplex with unspecified complication
C0392646|T047|AB|054.9|ICD9CM|Herpes simplex NOS|Herpes simplex NOS
C0392646|T047|PT|054.9|ICD9CM|Herpes simplex without mention of complication|Herpes simplex without mention of complication
C0025007|T047|HT|055|ICD9CM|Measles|Measles
C0153048|T047|AB|055.0|ICD9CM|Postmeasles encephalitis|Postmeasles encephalitis
C0153048|T047|PT|055.0|ICD9CM|Postmeasles encephalitis|Postmeasles encephalitis
C1112452|T047|AB|055.1|ICD9CM|Postmeasles pneumonia|Postmeasles pneumonia
C1112452|T047|PT|055.1|ICD9CM|Postmeasles pneumonia|Postmeasles pneumonia
C0153050|T047|AB|055.2|ICD9CM|Postmeasles otitis media|Postmeasles otitis media
C0153050|T047|PT|055.2|ICD9CM|Postmeasles otitis media|Postmeasles otitis media
C0153051|T047|HT|055.7|ICD9CM|Measles with other specified complications|Measles with other specified complications
C0153052|T047|AB|055.71|ICD9CM|Measles keratitis|Measles keratitis
C0153052|T047|PT|055.71|ICD9CM|Measles keratoconjunctivitis|Measles keratoconjunctivitis
C0153051|T047|AB|055.79|ICD9CM|Measles complication NEC|Measles complication NEC
C0153051|T047|PT|055.79|ICD9CM|Measles with other specified complications|Measles with other specified complications
C0153053|T047|AB|055.8|ICD9CM|Measles complication NOS|Measles complication NOS
C0153053|T047|PT|055.8|ICD9CM|Measles with unspecified complication|Measles with unspecified complication
C0392650|T047|AB|055.9|ICD9CM|Measles uncomplicated|Measles uncomplicated
C0392650|T047|PT|055.9|ICD9CM|Measles without mention of complication|Measles without mention of complication
C0035920|T047|HT|056|ICD9CM|Rubella|Rubella
C2937267|T047|HT|056.0|ICD9CM|Rubella with neurological complications|Rubella with neurological complications
C2937267|T047|AB|056.00|ICD9CM|Rubella nerve compl NOS|Rubella nerve compl NOS
C2937267|T047|PT|056.00|ICD9CM|Rubella with unspecified neurological complication|Rubella with unspecified neurological complication
C0033359|T047|PT|056.01|ICD9CM|Encephalomyelitis due to rubella|Encephalomyelitis due to rubella
C0033359|T047|AB|056.01|ICD9CM|Rubella encephalitis|Rubella encephalitis
C0153057|T047|AB|056.09|ICD9CM|Rubella nerve compl NEC|Rubella nerve compl NEC
C0153057|T047|PT|056.09|ICD9CM|Rubella with other neurological complications|Rubella with other neurological complications
C0153058|T047|HT|056.7|ICD9CM|Rubella with other specified complications|Rubella with other specified complications
C0276308|T047|AB|056.71|ICD9CM|Arthritis due to rubella|Arthritis due to rubella
C0276308|T047|PT|056.71|ICD9CM|Arthritis due to rubella|Arthritis due to rubella
C0153058|T047|AB|056.79|ICD9CM|Rubella complication NEC|Rubella complication NEC
C0153058|T047|PT|056.79|ICD9CM|Rubella with other specified complications|Rubella with other specified complications
C0153060|T047|AB|056.8|ICD9CM|Rubella complication NOS|Rubella complication NOS
C0153060|T047|PT|056.8|ICD9CM|Rubella with unspecified complications|Rubella with unspecified complications
C0348194|T047|AB|056.9|ICD9CM|Rubella uncomplicated|Rubella uncomplicated
C0348194|T047|PT|056.9|ICD9CM|Rubella without mention of complication|Rubella without mention of complication
C0153061|T047|HT|057|ICD9CM|Other viral exanthemata|Other viral exanthemata
C0085273|T047|AB|057.0|ICD9CM|Erythema infectiosum|Erythema infectiosum
C0085273|T047|PT|057.0|ICD9CM|Erythema infectiosum (fifth disease)|Erythema infectiosum (fifth disease)
C0029841|T047|PT|057.8|ICD9CM|Other specified viral exanthemata|Other specified viral exanthemata
C0029841|T047|AB|057.8|ICD9CM|Viral exanthemata NEC|Viral exanthemata NEC
C0153062|T047|PT|057.9|ICD9CM|Viral exanthem, unspecified|Viral exanthem, unspecified
C0153062|T047|AB|057.9|ICD9CM|Viral exanthemata NOS|Viral exanthemata NOS
C1955628|T047|HT|058|ICD9CM|Other human herpesvirus|Other human herpesvirus
C0015231|T047|HT|058.1|ICD9CM|Roseola infantum|Roseola infantum
C0015231|T047|AB|058.10|ICD9CM|Roseola infantum NOS|Roseola infantum NOS
C0015231|T047|PT|058.10|ICD9CM|Roseola infantum, unspecified|Roseola infantum, unspecified
C2240388|T047|AB|058.11|ICD9CM|Roseola infant d/t HHV-6|Roseola infant d/t HHV-6
C2240388|T047|PT|058.11|ICD9CM|Roseola infantum due to human herpesvirus 6|Roseola infantum due to human herpesvirus 6
C1274329|T047|AB|058.12|ICD9CM|Roseola infant d/t HHV-7|Roseola infant d/t HHV-7
C1274329|T047|PT|058.12|ICD9CM|Roseola infantum due to human herpesvirus 7|Roseola infantum due to human herpesvirus 7
C1955630|T047|HT|058.2|ICD9CM|Other human herpesvirus encephalitis|Other human herpesvirus encephalitis
C1955629|T047|AB|058.21|ICD9CM|Human herpesvir 6 enceph|Human herpesvir 6 enceph
C1955629|T047|PT|058.21|ICD9CM|Human herpesvirus 6 encephalitis|Human herpesvirus 6 encephalitis
C1955630|T047|AB|058.29|ICD9CM|Human herpesvr encph NEC|Human herpesvr encph NEC
C1955630|T047|PT|058.29|ICD9CM|Other human herpesvirus encephalitis|Other human herpesvirus encephalitis
C1955633|T047|HT|058.8|ICD9CM|Other human herpesvirus infections|Other human herpesvirus infections
C0854530|T047|AB|058.81|ICD9CM|Human herpesvirus 6 infc|Human herpesvirus 6 infc
C0854530|T047|PT|058.81|ICD9CM|Human herpesvirus 6 infection|Human herpesvirus 6 infection
C1504514|T047|AB|058.82|ICD9CM|Human herpesvirus 7 infc|Human herpesvirus 7 infc
C1504514|T047|PT|058.82|ICD9CM|Human herpesvirus 7 infection|Human herpesvirus 7 infection
C1955633|T047|AB|058.89|ICD9CM|Human herpesvirs inf NEC|Human herpesvirs inf NEC
C1955633|T047|PT|058.89|ICD9CM|Other human herpesvirus infection|Other human herpesvirus infection
C2349858|T047|HT|059|ICD9CM|Other poxvirus infections|Other poxvirus infections
C0348196|T047|HT|059.0|ICD9CM|Other orthopoxvirus infections|Other orthopoxvirus infections
C2349763|T047|AB|059.00|ICD9CM|Orthopoxvirus infect NOS|Orthopoxvirus infect NOS
C2349763|T047|PT|059.00|ICD9CM|Orthopoxvirus infection, unspecified|Orthopoxvirus infection, unspecified
C0276180|T047|PT|059.01|ICD9CM|Monkeypox|Monkeypox
C0276180|T047|AB|059.01|ICD9CM|Monkeypox|Monkeypox
C0348196|T047|AB|059.09|ICD9CM|Orthopoxvirus infect NEC|Orthopoxvirus infect NEC
C0348196|T047|PT|059.09|ICD9CM|Other orthopoxvirus infections|Other orthopoxvirus infections
C2349855|T047|HT|059.1|ICD9CM|Other parapoxvirus infections|Other parapoxvirus infections
C2368006|T047|PT|059.10|ICD9CM|Parapoxvirus infection, unspecified|Parapoxvirus infection, unspecified
C2368006|T047|AB|059.10|ICD9CM|Parapoxvirus infectn NOS|Parapoxvirus infectn NOS
C2349765|T047|PT|059.11|ICD9CM|Bovine stomatitis|Bovine stomatitis
C2349765|T047|AB|059.11|ICD9CM|Bovine stomatitis|Bovine stomatitis
C0276191|T047|PT|059.12|ICD9CM|Sealpox|Sealpox
C0276191|T047|AB|059.12|ICD9CM|Sealpox|Sealpox
C2349855|T047|PT|059.19|ICD9CM|Other parapoxvirus infections|Other parapoxvirus infections
C2349855|T047|AB|059.19|ICD9CM|Parapoxvirus infectn NEC|Parapoxvirus infectn NEC
C2349857|T047|HT|059.2|ICD9CM|Yatapoxvirus infections|Yatapoxvirus infections
C2349857|T047|PT|059.20|ICD9CM|Yatapoxvirus infection, unspecified|Yatapoxvirus infection, unspecified
C2349857|T047|AB|059.20|ICD9CM|Yatapoxvirus infectn NOS|Yatapoxvirus infectn NOS
C0276214|T047|PT|059.21|ICD9CM|Tanapox|Tanapox
C0276214|T047|AB|059.21|ICD9CM|Tanapox|Tanapox
C2349858|T047|PT|059.8|ICD9CM|Other poxvirus infections|Other poxvirus infections
C2349858|T047|AB|059.8|ICD9CM|Poxvirus infections NEC|Poxvirus infections NEC
C0032870|T047|AB|059.9|ICD9CM|Poxvirus infection NOS|Poxvirus infection NOS
C0032870|T047|PT|059.9|ICD9CM|Poxvirus infections, unspecified|Poxvirus infections, unspecified
C0043395|T047|HT|060|ICD9CM|Yellow fever|Yellow fever
C0003723|T047|HT|060-066.99|ICD9CM|ARTHROPOD-BORNE VIRAL DISEASES|ARTHROPOD-BORNE VIRAL DISEASES
C0043397|T047|AB|060.0|ICD9CM|Sylvatic yellow fever|Sylvatic yellow fever
C0043397|T047|PT|060.0|ICD9CM|Sylvatic yellow fever|Sylvatic yellow fever
C0043398|T047|AB|060.1|ICD9CM|Urban yellow fever|Urban yellow fever
C0043398|T047|PT|060.1|ICD9CM|Urban yellow fever|Urban yellow fever
C0043395|T047|AB|060.9|ICD9CM|Yellow fever NOS|Yellow fever NOS
C0043395|T047|PT|060.9|ICD9CM|Yellow fever, unspecified|Yellow fever, unspecified
C0011311|T047|AB|061|ICD9CM|Dengue|Dengue
C0011311|T047|PT|061|ICD9CM|Dengue|Dengue
C0751098|T047|HT|062|ICD9CM|Mosquito-borne viral encephalitis|Mosquito-borne viral encephalitis
C0014057|T047|AB|062.0|ICD9CM|Japanese encephalitis|Japanese encephalitis
C0014057|T047|PT|062.0|ICD9CM|Japanese encephalitis|Japanese encephalitis
C0153064|T047|AB|062.1|ICD9CM|West equine encephalitis|West equine encephalitis
C0153064|T047|PT|062.1|ICD9CM|Western equine encephalitis|Western equine encephalitis
C0153065|T047|AB|062.2|ICD9CM|East equine encephalitis|East equine encephalitis
C0153065|T047|PT|062.2|ICD9CM|Eastern equine encephalitis|Eastern equine encephalitis
C0014060|T047|AB|062.3|ICD9CM|St Louis encephalitis|St Louis encephalitis
C0014060|T047|PT|062.3|ICD9CM|St. Louis encephalitis|St. Louis encephalitis
C0153066|T047|AB|062.4|ICD9CM|Australian encephalitis|Australian encephalitis
C0153066|T047|PT|062.4|ICD9CM|Australian encephalitis|Australian encephalitis
C0014053|T047|AB|062.5|ICD9CM|California encephalitis|California encephalitis
C0014053|T047|PT|062.5|ICD9CM|California virus encephalitis|California virus encephalitis
C0348168|T047|AB|062.8|ICD9CM|Mosquit-borne enceph NEC|Mosquit-borne enceph NEC
C0348168|T047|PT|062.8|ICD9CM|Other specified mosquito-borne viral encephalitis|Other specified mosquito-borne viral encephalitis
C0751098|T047|AB|062.9|ICD9CM|Mosquit-borne enceph NOS|Mosquit-borne enceph NOS
C0751098|T047|PT|062.9|ICD9CM|Mosquito-borne viral encephalitis, unspecified|Mosquito-borne viral encephalitis, unspecified
C0014061|T047|HT|063|ICD9CM|Tick-borne viral encephalitis|Tick-borne viral encephalitis
C0015632|T047|AB|063.0|ICD9CM|Russia spr-summer enceph|Russia spr-summer enceph
C0015632|T047|PT|063.0|ICD9CM|Russian spring-summer [taiga] encephalitis|Russian spring-summer [taiga] encephalitis
C0024025|T047|AB|063.1|ICD9CM|Louping ill|Louping ill
C0024025|T047|PT|063.1|ICD9CM|Louping ill|Louping ill
C0014054|T047|AB|063.2|ICD9CM|Cent Europe encephalitis|Cent Europe encephalitis
C0014054|T047|PT|063.2|ICD9CM|Central european encephalitis|Central european encephalitis
C0029832|T047|PT|063.8|ICD9CM|Other specified tick-borne viral encephalitis|Other specified tick-borne viral encephalitis
C0029832|T047|AB|063.8|ICD9CM|Tick-borne enceph NEC|Tick-borne enceph NEC
C0014061|T047|AB|063.9|ICD9CM|Tick-borne enceph NOS|Tick-borne enceph NOS
C0014061|T047|PT|063.9|ICD9CM|Tick-borne viral encephalitis, unspecified|Tick-borne viral encephalitis, unspecified
C0153069|T047|AB|064|ICD9CM|Vir enceph arthropod NEC|Vir enceph arthropod NEC
C0153069|T047|PT|064|ICD9CM|Viral encephalitis transmitted by other and unspecified arthropods|Viral encephalitis transmitted by other and unspecified arthropods
C0003721|T047|HT|065|ICD9CM|Arthropod-borne hemorrhagic fever|Arthropod-borne hemorrhagic fever
C0019099|T047|AB|065.0|ICD9CM|Crimean hemorrhagic fev|Crimean hemorrhagic fev
C0019099|T047|PT|065.0|ICD9CM|Crimean hemorrhagic fever [CHF Congo virus]|Crimean hemorrhagic fever [CHF Congo virus]
C0019103|T047|AB|065.1|ICD9CM|Omsk hemorrhagic fever|Omsk hemorrhagic fever
C0019103|T047|PT|065.1|ICD9CM|Omsk hemorrhagic fever|Omsk hemorrhagic fever
C0022810|T047|AB|065.2|ICD9CM|Kyasanur forest disease|Kyasanur forest disease
C0022810|T047|PT|065.2|ICD9CM|Kyasanur forest disease|Kyasanur forest disease
C0153070|T047|PT|065.3|ICD9CM|Other tick-borne hemorrhagic fever|Other tick-borne hemorrhagic fever
C0153070|T047|AB|065.3|ICD9CM|Tick-borne hem fever NEC|Tick-borne hem fever NEC
C0153071|T047|AB|065.4|ICD9CM|Mosquito-borne hem fever|Mosquito-borne hem fever
C0153071|T047|PT|065.4|ICD9CM|Mosquito-borne hemorrhagic fever|Mosquito-borne hemorrhagic fever
C0153072|T047|AB|065.8|ICD9CM|Arthropod hem fever NEC|Arthropod hem fever NEC
C0153072|T047|PT|065.8|ICD9CM|Other specified arthropod-borne hemorrhagic fever|Other specified arthropod-borne hemorrhagic fever
C0003721|T047|AB|065.9|ICD9CM|Arthropod hem fever NOS|Arthropod hem fever NOS
C0003721|T047|PT|065.9|ICD9CM|Arthropod-borne hemorrhagic fever, unspecified|Arthropod-borne hemorrhagic fever, unspecified
C0153073|T047|HT|066|ICD9CM|Other arthropod-borne viral diseases|Other arthropod-borne viral diseases
C0030372|T047|AB|066.0|ICD9CM|Phlebotomus fever|Phlebotomus fever
C0030372|T047|PT|066.0|ICD9CM|Phlebotomus fever|Phlebotomus fever
C0040199|T047|AB|066.1|ICD9CM|Tick-borne fever|Tick-borne fever
C0040199|T047|PT|066.1|ICD9CM|Tick-borne fever|Tick-borne fever
C0014078|T047|AB|066.2|ICD9CM|Venezuelan equine fever|Venezuelan equine fever
C0014078|T047|PT|066.2|ICD9CM|Venezuelan equine fever|Venezuelan equine fever
C0029667|T047|AB|066.3|ICD9CM|Mosquito-borne fever NEC|Mosquito-borne fever NEC
C0029667|T047|PT|066.3|ICD9CM|Other mosquito-borne fever|Other mosquito-borne fever
C0043124|T047|HT|066.4|ICD9CM|West Nile fever|West Nile fever
C0043124|T047|AB|066.40|ICD9CM|West Nile Fever NOS|West Nile Fever NOS
C0043124|T047|PT|066.40|ICD9CM|West Nile Fever, unspecified|West Nile Fever, unspecified
C0751583|T047|AB|066.41|ICD9CM|West Nile Fever w/enceph|West Nile Fever w/enceph
C0751583|T047|PT|066.41|ICD9CM|West Nile Fever with encephalitis|West Nile Fever with encephalitis
C1456259|T047|PT|066.42|ICD9CM|West Nile Fever with other neurologic manifestation|West Nile Fever with other neurologic manifestation
C1456259|T047|AB|066.42|ICD9CM|West Nile neuro man NEC|West Nile neuro man NEC
C1456260|T047|PT|066.49|ICD9CM|West Nile Fever with other complications|West Nile Fever with other complications
C1456260|T047|AB|066.49|ICD9CM|West Nile w complic NEC|West Nile w complic NEC
C0153074|T047|AB|066.8|ICD9CM|Arthropod virus NEC|Arthropod virus NEC
C0153074|T047|PT|066.8|ICD9CM|Other specified arthropod-borne viral diseases|Other specified arthropod-borne viral diseases
C0003723|T047|AB|066.9|ICD9CM|Arthropod virus NOS|Arthropod virus NOS
C0003723|T047|PT|066.9|ICD9CM|Arthropod-borne viral disease, unspecified|Arthropod-borne viral disease, unspecified
C0042721|T047|HT|070|ICD9CM|Viral hepatitis|Viral hepatitis
C0153111|T047|HT|070-079.99|ICD9CM|OTHER DISEASES DUE TO VIRUSES AND CHLAMYDIAE|OTHER DISEASES DUE TO VIRUSES AND CHLAMYDIAE
C0153075|T047|AB|070.0|ICD9CM|Hepatitis A with coma|Hepatitis A with coma
C0153075|T047|PT|070.0|ICD9CM|Viral hepatitis A with hepatic coma|Viral hepatitis A with hepatic coma
C1290810|T047|AB|070.1|ICD9CM|Hepatitis A w/o coma|Hepatitis A w/o coma
C1290810|T047|PT|070.1|ICD9CM|Viral hepatitis A without mention of hepatic coma|Viral hepatitis A without mention of hepatic coma
C0153076|T047|HT|070.2|ICD9CM|Viral hepatitis B with hepatic coma|Viral hepatitis B with hepatic coma
C0375000|T047|AB|070.20|ICD9CM|Hpt B acte coma wo dlta|Hpt B acte coma wo dlta
C0375000|T047|PT|070.20|ICD9CM|Viral hepatitis B with hepatic coma, acute or unspecified, without mention of hepatitis delta|Viral hepatitis B with hepatic coma, acute or unspecified, without mention of hepatitis delta
C0375001|T047|AB|070.21|ICD9CM|Hpt B acte coma w dlta|Hpt B acte coma w dlta
C0375001|T047|PT|070.21|ICD9CM|Viral hepatitis B with hepatic coma, acute or unspecified, with hepatitis delta|Viral hepatitis B with hepatic coma, acute or unspecified, with hepatitis delta
C0375002|T047|PT|070.22|ICD9CM|Chronic viral hepatitis B with hepatic coma without hepatitis delta|Chronic viral hepatitis B with hepatic coma without hepatitis delta
C0375002|T047|AB|070.22|ICD9CM|Hpt B chrn coma wo dlta|Hpt B chrn coma wo dlta
C0375003|T047|PT|070.23|ICD9CM|Chronic viral hepatitis B with hepatic coma with hepatitis delta|Chronic viral hepatitis B with hepatic coma with hepatitis delta
C0375003|T047|AB|070.23|ICD9CM|Hpt B chrn coma w dlta|Hpt B chrn coma w dlta
C0700211|T047|HT|070.3|ICD9CM|Viral hepatitis B without mention of hepatic coma|Viral hepatitis B without mention of hepatic coma
C0375004|T047|AB|070.30|ICD9CM|Hpt B acte wo cm wo dlta|Hpt B acte wo cm wo dlta
C0375005|T047|AB|070.31|ICD9CM|Hpt B acte wo cm w dlta|Hpt B acte wo cm w dlta
C0375005|T047|PT|070.31|ICD9CM|Viral hepatitis B without mention of hepatic coma, acute or unspecified, with hepatitis delta|Viral hepatitis B without mention of hepatic coma, acute or unspecified, with hepatitis delta
C0375006|T047|PT|070.32|ICD9CM|Chronic viral hepatitis B without mention of hepatic coma without mention of hepatitis delta|Chronic viral hepatitis B without mention of hepatic coma without mention of hepatitis delta
C0375006|T047|AB|070.32|ICD9CM|Hpt B chrn wo cm wo dlta|Hpt B chrn wo cm wo dlta
C0375007|T047|PT|070.33|ICD9CM|Chronic viral hepatitis B without mention of hepatic coma with hepatitis delta|Chronic viral hepatitis B without mention of hepatic coma with hepatitis delta
C0375007|T047|AB|070.33|ICD9CM|Hpt B chrn wo cm w dlta|Hpt B chrn wo cm w dlta
C0153081|T047|HT|070.4|ICD9CM|Other specified viral hepatitis with hepatic coma|Other specified viral hepatitis with hepatic coma
C1456261|T047|PT|070.41|ICD9CM|Acute hepatitis C with hepatic coma|Acute hepatitis C with hepatic coma
C1456261|T047|AB|070.41|ICD9CM|Hpt C acute w hepat Coma|Hpt C acute w hepat Coma
C0153083|T047|PT|070.42|ICD9CM|Hepatitis delta without mention of active hepatitis B disease with hepatic coma|Hepatitis delta without mention of active hepatitis B disease with hepatic coma
C0153083|T047|AB|070.42|ICD9CM|Hpt dlt wo b w hpt coma|Hpt dlt wo b w hpt coma
C0153084|T047|PT|070.43|ICD9CM|Hepatitis E with hepatic coma|Hepatitis E with hepatic coma
C0153084|T047|AB|070.43|ICD9CM|Hpt E w hepat Coma|Hpt E w hepat Coma
C0375009|T047|AB|070.44|ICD9CM|Chrnc hpt C w hepat Coma|Chrnc hpt C w hepat Coma
C0375009|T047|PT|070.44|ICD9CM|Chronic hepatitis C with hepatic coma|Chronic hepatitis C with hepatic coma
C0153081|T047|AB|070.49|ICD9CM|Oth vrl hepat w hpt coma|Oth vrl hepat w hpt coma
C0153081|T047|PT|070.49|ICD9CM|Other specified viral hepatitis with hepatic coma|Other specified viral hepatitis with hepatic coma
C0153085|T047|HT|070.5|ICD9CM|Other specified viral hepatitis without mention of hepatic coma|Other specified viral hepatitis without mention of hepatic coma
C1456262|T047|PT|070.51|ICD9CM|Acute hepatitis C without mention of hepatic coma|Acute hepatitis C without mention of hepatic coma
C1456262|T047|AB|070.51|ICD9CM|Hpt C acute wo hpat coma|Hpt C acute wo hpat coma
C0375011|T047|PT|070.52|ICD9CM|Hepatitis delta without mention of active hepatitis B disease or hepatic coma|Hepatitis delta without mention of active hepatitis B disease or hepatic coma
C0375011|T047|AB|070.52|ICD9CM|Hpt dlt wo b wo hpt coma|Hpt dlt wo b wo hpt coma
C0153088|T047|PT|070.53|ICD9CM|Hepatitis E without mention of hepatic coma|Hepatitis E without mention of hepatic coma
C0153088|T047|AB|070.53|ICD9CM|Hpt E wo hepat Coma|Hpt E wo hepat Coma
C0375012|T047|AB|070.54|ICD9CM|Chrnc hpt C wo hpat coma|Chrnc hpt C wo hpat coma
C0375012|T047|PT|070.54|ICD9CM|Chronic hepatitis C without mention of hepatic coma|Chronic hepatitis C without mention of hepatic coma
C0153085|T047|AB|070.59|ICD9CM|Oth vrl hpat wo hpt coma|Oth vrl hpat wo hpt coma
C0153085|T047|PT|070.59|ICD9CM|Other specified viral hepatitis without mention of hepatic coma|Other specified viral hepatitis without mention of hepatic coma
C0153089|T047|PT|070.6|ICD9CM|Unspecified viral hepatitis with hepatic coma|Unspecified viral hepatitis with hepatic coma
C0153089|T047|AB|070.6|ICD9CM|Viral hepat NOS w coma|Viral hepat NOS w coma
C0019196|T047|HT|070.7|ICD9CM|Unspecified viral hepatitis C|Unspecified viral hepatitis C
C1456263|T047|AB|070.70|ICD9CM|Hpt C w/o hepat coma NOS|Hpt C w/o hepat coma NOS
C1456263|T047|PT|070.70|ICD9CM|Unspecified viral hepatitis C without hepatic coma|Unspecified viral hepatitis C without hepatic coma
C1456265|T047|AB|070.71|ICD9CM|Hpt C w hepatic coma NOS|Hpt C w hepatic coma NOS
C1456265|T047|PT|070.71|ICD9CM|Unspecified viral hepatitis C with hepatic coma|Unspecified viral hepatitis C with hepatic coma
C0489954|T047|PT|070.9|ICD9CM|Unspecified viral hepatitis without mention of hepatic coma|Unspecified viral hepatitis without mention of hepatic coma
C0489954|T047|AB|070.9|ICD9CM|Viral hepat NOS w/o coma|Viral hepat NOS w/o coma
C0034494|T047|AB|071|ICD9CM|Rabies|Rabies
C0034494|T047|PT|071|ICD9CM|Rabies|Rabies
C0026780|T047|HT|072|ICD9CM|Mumps|Mumps
C0153091|T047|AB|072.0|ICD9CM|Mumps orchitis|Mumps orchitis
C0153091|T047|PT|072.0|ICD9CM|Mumps orchitis|Mumps orchitis
C0153092|T047|AB|072.1|ICD9CM|Mumps meningitis|Mumps meningitis
C0153092|T047|PT|072.1|ICD9CM|Mumps meningitis|Mumps meningitis
C0153093|T047|AB|072.2|ICD9CM|Mumps encephalitis|Mumps encephalitis
C0153093|T047|PT|072.2|ICD9CM|Mumps encephalitis|Mumps encephalitis
C0153094|T047|AB|072.3|ICD9CM|Mumps pancreatitis|Mumps pancreatitis
C0153094|T047|PT|072.3|ICD9CM|Mumps pancreatitis|Mumps pancreatitis
C0153095|T047|HT|072.7|ICD9CM|Mumps with other specified complications|Mumps with other specified complications
C0153096|T047|AB|072.71|ICD9CM|Mumps hepatitis|Mumps hepatitis
C0153096|T047|PT|072.71|ICD9CM|Mumps hepatitis|Mumps hepatitis
C0153097|T047|AB|072.72|ICD9CM|Mumps polyneuropathy|Mumps polyneuropathy
C0153097|T047|PT|072.72|ICD9CM|Mumps polyneuropathy|Mumps polyneuropathy
C0153095|T047|AB|072.79|ICD9CM|Mumps complication NEC|Mumps complication NEC
C0153095|T047|PT|072.79|ICD9CM|Other mumps with other specified complications|Other mumps with other specified complications
C0153098|T047|AB|072.8|ICD9CM|Mumps complication NOS|Mumps complication NOS
C0153098|T047|PT|072.8|ICD9CM|Mumps with unspecified complication|Mumps with unspecified complication
C1306848|T047|AB|072.9|ICD9CM|Mumps uncomplicated|Mumps uncomplicated
C1306848|T047|PT|072.9|ICD9CM|Mumps without mention of complication|Mumps without mention of complication
C0029291|T047|HT|073|ICD9CM|Ornithosis|Ornithosis
C0153099|T047|AB|073.0|ICD9CM|Ornithosis pneumonia|Ornithosis pneumonia
C0153099|T047|PT|073.0|ICD9CM|Ornithosis with pneumonia|Ornithosis with pneumonia
C0153100|T047|AB|073.7|ICD9CM|Ornithosis complicat NEC|Ornithosis complicat NEC
C0153100|T047|PT|073.7|ICD9CM|Ornithosis with other specified complications|Ornithosis with other specified complications
C0153101|T047|AB|073.8|ICD9CM|Ornithosis complicat NOS|Ornithosis complicat NOS
C0153101|T047|PT|073.8|ICD9CM|Ornithosis with unspecified complication|Ornithosis with unspecified complication
C0029291|T047|AB|073.9|ICD9CM|Ornithosis NOS|Ornithosis NOS
C0029291|T047|PT|073.9|ICD9CM|Ornithosis, unspecified|Ornithosis, unspecified
C0728910|T047|HT|074|ICD9CM|Specific diseases due to Coxsackie virus|Specific diseases due to Coxsackie virus
C0019338|T047|AB|074.0|ICD9CM|Herpangina|Herpangina
C0019338|T047|PT|074.0|ICD9CM|Herpangina|Herpangina
C0032238|T047|AB|074.1|ICD9CM|Epidemic pleurodynia|Epidemic pleurodynia
C0032238|T047|PT|074.1|ICD9CM|Epidemic pleurodynia|Epidemic pleurodynia
C0153103|T047|HT|074.2|ICD9CM|Coxsackie carditis|Coxsackie carditis
C0153103|T047|AB|074.20|ICD9CM|Coxsackie carditis NOS|Coxsackie carditis NOS
C0153103|T047|PT|074.20|ICD9CM|Coxsackie carditis, unspecified|Coxsackie carditis, unspecified
C0153104|T047|AB|074.21|ICD9CM|Coxsackie pericarditis|Coxsackie pericarditis
C0153104|T047|PT|074.21|ICD9CM|Coxsackie pericarditis|Coxsackie pericarditis
C0153105|T047|AB|074.22|ICD9CM|Coxsackie endocarditis|Coxsackie endocarditis
C0153105|T047|PT|074.22|ICD9CM|Coxsackie endocarditis|Coxsackie endocarditis
C0153106|T047|AB|074.23|ICD9CM|Coxsackie myocarditis|Coxsackie myocarditis
C0153106|T047|PT|074.23|ICD9CM|Coxsackie myocarditis|Coxsackie myocarditis
C0018572|T047|AB|074.3|ICD9CM|Hand, foot & mouth dis|Hand, foot & mouth dis
C0018572|T047|PT|074.3|ICD9CM|Hand, foot, and mouth disease|Hand, foot, and mouth disease
C0343653|T047|AB|074.8|ICD9CM|Coxsackie virus NEC|Coxsackie virus NEC
C0343653|T047|PT|074.8|ICD9CM|Other specified diseases due to Coxsackie virus|Other specified diseases due to Coxsackie virus
C0021345|T047|AB|075|ICD9CM|Infectious mononucleosis|Infectious mononucleosis
C0021345|T047|PT|075|ICD9CM|Infectious mononucleosis|Infectious mononucleosis
C0040592|T047|HT|076|ICD9CM|Trachoma|Trachoma
C0153107|T047|AB|076.0|ICD9CM|Trachoma, initial stage|Trachoma, initial stage
C0153107|T047|PT|076.0|ICD9CM|Trachoma, initial stage|Trachoma, initial stage
C0153108|T047|AB|076.1|ICD9CM|Trachoma, active stage|Trachoma, active stage
C0153108|T047|PT|076.1|ICD9CM|Trachoma, active stage|Trachoma, active stage
C0040592|T047|AB|076.9|ICD9CM|Trachoma NOS|Trachoma NOS
C0040592|T047|PT|076.9|ICD9CM|Trachoma, unspecified|Trachoma, unspecified
C0153109|T047|HT|077|ICD9CM|Other diseases of conjunctiva due to viruses and Chlamydiae|Other diseases of conjunctiva due to viruses and Chlamydiae
C0009770|T047|AB|077.0|ICD9CM|Inclusion conjunctivitis|Inclusion conjunctivitis
C0009770|T047|PT|077.0|ICD9CM|Inclusion conjunctivitis|Inclusion conjunctivitis
C0014493|T047|AB|077.1|ICD9CM|Epidem keratoconjunctiv|Epidem keratoconjunctiv
C0014493|T047|PT|077.1|ICD9CM|Epidemic keratoconjunctivitis|Epidemic keratoconjunctivitis
C0031351|T047|AB|077.2|ICD9CM|Pharyngoconjunct fever|Pharyngoconjunct fever
C0031351|T047|PT|077.2|ICD9CM|Pharyngoconjunctival fever|Pharyngoconjunctival fever
C0153110|T047|AB|077.3|ICD9CM|Adenoviral conjunct NEC|Adenoviral conjunct NEC
C0153110|T047|PT|077.3|ICD9CM|Other adenoviral conjunctivitis|Other adenoviral conjunctivitis
C0009765|T047|AB|077.4|ICD9CM|Epidem hem conjunctivit|Epidem hem conjunctivit
C0009765|T047|PT|077.4|ICD9CM|Epidemic hemorrhagic conjunctivitis|Epidemic hemorrhagic conjunctivitis
C0029871|T047|PT|077.8|ICD9CM|Other viral conjunctivitis|Other viral conjunctivitis
C0029871|T047|AB|077.8|ICD9CM|Viral conjunctivitis NEC|Viral conjunctivitis NEC
C0041792|T047|HT|077.9|ICD9CM|Unspecified diseases of conjunctiva due to viruses and Chlamydiae|Unspecified diseases of conjunctiva due to viruses and Chlamydiae
C0376110|T047|AB|077.98|ICD9CM|Unsp ds conjuc chlamydia|Unsp ds conjuc chlamydia
C0376110|T047|PT|077.98|ICD9CM|Unspecified diseases of conjunctiva due to chlamydiae|Unspecified diseases of conjunctiva due to chlamydiae
C0376111|T047|AB|077.99|ICD9CM|Unsp ds conjuc viruses|Unsp ds conjuc viruses
C0376111|T047|PT|077.99|ICD9CM|Unspecified diseases of conjunctiva due to viruses|Unspecified diseases of conjunctiva due to viruses
C0153111|T047|HT|078|ICD9CM|Other diseases due to viruses and Chlamydiae|Other diseases due to viruses and Chlamydiae
C0026393|T047|AB|078.0|ICD9CM|Molluscum contagiosum|Molluscum contagiosum
C0026393|T047|PT|078.0|ICD9CM|Molluscum contagiosum|Molluscum contagiosum
C0043037|T047|HT|078.1|ICD9CM|Viral warts|Viral warts
C0343642|T047|AB|078.10|ICD9CM|Viral warts NOS|Viral warts NOS
C0343642|T047|PT|078.10|ICD9CM|Viral warts, unspecified|Viral warts, unspecified
C0009663|T047|AB|078.11|ICD9CM|Condyloma acuminatum|Condyloma acuminatum
C0009663|T047|PT|078.11|ICD9CM|Condyloma acuminatum|Condyloma acuminatum
C0042548|T047|PT|078.12|ICD9CM|Plantar wart|Plantar wart
C0042548|T047|AB|078.12|ICD9CM|Plantar wart|Plantar wart
C0375013|T047|AB|078.19|ICD9CM|Oth specfd viral warts|Oth specfd viral warts
C0375013|T047|PT|078.19|ICD9CM|Other specified viral warts|Other specified viral warts
C0038992|T047|AB|078.2|ICD9CM|Sweating fever|Sweating fever
C0038992|T047|PT|078.2|ICD9CM|Sweating fever|Sweating fever
C0007361|T047|AB|078.3|ICD9CM|Cat-scratch disease|Cat-scratch disease
C0007361|T047|PT|078.3|ICD9CM|Cat-scratch disease|Cat-scratch disease
C0016514|T047|AB|078.4|ICD9CM|Foot & mouth disease|Foot & mouth disease
C0016514|T047|PT|078.4|ICD9CM|Foot and mouth disease|Foot and mouth disease
C0010823|T047|AB|078.5|ICD9CM|Cytomegaloviral disease|Cytomegaloviral disease
C0010823|T047|PT|078.5|ICD9CM|Cytomegaloviral disease|Cytomegaloviral disease
C0019101|T047|AB|078.6|ICD9CM|Hem nephrosonephritis|Hem nephrosonephritis
C0019101|T047|PT|078.6|ICD9CM|Hemorrhagic nephrosonephritis|Hemorrhagic nephrosonephritis
C0153112|T047|AB|078.7|ICD9CM|Arenaviral hem fever|Arenaviral hem fever
C0153112|T047|PT|078.7|ICD9CM|Arenaviral hemorrhagic fever|Arenaviral hemorrhagic fever
C0029767|T047|HT|078.8|ICD9CM|Other specified diseases due to viruses and Chlamydiae|Other specified diseases due to viruses and Chlamydiae
C0751908|T047|AB|078.81|ICD9CM|Epidemic vertigo|Epidemic vertigo
C0751908|T047|PT|078.81|ICD9CM|Epidemic vertigo|Epidemic vertigo
C0014498|T047|AB|078.82|ICD9CM|Epidemic vomiting synd|Epidemic vomiting synd
C0014498|T047|PT|078.82|ICD9CM|Epidemic vomiting syndrome|Epidemic vomiting syndrome
C0375014|T047|AB|078.88|ICD9CM|Oth spec dis chlamydiae|Oth spec dis chlamydiae
C0375014|T047|PT|078.88|ICD9CM|Other specified diseases due to chlamydiae|Other specified diseases due to chlamydiae
C0859831|T047|AB|078.89|ICD9CM|Oth spec dis viruses|Oth spec dis viruses
C0859831|T047|PT|078.89|ICD9CM|Other specified diseases due to viruses|Other specified diseases due to viruses
C0375026|T047|HT|079|ICD9CM|Viral and chlamydial infection in conditions classified elsewhere and of unspecified site|Viral and chlamydial infection in conditions classified elsewhere and of unspecified site
C0001485|T047|AB|079.0|ICD9CM|Adenovirus infect NOS|Adenovirus infect NOS
C0001485|T047|PT|079.0|ICD9CM|Adenovirus infection in conditions classified elsewhere and of unspecified site|Adenovirus infection in conditions classified elsewhere and of unspecified site
C0013515|T047|AB|079.1|ICD9CM|Echo virus infect NOS|Echo virus infect NOS
C0013515|T047|PT|079.1|ICD9CM|Echo virus infection in conditions classified elsewhere and of unspecified site|Echo virus infection in conditions classified elsewhere and of unspecified site
C0010244|T047|AB|079.2|ICD9CM|Coxsackie virus inf NOS|Coxsackie virus inf NOS
C0010244|T047|PT|079.2|ICD9CM|Coxsackie virus infection in conditions classified elsewhere and of unspecified site|Coxsackie virus infection in conditions classified elsewhere and of unspecified site
C0153115|T047|AB|079.3|ICD9CM|Rhinovirus infect NOS|Rhinovirus infect NOS
C0153115|T047|PT|079.3|ICD9CM|Rhinovirus infection in conditions classified elsewhere and of unspecified site|Rhinovirus infection in conditions classified elsewhere and of unspecified site
C0375016|T047|AB|079.4|ICD9CM|Human papillomavirus|Human papillomavirus
C0375016|T047|PT|079.4|ICD9CM|Human papillomavirus in conditions classified elsewhere and of unspecified site|Human papillomavirus in conditions classified elsewhere and of unspecified site
C0375018|T047|HT|079.5|ICD9CM|Retrovirus infection in conditions classified elsewhere and of unspecified site|Retrovirus infection in conditions classified elsewhere and of unspecified site
C0375018|T047|AB|079.50|ICD9CM|Retrovirus, unspecified|Retrovirus, unspecified
C0375018|T047|PT|079.50|ICD9CM|Retrovirus, unspecified|Retrovirus, unspecified
C0375019|T047|AB|079.51|ICD9CM|Htlv-1 infection oth dis|Htlv-1 infection oth dis
C0375019|T047|PT|079.51|ICD9CM|Human T-cell lymphotrophic virus, type I [HTLV-I]|Human T-cell lymphotrophic virus, type I [HTLV-I]
C0375020|T047|AB|079.52|ICD9CM|Htlv-ii infectn oth dis|Htlv-ii infectn oth dis
C0375020|T047|PT|079.52|ICD9CM|Human T-cell lymphotrophic virus, type II [HTLV-II]|Human T-cell lymphotrophic virus, type II [HTLV-II]
C0375021|T047|AB|079.53|ICD9CM|Hiv-2 infection oth dis|Hiv-2 infection oth dis
C0375021|T047|PT|079.53|ICD9CM|Human immunodeficiency virus, type 2 [HIV-2]|Human immunodeficiency virus, type 2 [HIV-2]
C0375022|T047|AB|079.59|ICD9CM|Oth specfied retrovirus|Oth specfied retrovirus
C0375022|T047|PT|079.59|ICD9CM|Other specified retrovirus|Other specified retrovirus
C0375023|T047|PT|079.6|ICD9CM|Respiratory syncytial virus (RSV)|Respiratory syncytial virus (RSV)
C0375023|T047|AB|079.6|ICD9CM|Resprtry syncytial virus|Resprtry syncytial virus
C0375024|T047|AB|079.81|ICD9CM|Hantavirus infection|Hantavirus infection
C0375024|T047|PT|079.81|ICD9CM|Hantavirus infection|Hantavirus infection
C1175175|T047|AB|079.82|ICD9CM|SARS assoc coronavirus|SARS assoc coronavirus
C1175175|T047|PT|079.82|ICD9CM|SARS-associated coronavirus|SARS-associated coronavirus
C1959635|T047|AB|079.83|ICD9CM|Parvovirus B19|Parvovirus B19
C1959635|T047|PT|079.83|ICD9CM|Parvovirus B19|Parvovirus B19
C0375025|T047|AB|079.88|ICD9CM|Oth spcf chlamydial infc|Oth spcf chlamydial infc
C0375025|T047|PT|079.88|ICD9CM|Other specified chlamydial infection|Other specified chlamydial infection
C0029842|T047|AB|079.89|ICD9CM|Oth specf viral infectn|Oth specf viral infectn
C0029842|T047|PT|079.89|ICD9CM|Other specified viral infection|Other specified viral infection
C0375027|T047|AB|079.98|ICD9CM|Chlamydial infection NOS|Chlamydial infection NOS
C0375027|T047|PT|079.98|ICD9CM|Unspecified chlamydial infection|Unspecified chlamydial infection
C0153114|T047|PT|079.99|ICD9CM|Unspecified viral infection|Unspecified viral infection
C0153114|T047|AB|079.99|ICD9CM|Viral infection NOS|Viral infection NOS
C0041473|T047|PT|080|ICD9CM|Louse-borne (epidemic) typhus|Louse-borne (epidemic) typhus
C0041473|T047|AB|080|ICD9CM|Louse-borne typhus|Louse-borne typhus
C0178242|T047|HT|080-088.99|ICD9CM|RICKETTSIOSES AND OTHER ARTHROPOD-BORNE DISEASES|RICKETTSIOSES AND OTHER ARTHROPOD-BORNE DISEASES
C0153116|T047|HT|081|ICD9CM|Other typhus|Other typhus
C0041472|T047|PT|081.0|ICD9CM|Murine (endemic) typhus|Murine (endemic) typhus
C0041472|T047|AB|081.0|ICD9CM|Murine typhus|Murine typhus
C0006181|T047|AB|081.1|ICD9CM|Brill's disease|Brill's disease
C0006181|T047|PT|081.1|ICD9CM|Brill's disease|Brill's disease
C0036472|T047|AB|081.2|ICD9CM|Scrub typhus|Scrub typhus
C0036472|T047|PT|081.2|ICD9CM|Scrub typhus|Scrub typhus
C0041471|T047|AB|081.9|ICD9CM|Typhus NOS|Typhus NOS
C0041471|T047|PT|081.9|ICD9CM|Typhus, unspecified|Typhus, unspecified
C0153117|T047|HT|082|ICD9CM|Tick-borne rickettsioses|Tick-borne rickettsioses
C0038041|T047|AB|082.0|ICD9CM|Spotted fevers|Spotted fevers
C0038041|T047|PT|082.0|ICD9CM|Spotted fevers|Spotted fevers
C0006060|T047|AB|082.1|ICD9CM|Boutonneuse fever|Boutonneuse fever
C0006060|T047|PT|082.1|ICD9CM|Boutonneuse fever|Boutonneuse fever
C0549160|T047|PT|082.2|ICD9CM|North Asian tick fever|North Asian tick fever
C0549160|T047|AB|082.2|ICD9CM|North asian tick fever|North asian tick fever
C2979888|T047|AB|082.3|ICD9CM|Queensland tick typhus|Queensland tick typhus
C2979888|T047|PT|082.3|ICD9CM|Queensland tick typhus|Queensland tick typhus
C0085399|T047|HT|082.4|ICD9CM|Ehrlichiosis|Ehrlichiosis
C0085399|T047|AB|082.40|ICD9CM|Ehrlichiosis NOS|Ehrlichiosis NOS
C0085399|T047|PT|082.40|ICD9CM|Ehrlichiosis, unspecified|Ehrlichiosis, unspecified
C1282983|T047|AB|082.41|ICD9CM|Ehrlichiosis chafeensis|Ehrlichiosis chafeensis
C1282983|T047|PT|082.41|ICD9CM|Ehrlichiosis chafeensis [E. chafeensis]|Ehrlichiosis chafeensis [E. chafeensis]
C0878688|T047|AB|082.49|ICD9CM|Ehrlichiosis NEC|Ehrlichiosis NEC
C0878688|T047|PT|082.49|ICD9CM|Other ehrlichiosis|Other ehrlichiosis
C0153118|T047|PT|082.8|ICD9CM|Other specified tick-borne rickettsioses|Other specified tick-borne rickettsioses
C0153118|T047|AB|082.8|ICD9CM|Tick-borne ricketts NEC|Tick-borne ricketts NEC
C0153117|T047|AB|082.9|ICD9CM|Tick-borne ricketts NOS|Tick-borne ricketts NOS
C0153117|T047|PT|082.9|ICD9CM|Tick-borne rickettsiosis, unspecified|Tick-borne rickettsiosis, unspecified
C0153119|T047|HT|083|ICD9CM|Other rickettsioses|Other rickettsioses
C0034362|T047|AB|083.0|ICD9CM|Q fever|Q fever
C0034362|T047|PT|083.0|ICD9CM|Q fever|Q fever
C0040830|T047|AB|083.1|ICD9CM|Trench fever|Trench fever
C0040830|T047|PT|083.1|ICD9CM|Trench fever|Trench fever
C0035597|T047|AB|083.2|ICD9CM|Rickettsialpox|Rickettsialpox
C0035597|T047|PT|083.2|ICD9CM|Rickettsialpox|Rickettsialpox
C0153120|T047|PT|083.8|ICD9CM|Other specified rickettsioses|Other specified rickettsioses
C0153120|T047|AB|083.8|ICD9CM|Rickettsioses NEC|Rickettsioses NEC
C0035585|T047|AB|083.9|ICD9CM|Rickettsiosis NOS|Rickettsiosis NOS
C0035585|T047|PT|083.9|ICD9CM|Rickettsiosis, unspecified|Rickettsiosis, unspecified
C0024530|T047|HT|084|ICD9CM|Malaria|Malaria
C0024535|T047|AB|084.0|ICD9CM|Falciparum malaria|Falciparum malaria
C0024535|T047|PT|084.0|ICD9CM|Falciparum malaria [malignant tertian]|Falciparum malaria [malignant tertian]
C0024537|T047|AB|084.1|ICD9CM|Vivax malaria|Vivax malaria
C0024537|T047|PT|084.1|ICD9CM|Vivax malaria [benign tertian]|Vivax malaria [benign tertian]
C0024536|T047|AB|084.2|ICD9CM|Quartan malaria|Quartan malaria
C0024536|T047|PT|084.2|ICD9CM|Quartan malaria|Quartan malaria
C0152072|T047|AB|084.3|ICD9CM|Ovale malaria|Ovale malaria
C0152072|T047|PT|084.3|ICD9CM|Ovale malaria|Ovale malaria
C0029661|T047|AB|084.4|ICD9CM|Malaria NEC|Malaria NEC
C0029661|T047|PT|084.4|ICD9CM|Other malaria|Other malaria
C0153121|T047|AB|084.5|ICD9CM|Mixed malaria|Mixed malaria
C0153121|T047|PT|084.5|ICD9CM|Mixed malaria|Mixed malaria
C0024530|T047|AB|084.6|ICD9CM|Malaria NOS|Malaria NOS
C0024530|T047|PT|084.6|ICD9CM|Malaria, unspecified|Malaria, unspecified
C0153122|T047|AB|084.7|ICD9CM|Induced malaria|Induced malaria
C0153122|T047|PT|084.7|ICD9CM|Induced malaria|Induced malaria
C0005681|T047|AB|084.8|ICD9CM|Blackwater fever|Blackwater fever
C0005681|T047|PT|084.8|ICD9CM|Blackwater fever|Blackwater fever
C0153123|T047|AB|084.9|ICD9CM|Malaria complicated NEC|Malaria complicated NEC
C0153123|T047|PT|084.9|ICD9CM|Other pernicious complications of malaria|Other pernicious complications of malaria
C0023281|T047|HT|085|ICD9CM|Leishmaniasis|Leishmaniasis
C0023290|T047|PT|085.0|ICD9CM|Visceral [kala-azar] leishmaniasis|Visceral [kala-azar] leishmaniasis
C0023290|T047|AB|085.0|ICD9CM|Visceral leishmaniasis|Visceral leishmaniasis
C0086541|T047|AB|085.1|ICD9CM|Cutan leishmanias urban|Cutan leishmanias urban
C0086541|T047|PT|085.1|ICD9CM|Cutaneous leishmaniasis, urban|Cutaneous leishmaniasis, urban
C0023285|T047|AB|085.2|ICD9CM|Cutan leishmanias asian|Cutan leishmanias asian
C0023285|T047|PT|085.2|ICD9CM|Cutaneous leishmaniasis, Asian desert|Cutaneous leishmaniasis, Asian desert
C0152074|T047|AB|085.3|ICD9CM|Cutan leishmanias ethiop|Cutan leishmanias ethiop
C0152074|T047|PT|085.3|ICD9CM|Cutaneous leishmaniasis, Ethiopian|Cutaneous leishmaniasis, Ethiopian
C3495436|T047|AB|085.4|ICD9CM|Cutan leishmanias amer|Cutan leishmanias amer
C3495436|T047|PT|085.4|ICD9CM|Cutaneous leishmaniasis, American|Cutaneous leishmaniasis, American
C1328252|T047|AB|085.5|ICD9CM|Mucocutan leishmaniasis|Mucocutan leishmaniasis
C1328252|T047|PT|085.5|ICD9CM|Mucocutaneous leishmaniasis, (American)|Mucocutaneous leishmaniasis, (American)
C0023281|T047|AB|085.9|ICD9CM|Leishmaniasis NOS|Leishmaniasis NOS
C0023281|T047|PT|085.9|ICD9CM|Leishmaniasis, unspecified|Leishmaniasis, unspecified
C0041227|T047|HT|086|ICD9CM|Trypanosomiasis|Trypanosomiasis
C0007930|T047|AB|086.0|ICD9CM|Chagas disease of heart|Chagas disease of heart
C0007930|T047|PT|086.0|ICD9CM|Chagas' disease with heart involvement|Chagas' disease with heart involvement
C0153125|T047|AB|086.1|ICD9CM|Chagas dis of oth organ|Chagas dis of oth organ
C0153125|T047|PT|086.1|ICD9CM|Chagas' disease with other organ involvement|Chagas' disease with other organ involvement
C0007932|T047|AB|086.2|ICD9CM|Chagas disease NOS|Chagas disease NOS
C0007932|T047|PT|086.2|ICD9CM|Chagas' disease without mention of organ involvement|Chagas' disease without mention of organ involvement
C0041232|T047|AB|086.3|ICD9CM|Gambian trypanosomiasis|Gambian trypanosomiasis
C0041232|T047|PT|086.3|ICD9CM|Gambian trypanosomiasis|Gambian trypanosomiasis
C0041233|T047|AB|086.4|ICD9CM|Rhodesian trypanosomias|Rhodesian trypanosomias
C0041233|T047|PT|086.4|ICD9CM|Rhodesian trypanosomiasis|Rhodesian trypanosomiasis
C0041228|T047|AB|086.5|ICD9CM|African trypanosoma NOS|African trypanosoma NOS
C0041228|T047|PT|086.5|ICD9CM|African trypanosomiasis, unspecified|African trypanosomiasis, unspecified
C0041227|T047|AB|086.9|ICD9CM|Trypanosomiasis NOS|Trypanosomiasis NOS
C0041227|T047|PT|086.9|ICD9CM|Trypanosomiasis, unspecified|Trypanosomiasis, unspecified
C0035021|T047|HT|087|ICD9CM|Relapsing fever|Relapsing fever
C0152061|T047|AB|087.0|ICD9CM|Louse-borne relaps fever|Louse-borne relaps fever
C0152061|T047|PT|087.0|ICD9CM|Relapsing fever, louse-borne|Relapsing fever, louse-borne
C0035022|T047|PT|087.1|ICD9CM|Relapsing fever, tick-borne|Relapsing fever, tick-borne
C0035022|T047|AB|087.1|ICD9CM|Tick-borne relaps fever|Tick-borne relaps fever
C0035021|T047|AB|087.9|ICD9CM|Relapsing fever NOS|Relapsing fever NOS
C0035021|T047|PT|087.9|ICD9CM|Relapsing fever, unspecified|Relapsing fever, unspecified
C0153126|T047|HT|088|ICD9CM|Other arthropod-borne diseases|Other arthropod-borne diseases
C0004771|T047|AB|088.0|ICD9CM|Bartonellosis|Bartonellosis
C0004771|T047|PT|088.0|ICD9CM|Bartonellosis|Bartonellosis
C0029747|T047|HT|088.8|ICD9CM|Other specified arthropod-borne diseases|Other specified arthropod-borne diseases
C0024198|T047|PT|088.81|ICD9CM|Lyme Disease|Lyme Disease
C0024198|T047|AB|088.81|ICD9CM|Lyme disease|Lyme disease
C0004576|T047|AB|088.82|ICD9CM|Babesiosis|Babesiosis
C0004576|T047|PT|088.82|ICD9CM|Babesiosis|Babesiosis
C0029747|T047|AB|088.89|ICD9CM|Oth arthropod-borne dis|Oth arthropod-borne dis
C0029747|T047|PT|088.89|ICD9CM|Other specified arthropod-borne diseases, other|Other specified arthropod-borne diseases, other
C0521829|T047|AB|088.9|ICD9CM|Arthropod-borne dis NOS|Arthropod-borne dis NOS
C0521829|T047|PT|088.9|ICD9CM|Arthropod-borne disease, unspecified|Arthropod-borne disease, unspecified
C0039131|T047|HT|090|ICD9CM|Congenital syphilis|Congenital syphilis
C0178243|T047|HT|090-099.99|ICD9CM|SYPHILIS AND OTHER VENEREAL DISEASES|SYPHILIS AND OTHER VENEREAL DISEASES
C0343666|T047|AB|090.0|ICD9CM|Early cong syph symptom|Early cong syph symptom
C0343666|T047|PT|090.0|ICD9CM|Early congenital syphilis, symptomatic|Early congenital syphilis, symptomatic
C0153129|T047|AB|090.1|ICD9CM|Early congen syph latent|Early congen syph latent
C0153129|T047|PT|090.1|ICD9CM|Early congenital syphilis, latent|Early congenital syphilis, latent
C0275859|T019|AB|090.2|ICD9CM|Early congen syph NOS|Early congen syph NOS
C0275859|T047|AB|090.2|ICD9CM|Early congen syph NOS|Early congen syph NOS
C0275859|T019|PT|090.2|ICD9CM|Early congenital syphilis, unspecified|Early congenital syphilis, unspecified
C0275859|T047|PT|090.2|ICD9CM|Early congenital syphilis, unspecified|Early congenital syphilis, unspecified
C2039668|T019|PT|090.3|ICD9CM|Syphilitic interstitial keratitis|Syphilitic interstitial keratitis
C2039668|T047|PT|090.3|ICD9CM|Syphilitic interstitial keratitis|Syphilitic interstitial keratitis
C2039668|T019|AB|090.3|ICD9CM|Syphilitic keratitis|Syphilitic keratitis
C2039668|T047|AB|090.3|ICD9CM|Syphilitic keratitis|Syphilitic keratitis
C0153132|T047|HT|090.4|ICD9CM|Juvenile neurosyphilis|Juvenile neurosyphilis
C0153132|T047|AB|090.40|ICD9CM|Juvenile neurosyph NOS|Juvenile neurosyph NOS
C0153132|T047|PT|090.40|ICD9CM|Juvenile neurosyphilis, unspecified|Juvenile neurosyphilis, unspecified
C0153133|T047|AB|090.41|ICD9CM|Congen syph encephalitis|Congen syph encephalitis
C0153133|T047|PT|090.41|ICD9CM|Congenital syphilitic encephalitis|Congenital syphilitic encephalitis
C0153134|T047|AB|090.42|ICD9CM|Congen syph meningitis|Congen syph meningitis
C0153134|T047|PT|090.42|ICD9CM|Congenital syphilitic meningitis|Congenital syphilitic meningitis
C0153135|T047|AB|090.49|ICD9CM|Juvenile neurosyph NEC|Juvenile neurosyph NEC
C0153135|T047|PT|090.49|ICD9CM|Other juvenile neurosyphilis|Other juvenile neurosyphilis
C0153136|T047|AB|090.5|ICD9CM|Late congen syph symptom|Late congen syph symptom
C0153136|T047|PT|090.5|ICD9CM|Other late congenital syphilis, symptomatic|Other late congenital syphilis, symptomatic
C0275874|T047|AB|090.6|ICD9CM|Late congen syph latent|Late congen syph latent
C0275874|T047|PT|090.6|ICD9CM|Late congenital syphilis, latent|Late congenital syphilis, latent
C0554634|T047|AB|090.7|ICD9CM|Late congen syph NOS|Late congen syph NOS
C0554634|T047|PT|090.7|ICD9CM|Late congenital syphilis, unspecified|Late congenital syphilis, unspecified
C0039131|T047|AB|090.9|ICD9CM|Congenital syphilis NOS|Congenital syphilis NOS
C0039131|T047|PT|090.9|ICD9CM|Congenital syphilis, unspecified|Congenital syphilis, unspecified
C0153139|T047|HT|091|ICD9CM|Early syphilis, symptomatic|Early syphilis, symptomatic
C0017418|T047|PT|091.0|ICD9CM|Genital syphilis (primary)|Genital syphilis (primary)
C0017418|T047|AB|091.0|ICD9CM|Primary genital syphilis|Primary genital syphilis
C0153140|T047|AB|091.1|ICD9CM|Primary anal syphilis|Primary anal syphilis
C0153140|T047|PT|091.1|ICD9CM|Primary anal syphilis|Primary anal syphilis
C0153141|T047|PT|091.2|ICD9CM|Other primary syphilis|Other primary syphilis
C0153141|T047|AB|091.2|ICD9CM|Primary syphilis NEC|Primary syphilis NEC
C0343677|T047|AB|091.3|ICD9CM|Secondary syph skin|Secondary syph skin
C0343677|T047|PT|091.3|ICD9CM|Secondary syphilis of skin or mucous membranes|Secondary syphilis of skin or mucous membranes
C0275834|T047|PT|091.4|ICD9CM|Adenopathy due to secondary syphilis|Adenopathy due to secondary syphilis
C0275834|T047|AB|091.4|ICD9CM|Syphilitic adenopathy|Syphilitic adenopathy
C0275836|T047|HT|091.5|ICD9CM|Uveitis due to secondary syphilis|Uveitis due to secondary syphilis
C0275836|T047|AB|091.50|ICD9CM|Syphilitic uveitis NOS|Syphilitic uveitis NOS
C0275836|T047|PT|091.50|ICD9CM|Syphilitic uveitis, unspecified|Syphilitic uveitis, unspecified
C0153145|T047|AB|091.51|ICD9CM|Syphilit chorioretinitis|Syphilit chorioretinitis
C0153145|T047|PT|091.51|ICD9CM|Syphilitic chorioretinitis (secondary)|Syphilitic chorioretinitis (secondary)
C0153146|T047|AB|091.52|ICD9CM|Syphilitic iridocyclitis|Syphilitic iridocyclitis
C0153146|T047|PT|091.52|ICD9CM|Syphilitic iridocyclitis (secondary)|Syphilitic iridocyclitis (secondary)
C0343676|T047|HT|091.6|ICD9CM|Secondary syphilis of viscera and bone|Secondary syphilis of viscera and bone
C0153148|T047|PT|091.61|ICD9CM|Secondary syphilitic periostitis|Secondary syphilitic periostitis
C0153148|T047|AB|091.61|ICD9CM|Syphilitic periostitis|Syphilitic periostitis
C0153149|T047|PT|091.62|ICD9CM|Secondary syphilitic hepatitis|Secondary syphilitic hepatitis
C0153149|T047|AB|091.62|ICD9CM|Syphilitic hepatitis|Syphilitic hepatitis
C0153150|T047|AB|091.69|ICD9CM|Second syph viscera NEC|Second syph viscera NEC
C0153150|T047|PT|091.69|ICD9CM|Secondary syphilis of other viscera|Secondary syphilis of other viscera
C0153151|T047|AB|091.7|ICD9CM|Second syphilis relapse|Second syphilis relapse
C0153151|T047|PT|091.7|ICD9CM|Secondary syphilis, relapse|Secondary syphilis, relapse
C0348147|T047|HT|091.8|ICD9CM|Other forms of secondary syphilis|Other forms of secondary syphilis
C0851315|T047|AB|091.81|ICD9CM|Acute syphil meningitis|Acute syphil meningitis
C0851315|T047|PT|091.81|ICD9CM|Acute syphilitic meningitis (secondary)|Acute syphilitic meningitis (secondary)
C0002181|T047|AB|091.82|ICD9CM|Syphilitic alopecia|Syphilitic alopecia
C0002181|T047|PT|091.82|ICD9CM|Syphilitic alopecia|Syphilitic alopecia
C0348147|T047|PT|091.89|ICD9CM|Other forms of secondary syphilis|Other forms of secondary syphilis
C0348147|T047|AB|091.89|ICD9CM|Secondary syphilis NEC|Secondary syphilis NEC
C0149985|T047|AB|091.9|ICD9CM|Secondary syphilis NOS|Secondary syphilis NOS
C0149985|T047|PT|091.9|ICD9CM|Unspecified secondary syphilis|Unspecified secondary syphilis
C0275842|T047|HT|092|ICD9CM|Early syphilis, latent|Early syphilis, latent
C0153156|T047|AB|092.0|ICD9CM|Early syph latent relaps|Early syph latent relaps
C0153156|T047|PT|092.0|ICD9CM|Early syphilis, latent, serological relapse after treatment|Early syphilis, latent, serological relapse after treatment
C0275842|T047|AB|092.9|ICD9CM|Early syphil latent NOS|Early syphil latent NOS
C0275842|T047|PT|092.9|ICD9CM|Early syphilis, latent, unspecified|Early syphilis, latent, unspecified
C0039130|T047|HT|093|ICD9CM|Cardiovascular syphilis|Cardiovascular syphilis
C0275844|T047|PT|093.0|ICD9CM|Aneurysm of aorta, specified as syphilitic|Aneurysm of aorta, specified as syphilitic
C0275844|T047|AB|093.0|ICD9CM|Aortic aneurysm, syphil|Aortic aneurysm, syphil
C0003511|T047|AB|093.1|ICD9CM|Syphilitic aortitis|Syphilitic aortitis
C0003511|T047|PT|093.1|ICD9CM|Syphilitic aortitis|Syphilitic aortitis
C0153158|T047|HT|093.2|ICD9CM|Syphilitic endocarditis|Syphilitic endocarditis
C0340334|T047|AB|093.20|ICD9CM|Syphil endocarditis NOS|Syphil endocarditis NOS
C0340334|T047|PT|093.20|ICD9CM|Syphilitic endocarditis of valve, unspecified|Syphilitic endocarditis of valve, unspecified
C0153160|T047|PT|093.21|ICD9CM|Syphilitic endocarditis of mitral valve|Syphilitic endocarditis of mitral valve
C0153160|T047|AB|093.21|ICD9CM|Syphilitic mitral valve|Syphilitic mitral valve
C0153161|T047|AB|093.22|ICD9CM|Syphilitic aortic valve|Syphilitic aortic valve
C0153161|T047|PT|093.22|ICD9CM|Syphilitic endocarditis of aortic valve|Syphilitic endocarditis of aortic valve
C0153162|T047|AB|093.23|ICD9CM|Syphil tricuspid valve|Syphil tricuspid valve
C0153162|T047|PT|093.23|ICD9CM|Syphilitic endocarditis of tricuspid valve|Syphilitic endocarditis of tricuspid valve
C0153163|T047|AB|093.24|ICD9CM|Syphil pulmonary valve|Syphil pulmonary valve
C0153163|T047|PT|093.24|ICD9CM|Syphilitic endocarditis of pulmonary valve|Syphilitic endocarditis of pulmonary valve
C0029751|T047|HT|093.8|ICD9CM|Other specified cardiovascular syphilis|Other specified cardiovascular syphilis
C0153164|T047|AB|093.81|ICD9CM|Syphilitic pericarditis|Syphilitic pericarditis
C0153164|T047|PT|093.81|ICD9CM|Syphilitic pericarditis|Syphilitic pericarditis
C0153165|T047|AB|093.82|ICD9CM|Syphilitic myocarditis|Syphilitic myocarditis
C0153165|T047|PT|093.82|ICD9CM|Syphilitic myocarditis|Syphilitic myocarditis
C0029751|T047|AB|093.89|ICD9CM|Cardiovascular syph NEC|Cardiovascular syph NEC
C0029751|T047|PT|093.89|ICD9CM|Other specified cardiovascular syphilis|Other specified cardiovascular syphilis
C0039130|T047|AB|093.9|ICD9CM|Cardiovascular syph NOS|Cardiovascular syph NOS
C0039130|T047|PT|093.9|ICD9CM|Cardiovascular syphilis, unspecified|Cardiovascular syphilis, unspecified
C0027927|T047|HT|094|ICD9CM|Neurosyphilis|Neurosyphilis
C0039223|T047|AB|094.0|ICD9CM|Tabes dorsalis|Tabes dorsalis
C0039223|T047|PT|094.0|ICD9CM|Tabes dorsalis|Tabes dorsalis
C0205858|T047|AB|094.1|ICD9CM|General paresis|General paresis
C0205858|T047|PT|094.1|ICD9CM|General paresis|General paresis
C0153166|T047|AB|094.2|ICD9CM|Syphilitic meningitis|Syphilitic meningitis
C0153166|T047|PT|094.2|ICD9CM|Syphilitic meningitis|Syphilitic meningitis
C0153167|T047|AB|094.3|ICD9CM|Asymptomat neurosyphilis|Asymptomat neurosyphilis
C0153167|T047|PT|094.3|ICD9CM|Asymptomatic neurosyphilis|Asymptomatic neurosyphilis
C0029817|T047|HT|094.8|ICD9CM|Other specified neurosyphilis|Other specified neurosyphilis
C0153168|T047|AB|094.81|ICD9CM|Syphilitic encephalitis|Syphilitic encephalitis
C0153168|T047|PT|094.81|ICD9CM|Syphilitic encephalitis|Syphilitic encephalitis
C0153169|T047|AB|094.82|ICD9CM|Syphilitic parkinsonism|Syphilitic parkinsonism
C0153169|T047|PT|094.82|ICD9CM|Syphilitic parkinsonism|Syphilitic parkinsonism
C0153170|T047|AB|094.83|ICD9CM|Syph dissem retinitis|Syph dissem retinitis
C0153170|T047|PT|094.83|ICD9CM|Syphilitic disseminated retinochoroiditis|Syphilitic disseminated retinochoroiditis
C0153171|T047|AB|094.84|ICD9CM|Syphilitic optic atrophy|Syphilitic optic atrophy
C0153171|T047|PT|094.84|ICD9CM|Syphilitic optic atrophy|Syphilitic optic atrophy
C0153172|T047|AB|094.85|ICD9CM|Syph retrobulb neuritis|Syph retrobulb neuritis
C0153172|T047|PT|094.85|ICD9CM|Syphilitic retrobulbar neuritis|Syphilitic retrobulbar neuritis
C0153173|T047|AB|094.86|ICD9CM|Syphil acoustic neuritis|Syphil acoustic neuritis
C0153173|T047|PT|094.86|ICD9CM|Syphilitic acoustic neuritis|Syphilitic acoustic neuritis
C0153174|T047|AB|094.87|ICD9CM|Syph rupt cereb aneurysm|Syph rupt cereb aneurysm
C0153174|T047|PT|094.87|ICD9CM|Syphilitic ruptured cerebral aneurysm|Syphilitic ruptured cerebral aneurysm
C0029817|T047|AB|094.89|ICD9CM|Neurosyphilis NEC|Neurosyphilis NEC
C0029817|T047|PT|094.89|ICD9CM|Other specified neurosyphilis|Other specified neurosyphilis
C0027927|T047|AB|094.9|ICD9CM|Neurosyphilis NOS|Neurosyphilis NOS
C0027927|T047|PT|094.9|ICD9CM|Neurosyphilis, unspecified|Neurosyphilis, unspecified
C0348149|T047|HT|095|ICD9CM|Other forms of late syphilis, with symptoms|Other forms of late syphilis, with symptoms
C0153176|T047|AB|095.0|ICD9CM|Syphilitic episcleritis|Syphilitic episcleritis
C0153176|T047|PT|095.0|ICD9CM|Syphilitic episcleritis|Syphilitic episcleritis
C0153177|T047|AB|095.1|ICD9CM|Syphilis of lung|Syphilis of lung
C0153177|T047|PT|095.1|ICD9CM|Syphilis of lung|Syphilis of lung
C0153178|T047|AB|095.2|ICD9CM|Syphilitic peritonitis|Syphilitic peritonitis
C0153178|T047|PT|095.2|ICD9CM|Syphilitic peritonitis|Syphilitic peritonitis
C0153179|T047|AB|095.3|ICD9CM|Syphilis of liver|Syphilis of liver
C0153179|T047|PT|095.3|ICD9CM|Syphilis of liver|Syphilis of liver
C0153180|T047|AB|095.4|ICD9CM|Syphilis of kidney|Syphilis of kidney
C0153180|T047|PT|095.4|ICD9CM|Syphilis of kidney|Syphilis of kidney
C0153181|T047|AB|095.5|ICD9CM|Syphilis of bone|Syphilis of bone
C0153181|T047|PT|095.5|ICD9CM|Syphilis of bone|Syphilis of bone
C0153182|T047|AB|095.6|ICD9CM|Syphilis of muscle|Syphilis of muscle
C0153182|T047|PT|095.6|ICD9CM|Syphilis of muscle|Syphilis of muscle
C0153183|T047|PT|095.7|ICD9CM|Syphilis of synovium, tendon, and bursa|Syphilis of synovium, tendon, and bursa
C0153183|T047|AB|095.7|ICD9CM|Syphilis of tendon/bursa|Syphilis of tendon/bursa
C0343689|T047|AB|095.8|ICD9CM|Late sympt syphilis NEC|Late sympt syphilis NEC
C0343689|T047|PT|095.8|ICD9CM|Other specified forms of late symptomatic syphilis|Other specified forms of late symptomatic syphilis
C0153185|T047|AB|095.9|ICD9CM|Late sympt syphilis NOS|Late sympt syphilis NOS
C0153185|T047|PT|095.9|ICD9CM|Late symptomatic syphilis, unspecified|Late symptomatic syphilis, unspecified
C1260915|T047|AB|096|ICD9CM|Late syphilis latent|Late syphilis latent
C1260915|T047|PT|096|ICD9CM|Late syphilis, latent|Late syphilis, latent
C0558995|T047|HT|097|ICD9CM|Other and unspecified syphilis|Other and unspecified syphilis
C0153188|T047|AB|097.0|ICD9CM|Late syphilis NOS|Late syphilis NOS
C0153188|T047|PT|097.0|ICD9CM|Late syphilis, unspecified|Late syphilis, unspecified
C0039133|T047|AB|097.1|ICD9CM|Latent syphilis NOS|Latent syphilis NOS
C0039133|T047|PT|097.1|ICD9CM|Latent syphilis, unspecified|Latent syphilis, unspecified
C0039128|T047|AB|097.9|ICD9CM|Syphilis NOS|Syphilis NOS
C0039128|T047|PT|097.9|ICD9CM|Syphilis, unspecified|Syphilis, unspecified
C0018081|T047|HT|098|ICD9CM|Gonococcal infections|Gonococcal infections
C0018074|T047|AB|098.0|ICD9CM|Acute gc infect lower gu|Acute gc infect lower gu
C0018074|T047|PT|098.0|ICD9CM|Gonococcal infection (acute) of lower genitourinary tract|Gonococcal infection (acute) of lower genitourinary tract
C0375028|T047|HT|098.1|ICD9CM|Gonococcal infection (acute) of upper genitourinary tract|Gonococcal infection (acute) of upper genitourinary tract
C0375028|T047|AB|098.10|ICD9CM|Gc (acute) upper gu NOS|Gc (acute) upper gu NOS
C0375028|T047|PT|098.10|ICD9CM|Gonococcal infection (acute) of upper genitourinary tract, site unspecified|Gonococcal infection (acute) of upper genitourinary tract, site unspecified
C0153191|T047|AB|098.11|ICD9CM|Gc cystitis (acute)|Gc cystitis (acute)
C0153191|T047|PT|098.11|ICD9CM|Gonococcal cystitis (acute)|Gonococcal cystitis (acute)
C0153192|T047|AB|098.12|ICD9CM|Gc prostatitis (acute)|Gc prostatitis (acute)
C0153192|T047|PT|098.12|ICD9CM|Gonococcal prostatitis (acute)|Gonococcal prostatitis (acute)
C0153193|T047|AB|098.13|ICD9CM|Gc orchitis (acute)|Gc orchitis (acute)
C0153193|T047|PT|098.13|ICD9CM|Gonococcal epididymo-orchitis (acute)|Gonococcal epididymo-orchitis (acute)
C0153194|T047|AB|098.14|ICD9CM|Gc sem vesiculit (acute)|Gc sem vesiculit (acute)
C0153194|T047|PT|098.14|ICD9CM|Gonococcal seminal vesiculitis (acute)|Gonococcal seminal vesiculitis (acute)
C0153195|T047|AB|098.15|ICD9CM|Gc cervicitis (acute)|Gc cervicitis (acute)
C0153195|T047|PT|098.15|ICD9CM|Gonococcal cervicitis (acute)|Gonococcal cervicitis (acute)
C0153196|T047|AB|098.16|ICD9CM|Gc endometritis (acute)|Gc endometritis (acute)
C0153196|T047|PT|098.16|ICD9CM|Gonococcal endometritis (acute)|Gonococcal endometritis (acute)
C0275654|T047|AB|098.17|ICD9CM|Acute gc salpingitis|Acute gc salpingitis
C0275654|T047|PT|098.17|ICD9CM|Gonococcal salpingitis, specified as acute|Gonococcal salpingitis, specified as acute
C0153198|T047|AB|098.19|ICD9CM|Gc (acute) upper gu NEC|Gc (acute) upper gu NEC
C0153198|T047|PT|098.19|ICD9CM|Other gonococcal infection (acute) of upper genitourinary tract|Other gonococcal infection (acute) of upper genitourinary tract
C0153199|T047|AB|098.2|ICD9CM|Chr gc infect lower gu|Chr gc infect lower gu
C0153199|T047|PT|098.2|ICD9CM|Gonococcal infection, chronic, of lower genitourinary tract|Gonococcal infection, chronic, of lower genitourinary tract
C0375029|T047|HT|098.3|ICD9CM|Gonococcal infection, chronic, of upper genitourinary tract|Gonococcal infection, chronic, of upper genitourinary tract
C0375029|T047|AB|098.30|ICD9CM|Chr gc upper gu NOS|Chr gc upper gu NOS
C0375029|T047|PT|098.30|ICD9CM|Chronic gonococcal infection of upper genitourinary tract, site unspecified|Chronic gonococcal infection of upper genitourinary tract, site unspecified
C0153202|T047|AB|098.31|ICD9CM|Gc cystitis, chronic|Gc cystitis, chronic
C0153202|T047|PT|098.31|ICD9CM|Gonococcal cystitis, chronic|Gonococcal cystitis, chronic
C0153203|T047|AB|098.32|ICD9CM|Gc prostatitis, chronic|Gc prostatitis, chronic
C0153203|T047|PT|098.32|ICD9CM|Gonococcal prostatitis, chronic|Gonococcal prostatitis, chronic
C0153204|T047|AB|098.33|ICD9CM|Gc orchitis, chronic|Gc orchitis, chronic
C0153204|T047|PT|098.33|ICD9CM|Gonococcal epididymo-orchitis, chronic|Gonococcal epididymo-orchitis, chronic
C0153205|T047|AB|098.34|ICD9CM|Gc sem vesiculitis, chr|Gc sem vesiculitis, chr
C0153205|T047|PT|098.34|ICD9CM|Gonococcal seminal vesiculitis, chronic|Gonococcal seminal vesiculitis, chronic
C0153206|T047|AB|098.35|ICD9CM|Gc cervicitis, chronic|Gc cervicitis, chronic
C0153206|T047|PT|098.35|ICD9CM|Gonococcal cervicitis, chronic|Gonococcal cervicitis, chronic
C0153207|T047|AB|098.36|ICD9CM|Gc endometritis, chronic|Gc endometritis, chronic
C0153207|T047|PT|098.36|ICD9CM|Gonococcal endometritis, chronic|Gonococcal endometritis, chronic
C0153208|T047|AB|098.37|ICD9CM|Gc salpingitis (chronic)|Gc salpingitis (chronic)
C0153208|T047|PT|098.37|ICD9CM|Gonococcal salpingitis (chronic)|Gonococcal salpingitis (chronic)
C0153209|T047|AB|098.39|ICD9CM|Chr gc upper gu NEC|Chr gc upper gu NEC
C0153209|T047|PT|098.39|ICD9CM|Other chronic gonococcal infection of upper genitourinary tract|Other chronic gonococcal infection of upper genitourinary tract
C0153210|T047|HT|098.4|ICD9CM|Gonococcal infection of eye|Gonococcal infection of eye
C0339166|T047|AB|098.40|ICD9CM|Gonococcal conjunctivit|Gonococcal conjunctivit
C0339166|T047|PT|098.40|ICD9CM|Gonococcal conjunctivitis (neonatorum)|Gonococcal conjunctivitis (neonatorum)
C0153212|T047|AB|098.41|ICD9CM|Gonococcal iridocyclitis|Gonococcal iridocyclitis
C0153212|T047|PT|098.41|ICD9CM|Gonococcal iridocyclitis|Gonococcal iridocyclitis
C0153213|T047|AB|098.42|ICD9CM|Gonococcal endophthalmia|Gonococcal endophthalmia
C0153213|T047|PT|098.42|ICD9CM|Gonococcal endophthalmia|Gonococcal endophthalmia
C0153214|T047|AB|098.43|ICD9CM|Gonococcal keratitis|Gonococcal keratitis
C0153214|T047|PT|098.43|ICD9CM|Gonococcal keratitis|Gonococcal keratitis
C0153215|T047|AB|098.49|ICD9CM|Gonococcal eye NEC|Gonococcal eye NEC
C0153215|T047|PT|098.49|ICD9CM|Other gonococcal infection of eye|Other gonococcal infection of eye
C0153216|T047|HT|098.5|ICD9CM|Gonococcal infection of joint|Gonococcal infection of joint
C0153216|T047|AB|098.50|ICD9CM|Gonococcal arthritis|Gonococcal arthritis
C0153216|T047|PT|098.50|ICD9CM|Gonococcal arthritis|Gonococcal arthritis
C0343714|T047|AB|098.51|ICD9CM|Gonococcal synovitis|Gonococcal synovitis
C0343714|T047|PT|098.51|ICD9CM|Gonococcal synovitis and tenosynovitis|Gonococcal synovitis and tenosynovitis
C0153218|T047|AB|098.52|ICD9CM|Gonococcal bursitis|Gonococcal bursitis
C0153218|T047|PT|098.52|ICD9CM|Gonococcal bursitis|Gonococcal bursitis
C0153219|T047|AB|098.53|ICD9CM|Gonococcal spondylitis|Gonococcal spondylitis
C0153219|T047|PT|098.53|ICD9CM|Gonococcal spondylitis|Gonococcal spondylitis
C0153220|T047|AB|098.59|ICD9CM|Gc infect joint NEC|Gc infect joint NEC
C0153220|T047|PT|098.59|ICD9CM|Other gonococcal infection of joint|Other gonococcal infection of joint
C0149966|T047|AB|098.6|ICD9CM|Gonococcal infec pharynx|Gonococcal infec pharynx
C0149966|T047|PT|098.6|ICD9CM|Gonococcal infection of pharynx|Gonococcal infection of pharynx
C0153222|T047|AB|098.7|ICD9CM|Gc infect anus & rectum|Gc infect anus & rectum
C0153222|T047|PT|098.7|ICD9CM|Gonococcal infection of anus and rectum|Gonococcal infection of anus and rectum
C0153223|T047|HT|098.8|ICD9CM|Gonococcal infection of other specified sites|Gonococcal infection of other specified sites
C0018075|T047|AB|098.81|ICD9CM|Gonococcal keratosis|Gonococcal keratosis
C0018075|T047|PT|098.81|ICD9CM|Gonococcal keratosis (blennorrhagica)|Gonococcal keratosis (blennorrhagica)
C0153225|T047|AB|098.82|ICD9CM|Gonococcal meningitis|Gonococcal meningitis
C0153225|T047|PT|098.82|ICD9CM|Gonococcal meningitis|Gonococcal meningitis
C0153226|T047|AB|098.83|ICD9CM|Gonococcal pericarditis|Gonococcal pericarditis
C0153226|T047|PT|098.83|ICD9CM|Gonococcal pericarditis|Gonococcal pericarditis
C0153227|T047|AB|098.84|ICD9CM|Gonococcal endocarditis|Gonococcal endocarditis
C0153227|T047|PT|098.84|ICD9CM|Gonococcal endocarditis|Gonococcal endocarditis
C0153228|T047|AB|098.85|ICD9CM|Gonococcal heart dis NEC|Gonococcal heart dis NEC
C0153228|T047|PT|098.85|ICD9CM|Other gonococcal heart disease|Other gonococcal heart disease
C0018077|T047|AB|098.86|ICD9CM|Gonococcal peritonitis|Gonococcal peritonitis
C0018077|T047|PT|098.86|ICD9CM|Gonococcal peritonitis|Gonococcal peritonitis
C0153223|T047|AB|098.89|ICD9CM|Gonococcal inf site NEC|Gonococcal inf site NEC
C0153223|T047|PT|098.89|ICD9CM|Gonococcal infection of other specified sites|Gonococcal infection of other specified sites
C0153229|T047|HT|099|ICD9CM|Other venereal diseases|Other venereal diseases
C0007947|T047|AB|099.0|ICD9CM|Chancroid|Chancroid
C0007947|T047|PT|099.0|ICD9CM|Chancroid|Chancroid
C0024286|T047|AB|099.1|ICD9CM|Lymphogranuloma venereum|Lymphogranuloma venereum
C0024286|T047|PT|099.1|ICD9CM|Lymphogranuloma venereum|Lymphogranuloma venereum
C0018190|T047|AB|099.2|ICD9CM|Granuloma inguinale|Granuloma inguinale
C0018190|T047|PT|099.2|ICD9CM|Granuloma inguinale|Granuloma inguinale
C0035012|T047|AB|099.3|ICD9CM|Reiter's disease|Reiter's disease
C0035012|T047|PT|099.3|ICD9CM|Reiter's disease|Reiter's disease
C1112700|T047|HT|099.4|ICD9CM|Other nongonococcal urethritis [NGU]|Other nongonococcal urethritis [NGU]
C0375031|T047|PT|099.40|ICD9CM|Other nongonococcal urethritis, unspecified|Other nongonococcal urethritis, unspecified
C0375031|T047|AB|099.40|ICD9CM|Unspcf nongnccl urethrts|Unspcf nongnccl urethrts
C1278807|T047|AB|099.41|ICD9CM|Chlmyd trachomatis ureth|Chlmyd trachomatis ureth
C1278807|T047|PT|099.41|ICD9CM|Other nongonococcal urethritis, chlamydia trachomatis|Other nongonococcal urethritis, chlamydia trachomatis
C0375033|T047|AB|099.49|ICD9CM|Nongc urth oth spf orgsm|Nongc urth oth spf orgsm
C0375033|T047|PT|099.49|ICD9CM|Other nongonococcal urethritis, other specified organism|Other nongonococcal urethritis, other specified organism
C0375034|T047|HT|099.5|ICD9CM|Other venereal diseases due to Chlamydia trachomatis|Other venereal diseases due to Chlamydia trachomatis
C0375035|T047|AB|099.50|ICD9CM|Oth VD chlm trch unsp st|Oth VD chlm trch unsp st
C0375035|T047|PT|099.50|ICD9CM|Other venereal diseases due to chlamydia trachomatis, unspecified site|Other venereal diseases due to chlamydia trachomatis, unspecified site
C0375036|T047|AB|099.51|ICD9CM|Oth VD chlm trch pharynx|Oth VD chlm trch pharynx
C0375036|T047|PT|099.51|ICD9CM|Other venereal diseases due to chlamydia trachomatis, pharynx|Other venereal diseases due to chlamydia trachomatis, pharynx
C0348903|T047|AB|099.52|ICD9CM|Oth VD chlm trch ans rct|Oth VD chlm trch ans rct
C0348903|T047|PT|099.52|ICD9CM|Other venereal diseases due to chlamydia trachomatis, anus and rectum|Other venereal diseases due to chlamydia trachomatis, anus and rectum
C0348904|T047|AB|099.53|ICD9CM|Oth VD chlm trch lowr gu|Oth VD chlm trch lowr gu
C0348904|T047|PT|099.53|ICD9CM|Other venereal diseases due to chlamydia trachomatis, lower genitourinary sites|Other venereal diseases due to chlamydia trachomatis, lower genitourinary sites
C0375039|T047|AB|099.54|ICD9CM|Oth VD chlm trch oth gu|Oth VD chlm trch oth gu
C0375039|T047|PT|099.54|ICD9CM|Other venereal diseases due to chlamydia trachomatis, other genitourinary sites|Other venereal diseases due to chlamydia trachomatis, other genitourinary sites
C0348157|T047|AB|099.55|ICD9CM|Ot VD chlm trch unspf gu|Ot VD chlm trch unspf gu
C0348157|T047|PT|099.55|ICD9CM|Other venereal diseases due to chlamydia trachomatis, unspecified genitourinary site|Other venereal diseases due to chlamydia trachomatis, unspecified genitourinary site
C0375041|T047|AB|099.56|ICD9CM|Ot VD chlm trch prtoneum|Ot VD chlm trch prtoneum
C0375041|T047|PT|099.56|ICD9CM|Other venereal diseases due to chlamydia trachomatis, peritoneum|Other venereal diseases due to chlamydia trachomatis, peritoneum
C0375042|T047|AB|099.59|ICD9CM|Oth VD chlm trch spcf st|Oth VD chlm trch spcf st
C0375042|T047|PT|099.59|ICD9CM|Other venereal diseases due to chlamydia trachomatis, other specified site|Other venereal diseases due to chlamydia trachomatis, other specified site
C0029840|T047|PT|099.8|ICD9CM|Other specified venereal diseases|Other specified venereal diseases
C0029840|T047|AB|099.8|ICD9CM|Venereal disease NEC|Venereal disease NEC
C0036916|T047|AB|099.9|ICD9CM|Venereal disease NOS|Venereal disease NOS
C0036916|T047|PT|099.9|ICD9CM|Venereal disease, unspecified|Venereal disease, unspecified
C0023364|T047|HT|100|ICD9CM|Leptospirosis|Leptospirosis
C0178244|T047|HT|100-104.99|ICD9CM|OTHER SPIROCHETAL DISEASES|OTHER SPIROCHETAL DISEASES
C0043102|T047|AB|100.0|ICD9CM|Leptospiros icterohem|Leptospiros icterohem
C0043102|T047|PT|100.0|ICD9CM|Leptospirosis icterohemorrhagica|Leptospirosis icterohemorrhagica
C0153231|T047|HT|100.8|ICD9CM|Other specified leptospiral infections|Other specified leptospiral infections
C0153232|T047|AB|100.81|ICD9CM|Leptospiral meningitis|Leptospiral meningitis
C0153232|T047|PT|100.81|ICD9CM|Leptospiral meningitis (aseptic)|Leptospiral meningitis (aseptic)
C0153231|T047|AB|100.89|ICD9CM|Leptospiral infect NEC|Leptospiral infect NEC
C0153231|T047|PT|100.89|ICD9CM|Other specified leptospiral infections|Other specified leptospiral infections
C0023364|T047|AB|100.9|ICD9CM|Leptospirosis NOS|Leptospirosis NOS
C0023364|T047|PT|100.9|ICD9CM|Leptospirosis, unspecified|Leptospirosis, unspecified
C1527368|T047|AB|101|ICD9CM|Vincent's angina|Vincent's angina
C1527368|T047|PT|101|ICD9CM|Vincent's angina|Vincent's angina
C0043388|T047|HT|102|ICD9CM|Yaws|Yaws
C0275990|T047|PT|102.0|ICD9CM|Initial lesions of yaws|Initial lesions of yaws
C0275990|T047|AB|102.0|ICD9CM|Initial lesions yaws|Initial lesions yaws
C0153234|T047|AB|102.1|ICD9CM|Multiple papillomata|Multiple papillomata
C0153234|T047|PT|102.1|ICD9CM|Multiple papillomata due to yaws and wet crab yaws|Multiple papillomata due to yaws and wet crab yaws
C0153235|T047|AB|102.2|ICD9CM|Early skin yaws NEC|Early skin yaws NEC
C0153235|T047|PT|102.2|ICD9CM|Other early skin lesions of yaws|Other early skin lesions of yaws
C0276001|T047|PT|102.3|ICD9CM|Hyperkeratosis due to yaws|Hyperkeratosis due to yaws
C0276001|T047|AB|102.3|ICD9CM|Hyperkeratosis of yaws|Hyperkeratosis of yaws
C0276007|T047|PT|102.4|ICD9CM|Gummata and ulcers due to yaws|Gummata and ulcers due to yaws
C0276007|T047|AB|102.4|ICD9CM|Gummata and ulcers, yaws|Gummata and ulcers, yaws
C0276009|T047|AB|102.5|ICD9CM|Gangosa|Gangosa
C0276009|T047|PT|102.5|ICD9CM|Gangosa|Gangosa
C0343834|T047|PT|102.6|ICD9CM|Bone and joint lesions due to yaws|Bone and joint lesions due to yaws
C0343834|T047|AB|102.6|ICD9CM|Yaws of bone & joint|Yaws of bone & joint
C0153239|T047|PT|102.7|ICD9CM|Other manifestations of yaws|Other manifestations of yaws
C0153239|T047|AB|102.7|ICD9CM|Yaws manifestations NEC|Yaws manifestations NEC
C0153240|T047|AB|102.8|ICD9CM|Latent yaws|Latent yaws
C0153240|T047|PT|102.8|ICD9CM|Latent yaws|Latent yaws
C0043388|T047|AB|102.9|ICD9CM|Yaws NOS|Yaws NOS
C0043388|T047|PT|102.9|ICD9CM|Yaws, unspecified|Yaws, unspecified
C0031946|T047|HT|103|ICD9CM|Pinta|Pinta
C0153241|T047|AB|103.0|ICD9CM|Pinta primary lesions|Pinta primary lesions
C0153241|T047|PT|103.0|ICD9CM|Primary lesions of pinta|Primary lesions of pinta
C0153242|T047|PT|103.1|ICD9CM|Intermediate lesions of pinta|Intermediate lesions of pinta
C0153242|T047|AB|103.1|ICD9CM|Pinta intermed lesions|Pinta intermed lesions
C0153243|T047|PT|103.2|ICD9CM|Late lesions of pinta|Late lesions of pinta
C0153243|T047|AB|103.2|ICD9CM|Pinta late lesions|Pinta late lesions
C0153244|T047|PT|103.3|ICD9CM|Mixed lesions of pinta|Mixed lesions of pinta
C0153244|T047|AB|103.3|ICD9CM|Pinta mixed lesions|Pinta mixed lesions
C0031946|T047|AB|103.9|ICD9CM|Pinta NOS|Pinta NOS
C0031946|T047|PT|103.9|ICD9CM|Pinta, unspecified|Pinta, unspecified
C0153245|T047|HT|104|ICD9CM|Other spirochetal infection|Other spirochetal infection
C3537179|T047|AB|104.0|ICD9CM|Nonvenereal endemic syph|Nonvenereal endemic syph
C3537179|T047|PT|104.0|ICD9CM|Nonvenereal endemic syphilis|Nonvenereal endemic syphilis
C0029830|T047|PT|104.8|ICD9CM|Other specified spirochetal infections|Other specified spirochetal infections
C0029830|T047|AB|104.8|ICD9CM|Spirochetal infect NEC|Spirochetal infect NEC
C0037974|T047|AB|104.9|ICD9CM|Spirochetal infect NOS|Spirochetal infect NOS
C0037974|T047|PT|104.9|ICD9CM|Spirochetal infection, unspecified|Spirochetal infection, unspecified
C0011636|T047|HT|110|ICD9CM|Dermatophytosis|Dermatophytosis
C0026946|T047|HT|110-118.99|ICD9CM|MYCOSES|MYCOSES
C0011640|T047|AB|110.0|ICD9CM|Dermatophyt scalp/beard|Dermatophyt scalp/beard
C0011640|T047|PT|110.0|ICD9CM|Dermatophytosis of scalp and beard|Dermatophytosis of scalp and beard
C4082762|T047|AB|110.1|ICD9CM|Dermatophytosis of nail|Dermatophytosis of nail
C4082762|T047|PT|110.1|ICD9CM|Dermatophytosis of nail|Dermatophytosis of nail
C0153246|T047|AB|110.2|ICD9CM|Dermatophytosis of hand|Dermatophytosis of hand
C0153246|T047|PT|110.2|ICD9CM|Dermatophytosis of hand|Dermatophytosis of hand
C0011638|T047|AB|110.3|ICD9CM|Dermatophytosis of groin|Dermatophytosis of groin
C0011638|T047|PT|110.3|ICD9CM|Dermatophytosis of groin and perianal area|Dermatophytosis of groin and perianal area
C0040259|T047|AB|110.4|ICD9CM|Dermatophytosis of foot|Dermatophytosis of foot
C0040259|T047|PT|110.4|ICD9CM|Dermatophytosis of foot|Dermatophytosis of foot
C0546826|T047|AB|110.5|ICD9CM|Dermatophytosis of body|Dermatophytosis of body
C0546826|T047|PT|110.5|ICD9CM|Dermatophytosis of the body|Dermatophytosis of the body
C1395264|T047|AB|110.6|ICD9CM|Deep dermatophytosis|Deep dermatophytosis
C1395264|T047|PT|110.6|ICD9CM|Deep seated dermatophytosis|Deep seated dermatophytosis
C0153248|T047|PT|110.8|ICD9CM|Dermatophytosis of other specified sites|Dermatophytosis of other specified sites
C0153248|T047|AB|110.8|ICD9CM|Dermatophytosis site NEC|Dermatophytosis site NEC
C0011636|T047|PT|110.9|ICD9CM|Dermatophytosis of unspecified site|Dermatophytosis of unspecified site
C0011636|T047|AB|110.9|ICD9CM|Dermatophytosis site NOS|Dermatophytosis site NOS
C0011630|T047|HT|111|ICD9CM|Dermatomycosis, other and unspecified|Dermatomycosis, other and unspecified
C0040262|T047|AB|111.0|ICD9CM|Pityriasis versicolor|Pityriasis versicolor
C0040262|T047|PT|111.0|ICD9CM|Pityriasis versicolor|Pityriasis versicolor
C0152067|T047|AB|111.1|ICD9CM|Tinea nigra|Tinea nigra
C0152067|T047|PT|111.1|ICD9CM|Tinea nigra|Tinea nigra
C0040249|T047|AB|111.2|ICD9CM|Tinea blanca|Tinea blanca
C0040249|T047|PT|111.2|ICD9CM|Tinea blanca|Tinea blanca
C0153249|T047|AB|111.3|ICD9CM|Black piedra|Black piedra
C0153249|T047|PT|111.3|ICD9CM|Black piedra|Black piedra
C0029763|T047|AB|111.8|ICD9CM|Dermatomycoses NEC|Dermatomycoses NEC
C0029763|T047|PT|111.8|ICD9CM|Other specified dermatomycoses|Other specified dermatomycoses
C0011630|T047|AB|111.9|ICD9CM|Dermatomycosis NOS|Dermatomycosis NOS
C0011630|T047|PT|111.9|ICD9CM|Dermatomycosis, unspecified|Dermatomycosis, unspecified
C0006840|T047|HT|112|ICD9CM|Candidiasis|Candidiasis
C0006849|T047|PT|112.0|ICD9CM|Candidiasis of mouth|Candidiasis of mouth
C0006849|T047|AB|112.0|ICD9CM|Thrush|Thrush
C0700345|T047|AB|112.1|ICD9CM|Candidal vulvovaginitis|Candidal vulvovaginitis
C0700345|T047|PT|112.1|ICD9CM|Candidiasis of vulva and vagina|Candidiasis of vulva and vagina
C0153250|T047|AB|112.2|ICD9CM|Candidias urogenital NEC|Candidias urogenital NEC
C0153250|T047|PT|112.2|ICD9CM|Candidiasis of other urogenital sites|Candidiasis of other urogenital sites
C0006842|T047|PT|112.3|ICD9CM|Candidiasis of skin and nails|Candidiasis of skin and nails
C0006842|T047|AB|112.3|ICD9CM|Cutaneous candidiasis|Cutaneous candidiasis
C0153251|T047|AB|112.4|ICD9CM|Candidiasis of lung|Candidiasis of lung
C0153251|T047|PT|112.4|ICD9CM|Candidiasis of lung|Candidiasis of lung
C0153252|T047|AB|112.5|ICD9CM|Disseminated candidiasis|Disseminated candidiasis
C0153252|T047|PT|112.5|ICD9CM|Disseminated candidiasis|Disseminated candidiasis
C0153253|T047|HT|112.8|ICD9CM|Candidiasis of other specified sites|Candidiasis of other specified sites
C0153254|T047|AB|112.81|ICD9CM|Candidal endocarditis|Candidal endocarditis
C0153254|T047|PT|112.81|ICD9CM|Candidal endocarditis|Candidal endocarditis
C0153255|T047|AB|112.82|ICD9CM|Candidal otitis externa|Candidal otitis externa
C0153255|T047|PT|112.82|ICD9CM|Candidal otitis externa|Candidal otitis externa
C0153256|T047|AB|112.83|ICD9CM|Candidal meningitis|Candidal meningitis
C0153256|T047|PT|112.83|ICD9CM|Candidal meningitis|Candidal meningitis
C0239295|T047|AB|112.84|ICD9CM|Candidal esophagitis|Candidal esophagitis
C0239295|T047|PT|112.84|ICD9CM|Candidal esophagitis|Candidal esophagitis
C0858895|T047|AB|112.85|ICD9CM|Candidal enteritis|Candidal enteritis
C0858895|T047|PT|112.85|ICD9CM|Candidal enteritis|Candidal enteritis
C3665466|T047|AB|112.89|ICD9CM|Candidiasis site NEC|Candidiasis site NEC
C3665466|T047|PT|112.89|ICD9CM|Other candidiasis of other specified sites|Other candidiasis of other specified sites
C0006840|T047|PT|112.9|ICD9CM|Candidiasis of unspecified site|Candidiasis of unspecified site
C0006840|T047|AB|112.9|ICD9CM|Candidiasis site NOS|Candidiasis site NOS
C0009186|T047|HT|114|ICD9CM|Coccidioidomycosis|Coccidioidomycosis
C0153257|T047|AB|114.0|ICD9CM|Primary coccidioidomycos|Primary coccidioidomycos
C0153257|T047|PT|114.0|ICD9CM|Primary coccidioidomycosis (pulmonary)|Primary coccidioidomycosis (pulmonary)
C0700644|T047|AB|114.1|ICD9CM|Prim cutan coccidioid|Prim cutan coccidioid
C0700644|T047|PT|114.1|ICD9CM|Primary extrapulmonary coccidioidomycosis|Primary extrapulmonary coccidioidomycosis
C0153259|T047|AB|114.2|ICD9CM|Coccidioidal meningitis|Coccidioidal meningitis
C0153259|T047|PT|114.2|ICD9CM|Coccidioidal meningitis|Coccidioidal meningitis
C0343891|T047|PT|114.3|ICD9CM|Other forms of progressive coccidioidomycosis|Other forms of progressive coccidioidomycosis
C0343891|T047|AB|114.3|ICD9CM|Progress coccidioid NEC|Progress coccidioid NEC
C0339963|T047|AB|114.4|ICD9CM|Ch pl coccidioidomycosis|Ch pl coccidioidomycosis
C0339963|T047|PT|114.4|ICD9CM|Chronic pulmonary coccidioidomycosis|Chronic pulmonary coccidioidomycosis
C0375046|T047|AB|114.5|ICD9CM|Pl cocidioidomycosis NOS|Pl cocidioidomycosis NOS
C0375046|T047|PT|114.5|ICD9CM|Pulmonary coccidioidomycosis, unspecified|Pulmonary coccidioidomycosis, unspecified
C0009186|T047|AB|114.9|ICD9CM|Coccidioidomycosis NOS|Coccidioidomycosis NOS
C0009186|T047|PT|114.9|ICD9CM|Coccidioidomycosis, unspecified|Coccidioidomycosis, unspecified
C0019655|T047|HT|115|ICD9CM|Histoplasmosis|Histoplasmosis
C0153261|T047|HT|115.0|ICD9CM|Infection by Histoplasma capsulatum|Infection by Histoplasma capsulatum
C0153262|T047|AB|115.00|ICD9CM|Histoplasma capsulat NOS|Histoplasma capsulat NOS
C0153262|T047|PT|115.00|ICD9CM|Infection by Histoplasma capsulatum, without mention of manifestation|Infection by Histoplasma capsulatum, without mention of manifestation
C0153263|T047|AB|115.01|ICD9CM|Histoplasm capsul mening|Histoplasm capsul mening
C0153263|T047|PT|115.01|ICD9CM|Infection by Histoplasma capsulatum, meningitis|Infection by Histoplasma capsulatum, meningitis
C0153264|T047|AB|115.02|ICD9CM|Histoplasm capsul retina|Histoplasm capsul retina
C0153264|T047|PT|115.02|ICD9CM|Infection by Histoplasma capsulatum, retinitis|Infection by Histoplasma capsulatum, retinitis
C0153265|T047|AB|115.03|ICD9CM|Histoplasm caps pericard|Histoplasm caps pericard
C0153265|T047|PT|115.03|ICD9CM|Infection by Histoplasma capsulatum, pericarditis|Infection by Histoplasma capsulatum, pericarditis
C0153266|T047|AB|115.04|ICD9CM|Histoplasm caps endocard|Histoplasm caps endocard
C0153266|T047|PT|115.04|ICD9CM|Infection by Histoplasma capsulatum, endocarditis|Infection by Histoplasma capsulatum, endocarditis
C1261318|T047|AB|115.05|ICD9CM|Histoplasm caps pneumon|Histoplasm caps pneumon
C1261318|T047|PT|115.05|ICD9CM|Infection by Histoplasma capsulatum, pneumonia|Infection by Histoplasma capsulatum, pneumonia
C0153268|T047|AB|115.09|ICD9CM|Histoplasma capsulat NEC|Histoplasma capsulat NEC
C0153268|T047|PT|115.09|ICD9CM|Infection by Histoplasma capsulatum, other|Infection by Histoplasma capsulatum, other
C0220977|T047|HT|115.1|ICD9CM|Infection by Histoplasma duboisii|Infection by Histoplasma duboisii
C0153270|T047|AB|115.10|ICD9CM|Histoplasma duboisii NOS|Histoplasma duboisii NOS
C0153270|T047|PT|115.10|ICD9CM|Infection by Histoplasma duboisii, without mention of manifestation|Infection by Histoplasma duboisii, without mention of manifestation
C0153271|T047|AB|115.11|ICD9CM|Histoplasm dubois mening|Histoplasm dubois mening
C0153271|T047|PT|115.11|ICD9CM|Infection by Histoplasma duboisii, meningitis|Infection by Histoplasma duboisii, meningitis
C0153272|T047|AB|115.12|ICD9CM|Histoplasm dubois retina|Histoplasm dubois retina
C0153272|T047|PT|115.12|ICD9CM|Infection by Histoplasma duboisii, retinitis|Infection by Histoplasma duboisii, retinitis
C0153273|T047|AB|115.13|ICD9CM|Histoplasm dub pericard|Histoplasm dub pericard
C0153273|T047|PT|115.13|ICD9CM|Infection by Histoplasma duboisii, pericarditis|Infection by Histoplasma duboisii, pericarditis
C0153274|T047|AB|115.14|ICD9CM|Histoplasm dub endocard|Histoplasm dub endocard
C0153274|T047|PT|115.14|ICD9CM|Infection by Histoplasma duboisii, endocarditis|Infection by Histoplasma duboisii, endocarditis
C0153275|T047|AB|115.15|ICD9CM|Histoplasm dub pneumonia|Histoplasm dub pneumonia
C0153275|T047|PT|115.15|ICD9CM|Infection by Histoplasma duboisii, pneumonia|Infection by Histoplasma duboisii, pneumonia
C0153276|T047|AB|115.19|ICD9CM|Histoplasma duboisii NEC|Histoplasma duboisii NEC
C0153276|T047|PT|115.19|ICD9CM|Infection by Histoplasma duboisii, other|Infection by Histoplasma duboisii, other
C0019655|T047|HT|115.9|ICD9CM|Histoplasmosis, unspecified|Histoplasmosis, unspecified
C0677640|T047|AB|115.90|ICD9CM|Histoplasmosis NOS|Histoplasmosis NOS
C0677640|T047|PT|115.90|ICD9CM|Histoplasmosis, unspecified, without mention of manifestation|Histoplasmosis, unspecified, without mention of manifestation
C0153277|T047|AB|115.91|ICD9CM|Histoplasmosis meningit|Histoplasmosis meningit
C0153277|T047|PT|115.91|ICD9CM|Histoplasmosis, unspecified, meningitis|Histoplasmosis, unspecified, meningitis
C0153278|T047|AB|115.92|ICD9CM|Histoplasmosis retinitis|Histoplasmosis retinitis
C0153278|T047|PT|115.92|ICD9CM|Histoplasmosis, unspecified, retinitis|Histoplasmosis, unspecified, retinitis
C0153279|T047|AB|115.93|ICD9CM|Histoplasmosis pericard|Histoplasmosis pericard
C0153279|T047|PT|115.93|ICD9CM|Histoplasmosis, unspecified, pericarditis|Histoplasmosis, unspecified, pericarditis
C0153266|T047|AB|115.94|ICD9CM|Histoplasmosis endocard|Histoplasmosis endocard
C0153266|T047|PT|115.94|ICD9CM|Histoplasmosis, unspecified, endocarditis|Histoplasmosis, unspecified, endocarditis
C0153281|T047|AB|115.95|ICD9CM|Histoplasmosis pneumonia|Histoplasmosis pneumonia
C0153281|T047|PT|115.95|ICD9CM|Histoplasmosis, unspecified, pneumonia|Histoplasmosis, unspecified, pneumonia
C0019657|T047|AB|115.99|ICD9CM|Histoplasmosis NEC|Histoplasmosis NEC
C0019657|T047|PT|115.99|ICD9CM|Histoplasmosis, unspecified, other|Histoplasmosis, unspecified, other
C0005716|T047|HT|116|ICD9CM|Blastomycotic infection|Blastomycotic infection
C0005716|T047|AB|116.0|ICD9CM|Blastomycosis|Blastomycosis
C0005716|T047|PT|116.0|ICD9CM|Blastomycosis|Blastomycosis
C0030409|T047|AB|116.1|ICD9CM|Paracoccidioidomycosis|Paracoccidioidomycosis
C0030409|T047|PT|116.1|ICD9CM|Paracoccidioidomycosis|Paracoccidioidomycosis
C0152066|T047|AB|116.2|ICD9CM|Lobomycosis|Lobomycosis
C0152066|T047|PT|116.2|ICD9CM|Lobomycosis|Lobomycosis
C0343846|T047|HT|117|ICD9CM|Other mycoses|Other mycoses
C0035469|T047|AB|117.0|ICD9CM|Rhinosporidiosis|Rhinosporidiosis
C0035469|T047|PT|117.0|ICD9CM|Rhinosporidiosis|Rhinosporidiosis
C0038034|T047|AB|117.1|ICD9CM|Sporotrichosis|Sporotrichosis
C0038034|T047|PT|117.1|ICD9CM|Sporotrichosis|Sporotrichosis
C0008582|T047|AB|117.2|ICD9CM|Chromoblastomycosis|Chromoblastomycosis
C0008582|T047|PT|117.2|ICD9CM|Chromoblastomycosis|Chromoblastomycosis
C0004030|T047|AB|117.3|ICD9CM|Aspergillosis|Aspergillosis
C0004030|T047|PT|117.3|ICD9CM|Aspergillosis|Aspergillosis
C2350621|T047|AB|117.4|ICD9CM|Mycotic mycetomas|Mycotic mycetomas
C2350621|T047|PT|117.4|ICD9CM|Mycotic mycetomas|Mycotic mycetomas
C0010414|T047|AB|117.5|ICD9CM|Cryptococcosis|Cryptococcosis
C0010414|T047|PT|117.5|ICD9CM|Cryptococcosis|Cryptococcosis
C0153285|T047|AB|117.6|ICD9CM|Allescheriosis|Allescheriosis
C0153285|T047|PT|117.6|ICD9CM|Allescheriosis [Petriellidosis]|Allescheriosis [Petriellidosis]
C0043541|T047|AB|117.7|ICD9CM|Zygomycosis|Zygomycosis
C0043541|T047|PT|117.7|ICD9CM|Zygomycosis [Phycomycosis or Mucormycosis]|Zygomycosis [Phycomycosis or Mucormycosis]
C0276721|T047|AB|117.8|ICD9CM|Dematiacious fungi inf|Dematiacious fungi inf
C0276721|T047|PT|117.8|ICD9CM|Infection by dematiacious fungi [Phaehyphomycosis]|Infection by dematiacious fungi [Phaehyphomycosis]
C0029511|T047|AB|117.9|ICD9CM|Mycoses NEC & NOS|Mycoses NEC & NOS
C0029511|T047|PT|117.9|ICD9CM|Other and unspecified mycoses|Other and unspecified mycoses
C0029119|T047|AB|118|ICD9CM|Opportunistic mycoses|Opportunistic mycoses
C0029119|T047|PT|118|ICD9CM|Opportunistic mycoses|Opportunistic mycoses
C0036323|T047|HT|120|ICD9CM|Schistosomiasis [bilharziasis]|Schistosomiasis [bilharziasis]
C0018889|T047|HT|120-129.99|ICD9CM|HELMINTHIASES|HELMINTHIASES
C0276926|T047|AB|120.0|ICD9CM|Schistosoma haematobium|Schistosoma haematobium
C0276926|T047|PT|120.0|ICD9CM|Schistosomiasis due to schistosoma haematobium|Schistosomiasis due to schistosoma haematobium
C0036330|T047|AB|120.1|ICD9CM|Schistosoma mansoni|Schistosoma mansoni
C0036330|T047|PT|120.1|ICD9CM|Schistosomiasis due to schistosoma mansoni|Schistosomiasis due to schistosoma mansoni
C0036329|T047|AB|120.2|ICD9CM|Schistosoma japonicum|Schistosoma japonicum
C0036329|T047|PT|120.2|ICD9CM|Schistosomiasis due to schistosoma japonicum|Schistosomiasis due to schistosoma japonicum
C0546996|T047|AB|120.3|ICD9CM|Cutaneous schistosoma|Cutaneous schistosoma
C0546996|T047|PT|120.3|ICD9CM|Cutaneous schistosomiasis|Cutaneous schistosomiasis
C0029827|T047|PT|120.8|ICD9CM|Other specified schistosomiasis|Other specified schistosomiasis
C0029827|T047|AB|120.8|ICD9CM|Schistosomiasis NEC|Schistosomiasis NEC
C0036323|T047|AB|120.9|ICD9CM|Schistosomiasis NOS|Schistosomiasis NOS
C0036323|T047|PT|120.9|ICD9CM|Schistosomiasis, unspecified|Schistosomiasis, unspecified
C0153288|T047|HT|121|ICD9CM|Other trematode infections|Other trematode infections
C0029106|T047|AB|121.0|ICD9CM|Opisthorchiasis|Opisthorchiasis
C0029106|T047|PT|121.0|ICD9CM|Opisthorchiasis|Opisthorchiasis
C0009021|T047|AB|121.1|ICD9CM|Clonorchiasis|Clonorchiasis
C0009021|T047|PT|121.1|ICD9CM|Clonorchiasis|Clonorchiasis
C0030424|T047|AB|121.2|ICD9CM|Paragonimiasis|Paragonimiasis
C0030424|T047|PT|121.2|ICD9CM|Paragonimiasis|Paragonimiasis
C0015652|T047|AB|121.3|ICD9CM|Fascioliasis|Fascioliasis
C0015652|T047|PT|121.3|ICD9CM|Fascioliasis|Fascioliasis
C0015656|T047|AB|121.4|ICD9CM|Fasciolopsiasis|Fasciolopsiasis
C0015656|T047|PT|121.4|ICD9CM|Fasciolopsiasis|Fasciolopsiasis
C0025530|T047|AB|121.5|ICD9CM|Metagonimiasis|Metagonimiasis
C0025530|T047|PT|121.5|ICD9CM|Metagonimiasis|Metagonimiasis
C0152071|T047|AB|121.6|ICD9CM|Heterophyiasis|Heterophyiasis
C0152071|T047|PT|121.6|ICD9CM|Heterophyiasis|Heterophyiasis
C0029833|T047|PT|121.8|ICD9CM|Other specified trematode infections|Other specified trematode infections
C0029833|T047|AB|121.8|ICD9CM|Trematode infection NEC|Trematode infection NEC
C0040820|T047|AB|121.9|ICD9CM|Trematode infection NOS|Trematode infection NOS
C0040820|T047|PT|121.9|ICD9CM|Trematode infection, unspecified|Trematode infection, unspecified
C0013502|T047|HT|122|ICD9CM|Echinococcosis|Echinococcosis
C0153289|T047|AB|122.0|ICD9CM|Echinococc granul liver|Echinococc granul liver
C0153289|T047|PT|122.0|ICD9CM|Echinococcus granulosus infection of liver|Echinococcus granulosus infection of liver
C0153290|T047|AB|122.1|ICD9CM|Echinococc granul lung|Echinococc granul lung
C0153290|T047|PT|122.1|ICD9CM|Echinococcus granulosus infection of lung|Echinococcus granulosus infection of lung
C0153291|T047|AB|122.2|ICD9CM|Echinococc gran thyroid|Echinococc gran thyroid
C0153291|T047|PT|122.2|ICD9CM|Echinococcus granulosus infection of thyroid|Echinococcus granulosus infection of thyroid
C0153292|T047|AB|122.3|ICD9CM|Echinococc granul NEC|Echinococc granul NEC
C0153292|T047|PT|122.3|ICD9CM|Echinococcus granulosus infection, other|Echinococcus granulosus infection, other
C0152068|T047|AB|122.4|ICD9CM|Echinococc granul NOS|Echinococc granul NOS
C0152068|T047|PT|122.4|ICD9CM|Echinococcus granulosus infection, unspecified|Echinococcus granulosus infection, unspecified
C0153293|T047|AB|122.5|ICD9CM|Echinococ multiloc liver|Echinococ multiloc liver
C0153293|T047|PT|122.5|ICD9CM|Echinococcus multilocularis infection of liver|Echinococcus multilocularis infection of liver
C0277056|T047|AB|122.6|ICD9CM|Echinococc multiloc NEC|Echinococc multiloc NEC
C0277056|T047|PT|122.6|ICD9CM|Echinococcus multilocularis infection, other|Echinococcus multilocularis infection, other
C0152069|T047|AB|122.7|ICD9CM|Echinococc multiloc NOS|Echinococc multiloc NOS
C0152069|T047|PT|122.7|ICD9CM|Echinococcus multilocularis infection, unspecified|Echinococcus multilocularis infection, unspecified
C0013504|T047|AB|122.8|ICD9CM|Echinococcosis NOS liver|Echinococcosis NOS liver
C0013504|T047|PT|122.8|ICD9CM|Echinococcosis, unspecified, of liver|Echinococcosis, unspecified, of liver
C0348276|T047|AB|122.9|ICD9CM|Echinococcosis NEC/NOS|Echinococcosis NEC/NOS
C0348276|T047|PT|122.9|ICD9CM|Echinococcosis, other and unspecified|Echinococcosis, other and unspecified
C0153296|T047|HT|123|ICD9CM|Other cestode infection|Other cestode infection
C0473878|T047|PT|123.0|ICD9CM|Taenia solium infection, intestinal form|Taenia solium infection, intestinal form
C0473878|T047|AB|123.0|ICD9CM|Taenia solium intestine|Taenia solium intestine
C0010678|T047|AB|123.1|ICD9CM|Cysticercosis|Cysticercosis
C0010678|T047|PT|123.1|ICD9CM|Cysticercosis|Cysticercosis
C0152073|T047|AB|123.2|ICD9CM|Taenia saginata infect|Taenia saginata infect
C0152073|T047|PT|123.2|ICD9CM|Taenia saginata infection|Taenia saginata infection
C0039254|T047|AB|123.3|ICD9CM|Taeniasis NOS|Taeniasis NOS
C0039254|T047|PT|123.3|ICD9CM|Taeniasis, unspecified|Taeniasis, unspecified
C0012561|T047|AB|123.4|ICD9CM|Diphyllobothrias intest|Diphyllobothrias intest
C0012561|T047|PT|123.4|ICD9CM|Diphyllobothriasis, intestinal|Diphyllobothriasis, intestinal
C0037753|T047|AB|123.5|ICD9CM|Sparganosis|Sparganosis
C0037753|T047|PT|123.5|ICD9CM|Sparganosis [larval diphyllobothriasis]|Sparganosis [larval diphyllobothriasis]
C0020413|T047|AB|123.6|ICD9CM|Hymenolepiasis|Hymenolepiasis
C0020413|T047|PT|123.6|ICD9CM|Hymenolepiasis|Hymenolepiasis
C0029754|T047|AB|123.8|ICD9CM|Cestode infection NEC|Cestode infection NEC
C0029754|T047|PT|123.8|ICD9CM|Other specified cestode infection|Other specified cestode infection
C0007894|T047|AB|123.9|ICD9CM|Cestode infection NOS|Cestode infection NOS
C0007894|T047|PT|123.9|ICD9CM|Cestode infection, unspecified|Cestode infection, unspecified
C0040896|T047|AB|124|ICD9CM|Trichinosis|Trichinosis
C0040896|T047|PT|124|ICD9CM|Trichinosis|Trichinosis
C0153298|T047|HT|125|ICD9CM|Filarial infection and dracontiasis|Filarial infection and dracontiasis
C0392663|T047|AB|125.0|ICD9CM|Bancroftian filariasis|Bancroftian filariasis
C0392663|T047|PT|125.0|ICD9CM|Bancroftian filariasis|Bancroftian filariasis
C0152070|T047|AB|125.1|ICD9CM|Malayan filariasis|Malayan filariasis
C0152070|T047|PT|125.1|ICD9CM|Malayan filariasis|Malayan filariasis
C0023968|T047|AB|125.2|ICD9CM|Loiasis|Loiasis
C0023968|T047|PT|125.2|ICD9CM|Loiasis|Loiasis
C0029001|T047|AB|125.3|ICD9CM|Onchocerciasis|Onchocerciasis
C0029001|T047|PT|125.3|ICD9CM|Onchocerciasis|Onchocerciasis
C0012517|T047|AB|125.4|ICD9CM|Dipetalonemiasis|Dipetalonemiasis
C0012517|T047|PT|125.4|ICD9CM|Dipetalonemiasis|Dipetalonemiasis
C0016089|T047|AB|125.5|ICD9CM|Mansonella ozzardi infec|Mansonella ozzardi infec
C0016089|T047|PT|125.5|ICD9CM|Mansonella ozzardi infection|Mansonella ozzardi infection
C0029796|T047|AB|125.6|ICD9CM|Filariasis NEC|Filariasis NEC
C0029796|T047|PT|125.6|ICD9CM|Other specified filariasis|Other specified filariasis
C0013100|T047|AB|125.7|ICD9CM|Dracontiasis|Dracontiasis
C0013100|T047|PT|125.7|ICD9CM|Dracontiasis|Dracontiasis
C0016085|T047|AB|125.9|ICD9CM|Filariasis NOS|Filariasis NOS
C0016085|T047|PT|125.9|ICD9CM|Unspecified filariasis|Unspecified filariasis
C0411279|T047|HT|126|ICD9CM|Ancylostomiasis and necatoriasis|Ancylostomiasis and necatoriasis
C1384687|T047|AB|126.0|ICD9CM|Ancylostoma duodenale|Ancylostoma duodenale
C1384687|T047|PT|126.0|ICD9CM|Ancylostomiasis due to ancylostoma duodenale|Ancylostomiasis due to ancylostoma duodenale
C0027529|T047|AB|126.1|ICD9CM|Necator Americanus|Necator Americanus
C0027529|T047|PT|126.1|ICD9CM|Necatoriasis due to necator americanus|Necatoriasis due to necator americanus
C0153299|T047|AB|126.2|ICD9CM|Ancylostoma braziliense|Ancylostoma braziliense
C0153299|T047|PT|126.2|ICD9CM|Ancylostomiasis due to ancylostoma braziliense|Ancylostomiasis due to ancylostoma braziliense
C0277120|T047|AB|126.3|ICD9CM|Ancylostoma ceylanicum|Ancylostoma ceylanicum
C0277120|T047|PT|126.3|ICD9CM|Ancylostomiasis due to ancylostoma ceylanicum|Ancylostomiasis due to ancylostoma ceylanicum
C0546827|T047|AB|126.8|ICD9CM|Ancylostoma NEC|Ancylostoma NEC
C0546827|T047|PT|126.8|ICD9CM|Other specified ancylostoma|Other specified ancylostoma
C0411279|T047|PT|126.9|ICD9CM|Ancylostomiasis and necatoriasis, unspecified|Ancylostomiasis and necatoriasis, unspecified
C0411279|T047|AB|126.9|ICD9CM|Ancylostomiasis NOS|Ancylostomiasis NOS
C0153302|T047|HT|127|ICD9CM|Other intestinal helminthiases|Other intestinal helminthiases
C0003950|T047|AB|127.0|ICD9CM|Ascariasis|Ascariasis
C0003950|T047|PT|127.0|ICD9CM|Ascariasis|Ascariasis
C0162576|T047|AB|127.1|ICD9CM|Anisakiasis|Anisakiasis
C0162576|T047|PT|127.1|ICD9CM|Anisakiasis|Anisakiasis
C0038463|T047|AB|127.2|ICD9CM|Strongyloidiasis|Strongyloidiasis
C0038463|T047|PT|127.2|ICD9CM|Strongyloidiasis|Strongyloidiasis
C0040954|T047|AB|127.3|ICD9CM|Trichuriasis|Trichuriasis
C0040954|T047|PT|127.3|ICD9CM|Trichuriasis|Trichuriasis
C0086227|T047|AB|127.4|ICD9CM|Enterobiasis|Enterobiasis
C0086227|T047|PT|127.4|ICD9CM|Enterobiasis|Enterobiasis
C0006897|T047|AB|127.5|ICD9CM|Capillariasis|Capillariasis
C0006897|T047|PT|127.5|ICD9CM|Capillariasis|Capillariasis
C0040948|T047|AB|127.6|ICD9CM|Trichostrongyliasis|Trichostrongyliasis
C0040948|T047|PT|127.6|ICD9CM|Trichostrongyliasis|Trichostrongyliasis
C0029808|T047|AB|127.7|ICD9CM|Intest helminthiasis NEC|Intest helminthiasis NEC
C0029808|T047|PT|127.7|ICD9CM|Other specified intestinal helminthiasis|Other specified intestinal helminthiasis
C0153303|T047|PT|127.8|ICD9CM|Mixed intestinal helminthiasis|Mixed intestinal helminthiasis
C0153303|T047|AB|127.8|ICD9CM|Mixed intestine helminth|Mixed intestine helminth
C0348287|T047|AB|127.9|ICD9CM|Intest helminthiasis NOS|Intest helminthiasis NOS
C0348287|T047|PT|127.9|ICD9CM|Intestinal helminthiasis, unspecified|Intestinal helminthiasis, unspecified
C0494126|T047|HT|128|ICD9CM|Other and unspecified helminthiases|Other and unspecified helminthiases
C0040553|T047|AB|128.0|ICD9CM|Toxocariasis|Toxocariasis
C0040553|T047|PT|128.0|ICD9CM|Toxocariasis|Toxocariasis
C0018013|T047|AB|128.1|ICD9CM|Gnathostomiasis|Gnathostomiasis
C0018013|T047|PT|128.1|ICD9CM|Gnathostomiasis|Gnathostomiasis
C0029803|T047|AB|128.8|ICD9CM|Helminthiasis NEC|Helminthiasis NEC
C0029803|T047|PT|128.8|ICD9CM|Other specified helminthiasis|Other specified helminthiasis
C0018889|T047|PT|128.9|ICD9CM|Helminth infection, unspecified|Helminth infection, unspecified
C0018889|T047|AB|128.9|ICD9CM|Helminthiasis NOS|Helminthiasis NOS
C0021832|T047|AB|129|ICD9CM|Intestin parasitism NOS|Intestin parasitism NOS
C0021832|T047|PT|129|ICD9CM|Intestinal parasitism, unspecified|Intestinal parasitism, unspecified
C0040558|T047|HT|130|ICD9CM|Toxoplasmosis|Toxoplasmosis
C0153325|T047|HT|130-136.99|ICD9CM|OTHER INFECTIOUS AND PARASITIC DISEASES|OTHER INFECTIOUS AND PARASITIC DISEASES
C0085315|T047|PT|130.0|ICD9CM|Meningoencephalitis due to toxoplasmosis|Meningoencephalitis due to toxoplasmosis
C0085315|T047|AB|130.0|ICD9CM|Toxoplasm meningoenceph|Toxoplasm meningoenceph
C0153307|T047|PT|130.1|ICD9CM|Conjunctivitis due to toxoplasmosis|Conjunctivitis due to toxoplasmosis
C0153307|T047|AB|130.1|ICD9CM|Toxoplasm conjunctivitis|Toxoplasm conjunctivitis
C0153308|T047|PT|130.2|ICD9CM|Chorioretinitis due to toxoplasmosis|Chorioretinitis due to toxoplasmosis
C0153308|T047|AB|130.2|ICD9CM|Toxoplasm chorioretinit|Toxoplasm chorioretinit
C0276804|T047|PT|130.3|ICD9CM|Myocarditis due to toxoplasmosis|Myocarditis due to toxoplasmosis
C0276804|T047|AB|130.3|ICD9CM|Toxoplasma myocarditis|Toxoplasma myocarditis
C0339950|T047|PT|130.4|ICD9CM|Pneumonitis due to toxoplasmosis|Pneumonitis due to toxoplasmosis
C0339950|T047|AB|130.4|ICD9CM|Toxoplasma pneumonitis|Toxoplasma pneumonitis
C0400895|T047|PT|130.5|ICD9CM|Hepatitis due to toxoplasmosis|Hepatitis due to toxoplasmosis
C0400895|T047|AB|130.5|ICD9CM|Toxoplasma hepatitis|Toxoplasma hepatitis
C0153312|T047|PT|130.7|ICD9CM|Toxoplasmosis of other specified sites|Toxoplasmosis of other specified sites
C0153312|T047|AB|130.7|ICD9CM|Toxoplasmosis site NEC|Toxoplasmosis site NEC
C0343816|T047|AB|130.8|ICD9CM|Multisystem toxoplasmos|Multisystem toxoplasmos
C0343816|T047|PT|130.8|ICD9CM|Multisystemic disseminated toxoplasmosis|Multisystemic disseminated toxoplasmosis
C0040558|T047|AB|130.9|ICD9CM|Toxoplasmosis NOS|Toxoplasmosis NOS
C0040558|T047|PT|130.9|ICD9CM|Toxoplasmosis, unspecified|Toxoplasmosis, unspecified
C0040921|T047|HT|131|ICD9CM|Trichomoniasis|Trichomoniasis
C0040928|T047|HT|131.0|ICD9CM|Urogenital trichomoniasis|Urogenital trichomoniasis
C0040928|T047|AB|131.00|ICD9CM|Urogenital trichomon NOS|Urogenital trichomon NOS
C0040928|T047|PT|131.00|ICD9CM|Urogenital trichomoniasis, unspecified|Urogenital trichomoniasis, unspecified
C2945558|T047|AB|131.01|ICD9CM|Trichomonal vaginitis|Trichomonal vaginitis
C2945558|T047|PT|131.01|ICD9CM|Trichomonal vulvovaginitis|Trichomonal vulvovaginitis
C0153314|T047|AB|131.02|ICD9CM|Trichomonal urethritis|Trichomonal urethritis
C0153314|T047|PT|131.02|ICD9CM|Trichomonal urethritis|Trichomonal urethritis
C0153315|T047|AB|131.03|ICD9CM|Trichomonal prostatitis|Trichomonal prostatitis
C0153315|T047|PT|131.03|ICD9CM|Trichomonal prostatitis|Trichomonal prostatitis
C0153316|T047|PT|131.09|ICD9CM|Other urogenital trichomoniasis|Other urogenital trichomoniasis
C0153316|T047|AB|131.09|ICD9CM|Urogenital trichomon NEC|Urogenital trichomon NEC
C0040926|T047|AB|131.8|ICD9CM|Trichomoniasis NEC|Trichomoniasis NEC
C0040926|T047|PT|131.8|ICD9CM|Trichomoniasis of other specified sites|Trichomoniasis of other specified sites
C0040921|T047|AB|131.9|ICD9CM|Trichomoniasis NOS|Trichomoniasis NOS
C0040921|T047|PT|131.9|ICD9CM|Trichomoniasis, unspecified|Trichomoniasis, unspecified
C0153317|T047|HT|132|ICD9CM|Pediculosis and phthirus infestation|Pediculosis and phthirus infestation
C0030757|T047|AB|132.0|ICD9CM|Pediculus capitis|Pediculus capitis
C0030757|T047|PT|132.0|ICD9CM|Pediculus capitis [head louse]|Pediculus capitis [head louse]
C0030758|T047|AB|132.1|ICD9CM|Pediculus corporis|Pediculus corporis
C0030758|T047|PT|132.1|ICD9CM|Pediculus corporis [body louse]|Pediculus corporis [body louse]
C0030759|T047|AB|132.2|ICD9CM|Phthirus pubis|Phthirus pubis
C0030759|T047|PT|132.2|ICD9CM|Phthirus pubis [pubic louse]|Phthirus pubis [pubic louse]
C0277351|T047|AB|132.3|ICD9CM|Mixed pedicul & phthirus|Mixed pedicul & phthirus
C0277351|T047|PT|132.3|ICD9CM|Mixed pediculosis infestation|Mixed pediculosis infestation
C0030756|T047|AB|132.9|ICD9CM|Pediculosis NOS|Pediculosis NOS
C0030756|T047|PT|132.9|ICD9CM|Pediculosis, unspecified|Pediculosis, unspecified
C0026229|T047|HT|133|ICD9CM|Acariasis|Acariasis
C0036262|T047|AB|133.0|ICD9CM|Scabies|Scabies
C0036262|T047|PT|133.0|ICD9CM|Scabies|Scabies
C0029482|T047|AB|133.8|ICD9CM|Acariasis NEC|Acariasis NEC
C0029482|T047|PT|133.8|ICD9CM|Other acariasis|Other acariasis
C0026229|T047|AB|133.9|ICD9CM|Acariasis NOS|Acariasis NOS
C0026229|T047|PT|133.9|ICD9CM|Acariasis, unspecified|Acariasis, unspecified
C0153322|T047|HT|134|ICD9CM|Other infestation|Other infestation
C0027030|T047|AB|134.0|ICD9CM|Myiasis|Myiasis
C0027030|T047|PT|134.0|ICD9CM|Myiasis|Myiasis
C0153323|T047|AB|134.1|ICD9CM|Arthropod infest NEC|Arthropod infest NEC
C0153323|T047|PT|134.1|ICD9CM|Other arthropod infestation|Other arthropod infestation
C0019575|T047|AB|134.2|ICD9CM|Hirudiniasis|Hirudiniasis
C0019575|T047|PT|134.2|ICD9CM|Hirudiniasis|Hirudiniasis
C0153324|T047|AB|134.8|ICD9CM|Infestation NEC|Infestation NEC
C0153324|T047|PT|134.8|ICD9CM|Other specified infestations|Other specified infestations
C0851341|T047|AB|134.9|ICD9CM|Infestation NOS|Infestation NOS
C0851341|T047|PT|134.9|ICD9CM|Infestation, unspecified|Infestation, unspecified
C0036202|T047|AB|135|ICD9CM|Sarcoidosis|Sarcoidosis
C0036202|T047|PT|135|ICD9CM|Sarcoidosis|Sarcoidosis
C0153325|T047|HT|136|ICD9CM|Other and unspecified infectious and parasitic diseases|Other and unspecified infectious and parasitic diseases
C0001860|T047|AB|136.0|ICD9CM|Ainhum|Ainhum
C0001860|T047|PT|136.0|ICD9CM|Ainhum|Ainhum
C0004943|T047|AB|136.1|ICD9CM|Behcet's syndrome|Behcet's syndrome
C0004943|T047|PT|136.1|ICD9CM|Behcet's syndrome|Behcet's syndrome
C0153326|T047|HT|136.2|ICD9CM|Specific infections by free-living amebae|Specific infections by free-living amebae
C2349230|T047|AB|136.21|ICD9CM|Infectn d/t acanthamoeba|Infectn d/t acanthamoeba
C2349230|T047|PT|136.21|ICD9CM|Specific infection due to acanthamoeba|Specific infection due to acanthamoeba
C2349231|T047|AB|136.29|ICD9CM|Infc free-liv amebae NEC|Infc free-liv amebae NEC
C2349231|T047|PT|136.29|ICD9CM|Other specific infections by free-living amebae|Other specific infections by free-living amebae
C1535939|T047|AB|136.3|ICD9CM|Pneumocystosis|Pneumocystosis
C1535939|T047|PT|136.3|ICD9CM|Pneumocystosis|Pneumocystosis
C0153327|T047|AB|136.4|ICD9CM|Psorospermiasis|Psorospermiasis
C0153327|T047|PT|136.4|ICD9CM|Psorospermiasis|Psorospermiasis
C0036231|T047|AB|136.5|ICD9CM|Sarcosporidiosis|Sarcosporidiosis
C0036231|T047|PT|136.5|ICD9CM|Sarcosporidiosis|Sarcosporidiosis
C0153328|T047|AB|136.8|ICD9CM|Infect/parasite dis NEC|Infect/parasite dis NEC
C0153328|T047|PT|136.8|ICD9CM|Other specified infectious and parasitic diseases|Other specified infectious and parasitic diseases
C0041849|T047|AB|136.9|ICD9CM|Infect/parasite dis NOS|Infect/parasite dis NOS
C0041849|T047|PT|136.9|ICD9CM|Unspecified infectious and parasitic diseases|Unspecified infectious and parasitic diseases
C0153329|T046|HT|137|ICD9CM|Late effects of tuberculosis|Late effects of tuberculosis
C0348296|T047|HT|137-139.99|ICD9CM|LATE EFFECTS OF INFECTIOUS AND PARASITIC DISEASES|LATE EFFECTS OF INFECTIOUS AND PARASITIC DISEASES
C0343413|T047|AB|137.0|ICD9CM|Late effect tb, resp/NOS|Late effect tb, resp/NOS
C0343413|T047|PT|137.0|ICD9CM|Late effects of respiratory or unspecified tuberculosis|Late effects of respiratory or unspecified tuberculosis
C0153331|T046|AB|137.1|ICD9CM|Late effect cns TB|Late effect cns TB
C0153331|T046|PT|137.1|ICD9CM|Late effects of central nervous system tuberculosis|Late effects of central nervous system tuberculosis
C0343422|T046|AB|137.2|ICD9CM|Late effect gu TB|Late effect gu TB
C0343422|T046|PT|137.2|ICD9CM|Late effects of genitourinary tuberculosis|Late effects of genitourinary tuberculosis
C0153333|T046|AB|137.3|ICD9CM|Late eff bone & joint TB|Late eff bone & joint TB
C0153333|T046|PT|137.3|ICD9CM|Late effects of tuberculosis of bones and joints|Late effects of tuberculosis of bones and joints
C0153334|T046|AB|137.4|ICD9CM|Late effect TB NEC|Late effect TB NEC
C0153334|T046|PT|137.4|ICD9CM|Late effects of tuberculosis of other specified organs|Late effects of tuberculosis of other specified organs
C0362050|T046|AB|138|ICD9CM|Late effect acute polio|Late effect acute polio
C0362050|T046|PT|138|ICD9CM|Late effects of acute poliomyelitis|Late effects of acute poliomyelitis
C0153336|T046|HT|139|ICD9CM|Late effects of other infectious and parasitic diseases|Late effects of other infectious and parasitic diseases
C0153337|T046|AB|139.0|ICD9CM|Late eff viral encephal|Late eff viral encephal
C0153337|T046|PT|139.0|ICD9CM|Late effects of viral encephalitis|Late effects of viral encephalitis
C0153338|T047|AB|139.1|ICD9CM|Late effect of trachoma|Late effect of trachoma
C0153338|T047|PT|139.1|ICD9CM|Late effects of trachoma|Late effects of trachoma
C0153336|T046|AB|139.8|ICD9CM|Late eff infect dis NEC|Late eff infect dis NEC
C0153336|T046|PT|139.8|ICD9CM|Late effects of other and unspecified infectious and parasitic diseases|Late effects of other and unspecified infectious and parasitic diseases
C0153340|T191|HT|140|ICD9CM|Malignant neoplasm of lip|Malignant neoplasm of lip
C0178247|T191|HT|140-149.99|ICD9CM|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY, AND PHARYNX|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY, AND PHARYNX
C0027651|T191|HT|140-239.99|ICD9CM|NEOPLASMS|NEOPLASMS
C0474962|T191|AB|140.0|ICD9CM|Mal neo upper vermilion|Mal neo upper vermilion
C0474962|T191|PT|140.0|ICD9CM|Malignant neoplasm of upper lip, vermilion border|Malignant neoplasm of upper lip, vermilion border
C0432520|T191|AB|140.1|ICD9CM|Mal neo lower vermilion|Mal neo lower vermilion
C0432520|T191|PT|140.1|ICD9CM|Malignant neoplasm of lower lip, vermilion border|Malignant neoplasm of lower lip, vermilion border
C0432579|T191|AB|140.3|ICD9CM|Mal neo upper lip, inner|Mal neo upper lip, inner
C0432579|T191|PT|140.3|ICD9CM|Malignant neoplasm of upper lip, inner aspect|Malignant neoplasm of upper lip, inner aspect
C0733940|T191|AB|140.4|ICD9CM|Mal neo lower lip, inner|Mal neo lower lip, inner
C0733940|T191|PT|140.4|ICD9CM|Malignant neoplasm of lower lip, inner aspect|Malignant neoplasm of lower lip, inner aspect
C0474971|T191|AB|140.5|ICD9CM|Mal neo lip, inner NOS|Mal neo lip, inner NOS
C0474971|T191|PT|140.5|ICD9CM|Malignant neoplasm of lip, unspecified, inner aspect|Malignant neoplasm of lip, unspecified, inner aspect
C0153346|T191|AB|140.6|ICD9CM|Mal neo lip, commissure|Mal neo lip, commissure
C0153346|T191|PT|140.6|ICD9CM|Malignant neoplasm of commissure of lip|Malignant neoplasm of commissure of lip
C0153347|T191|AB|140.8|ICD9CM|Mal neo lip NEC|Mal neo lip NEC
C0153347|T191|PT|140.8|ICD9CM|Malignant neoplasm of other sites of lip|Malignant neoplasm of other sites of lip
C0546836|T191|AB|140.9|ICD9CM|Mal neo lip/vermil NOS|Mal neo lip/vermil NOS
C0546836|T191|PT|140.9|ICD9CM|Malignant neoplasm of lip, unspecified, vermilion border|Malignant neoplasm of lip, unspecified, vermilion border
C0153349|T191|HT|141|ICD9CM|Malignant neoplasm of tongue|Malignant neoplasm of tongue
C0153350|T191|AB|141.0|ICD9CM|Mal neo tongue base|Mal neo tongue base
C0153350|T191|PT|141.0|ICD9CM|Malignant neoplasm of base of tongue|Malignant neoplasm of base of tongue
C0153351|T191|AB|141.1|ICD9CM|Mal neo dorsal tongue|Mal neo dorsal tongue
C0153351|T191|PT|141.1|ICD9CM|Malignant neoplasm of dorsal surface of tongue|Malignant neoplasm of dorsal surface of tongue
C0496755|T191|AB|141.2|ICD9CM|Mal neo tip/lat tongue|Mal neo tip/lat tongue
C0496755|T191|PT|141.2|ICD9CM|Malignant neoplasm of tip and lateral border of tongue|Malignant neoplasm of tip and lateral border of tongue
C0684333|T191|AB|141.3|ICD9CM|Mal neo ventral tongue|Mal neo ventral tongue
C0684333|T191|PT|141.3|ICD9CM|Malignant neoplasm of ventral surface of tongue|Malignant neoplasm of ventral surface of tongue
C0153354|T191|AB|141.4|ICD9CM|Mal neo ant 2/3 tongue|Mal neo ant 2/3 tongue
C0153354|T191|PT|141.4|ICD9CM|Malignant neoplasm of anterior two-thirds of tongue, part unspecified|Malignant neoplasm of anterior two-thirds of tongue, part unspecified
C0474963|T191|AB|141.5|ICD9CM|Mal neo tongue junction|Mal neo tongue junction
C0474963|T191|PT|141.5|ICD9CM|Malignant neoplasm of junctional zone of tongue|Malignant neoplasm of junctional zone of tongue
C0153356|T191|AB|141.6|ICD9CM|Mal neo lingual tonsil|Mal neo lingual tonsil
C0153356|T191|PT|141.6|ICD9CM|Malignant neoplasm of lingual tonsil|Malignant neoplasm of lingual tonsil
C0153357|T191|AB|141.8|ICD9CM|Malig neo tongue NEC|Malig neo tongue NEC
C0153357|T191|PT|141.8|ICD9CM|Malignant neoplasm of other sites of tongue|Malignant neoplasm of other sites of tongue
C0153349|T191|AB|141.9|ICD9CM|Malig neo tongue NOS|Malig neo tongue NOS
C0153349|T191|PT|141.9|ICD9CM|Malignant neoplasm of tongue, unspecified|Malignant neoplasm of tongue, unspecified
C0496763|T191|HT|142|ICD9CM|Malignant neoplasm of major salivary glands|Malignant neoplasm of major salivary glands
C0747273|T191|AB|142.0|ICD9CM|Malig neo parotid|Malig neo parotid
C0747273|T191|PT|142.0|ICD9CM|Malignant neoplasm of parotid gland|Malignant neoplasm of parotid gland
C0153360|T191|AB|142.1|ICD9CM|Malig neo submandibular|Malig neo submandibular
C0153360|T191|PT|142.1|ICD9CM|Malignant neoplasm of submandibular gland|Malignant neoplasm of submandibular gland
C0153361|T191|AB|142.2|ICD9CM|Malig neo sublingual|Malig neo sublingual
C0153361|T191|PT|142.2|ICD9CM|Malignant neoplasm of sublingual gland|Malignant neoplasm of sublingual gland
C0153362|T191|AB|142.8|ICD9CM|Mal neo maj salivary NEC|Mal neo maj salivary NEC
C0153362|T191|PT|142.8|ICD9CM|Malignant neoplasm of other major salivary glands|Malignant neoplasm of other major salivary glands
C0220636|T191|AB|142.9|ICD9CM|Mal neo salivary NOS|Mal neo salivary NOS
C0220636|T191|PT|142.9|ICD9CM|Malignant neoplasm of salivary gland, unspecified|Malignant neoplasm of salivary gland, unspecified
C0153364|T191|HT|143|ICD9CM|Malignant neoplasm of gum|Malignant neoplasm of gum
C0153365|T191|AB|143.0|ICD9CM|Malig neo upper gum|Malig neo upper gum
C0153365|T191|PT|143.0|ICD9CM|Malignant neoplasm of upper gum|Malignant neoplasm of upper gum
C0432581|T191|AB|143.1|ICD9CM|Malig neo lower gum|Malig neo lower gum
C0432581|T191|PT|143.1|ICD9CM|Malignant neoplasm of lower gum|Malignant neoplasm of lower gum
C0153367|T191|AB|143.8|ICD9CM|Malig neo gum NEC|Malig neo gum NEC
C0153367|T191|PT|143.8|ICD9CM|Malignant neoplasm of other sites of gum|Malignant neoplasm of other sites of gum
C0153364|T191|AB|143.9|ICD9CM|Malig neo gum NOS|Malig neo gum NOS
C0153364|T191|PT|143.9|ICD9CM|Malignant neoplasm of gum, unspecified|Malignant neoplasm of gum, unspecified
C0153368|T191|HT|144|ICD9CM|Malignant neoplasm of floor of mouth|Malignant neoplasm of floor of mouth
C0153369|T191|AB|144.0|ICD9CM|Mal neo ant floor mouth|Mal neo ant floor mouth
C0153369|T191|PT|144.0|ICD9CM|Malignant neoplasm of anterior portion of floor of mouth|Malignant neoplasm of anterior portion of floor of mouth
C0496758|T191|AB|144.1|ICD9CM|Mal neo lat floor mouth|Mal neo lat floor mouth
C0496758|T191|PT|144.1|ICD9CM|Malignant neoplasm of lateral portion of floor of mouth|Malignant neoplasm of lateral portion of floor of mouth
C0153371|T191|AB|144.8|ICD9CM|Mal neo mouth floor NEC|Mal neo mouth floor NEC
C0153371|T191|PT|144.8|ICD9CM|Malignant neoplasm of other sites of floor of mouth|Malignant neoplasm of other sites of floor of mouth
C0153368|T191|AB|144.9|ICD9CM|Mal neo mouth floor NOS|Mal neo mouth floor NOS
C0153368|T191|PT|144.9|ICD9CM|Malignant neoplasm of floor of mouth, part unspecified|Malignant neoplasm of floor of mouth, part unspecified
C0153372|T191|HT|145|ICD9CM|Malignant neoplasm of other and unspecified parts of mouth|Malignant neoplasm of other and unspecified parts of mouth
C0153373|T191|AB|145.0|ICD9CM|Mal neo cheek mucosa|Mal neo cheek mucosa
C0153373|T191|PT|145.0|ICD9CM|Malignant neoplasm of cheek mucosa|Malignant neoplasm of cheek mucosa
C0153374|T191|AB|145.1|ICD9CM|Mal neo mouth vestibule|Mal neo mouth vestibule
C0153374|T191|PT|145.1|ICD9CM|Malignant neoplasm of vestibule of mouth|Malignant neoplasm of vestibule of mouth
C0153375|T191|AB|145.2|ICD9CM|Malig neo hard palate|Malig neo hard palate
C0153375|T191|PT|145.2|ICD9CM|Malignant neoplasm of hard palate|Malignant neoplasm of hard palate
C0153376|T191|AB|145.3|ICD9CM|Malig neo soft palate|Malig neo soft palate
C0153376|T191|PT|145.3|ICD9CM|Malignant neoplasm of soft palate|Malignant neoplasm of soft palate
C0153377|T191|PT|145.4|ICD9CM|Malignant neoplasm of uvula|Malignant neoplasm of uvula
C0153377|T191|AB|145.4|ICD9CM|Malignant neoplasm uvula|Malignant neoplasm uvula
C0153378|T191|AB|145.5|ICD9CM|Malignant neo palate NOS|Malignant neo palate NOS
C0153378|T191|PT|145.5|ICD9CM|Malignant neoplasm of palate, unspecified|Malignant neoplasm of palate, unspecified
C0153379|T191|AB|145.6|ICD9CM|Malig neo retromolar|Malig neo retromolar
C0153379|T191|PT|145.6|ICD9CM|Malignant neoplasm of retromolar area|Malignant neoplasm of retromolar area
C0153380|T191|AB|145.8|ICD9CM|Malig neoplasm mouth NEC|Malig neoplasm mouth NEC
C0153380|T191|PT|145.8|ICD9CM|Malignant neoplasm of other specified parts of mouth|Malignant neoplasm of other specified parts of mouth
C0153381|T191|AB|145.9|ICD9CM|Malig neoplasm mouth NOS|Malig neoplasm mouth NOS
C0153381|T191|PT|145.9|ICD9CM|Malignant neoplasm of mouth, unspecified|Malignant neoplasm of mouth, unspecified
C0153382|T191|HT|146|ICD9CM|Malignant neoplasm of oropharynx|Malignant neoplasm of oropharynx
C0751560|T191|AB|146.0|ICD9CM|Malignant neopl tonsil|Malignant neopl tonsil
C0751560|T191|PT|146.0|ICD9CM|Malignant neoplasm of tonsil|Malignant neoplasm of tonsil
C0153384|T191|AB|146.1|ICD9CM|Mal neo tonsillar fossa|Mal neo tonsillar fossa
C0153384|T191|PT|146.1|ICD9CM|Malignant neoplasm of tonsillar fossa|Malignant neoplasm of tonsillar fossa
C0153385|T191|AB|146.2|ICD9CM|Mal neo tonsil pillars|Mal neo tonsil pillars
C0153385|T191|PT|146.2|ICD9CM|Malignant neoplasm of tonsillar pillars (anterior) (posterior)|Malignant neoplasm of tonsillar pillars (anterior) (posterior)
C0153386|T191|AB|146.3|ICD9CM|Malign neopl vallecula|Malign neopl vallecula
C0153386|T191|PT|146.3|ICD9CM|Malignant neoplasm of vallecula epiglottica|Malignant neoplasm of vallecula epiglottica
C0496765|T191|AB|146.4|ICD9CM|Mal neo ant epiglottis|Mal neo ant epiglottis
C0496765|T191|PT|146.4|ICD9CM|Malignant neoplasm of anterior aspect of epiglottis|Malignant neoplasm of anterior aspect of epiglottis
C0153388|T191|AB|146.5|ICD9CM|Mal neo epiglottis junct|Mal neo epiglottis junct
C0153388|T191|PT|146.5|ICD9CM|Malignant neoplasm of junctional region of oropharynx|Malignant neoplasm of junctional region of oropharynx
C0153389|T191|AB|146.6|ICD9CM|Mal neo lat oropharynx|Mal neo lat oropharynx
C0153389|T191|PT|146.6|ICD9CM|Malignant neoplasm of lateral wall of oropharynx|Malignant neoplasm of lateral wall of oropharynx
C0153390|T191|AB|146.7|ICD9CM|Mal neo post oropharynx|Mal neo post oropharynx
C0153390|T191|PT|146.7|ICD9CM|Malignant neoplasm of posterior wall of oropharynx|Malignant neoplasm of posterior wall of oropharynx
C0153391|T191|AB|146.8|ICD9CM|Mal neo oropharynx NEC|Mal neo oropharynx NEC
C0153391|T191|PT|146.8|ICD9CM|Malignant neoplasm of other specified sites of oropharynx|Malignant neoplasm of other specified sites of oropharynx
C0153382|T191|AB|146.9|ICD9CM|Malig neo oropharynx NOS|Malig neo oropharynx NOS
C0153382|T191|PT|146.9|ICD9CM|Malignant neoplasm of oropharynx, unspecified site|Malignant neoplasm of oropharynx, unspecified site
C0153392|T191|HT|147|ICD9CM|Malignant neoplasm of nasopharynx|Malignant neoplasm of nasopharynx
C0153393|T191|AB|147.0|ICD9CM|Mal neo super nasopharyn|Mal neo super nasopharyn
C0153393|T191|PT|147.0|ICD9CM|Malignant neoplasm of superior wall of nasopharynx|Malignant neoplasm of superior wall of nasopharynx
C0153394|T191|AB|147.1|ICD9CM|Mal neo post nasopharynx|Mal neo post nasopharynx
C0153394|T191|PT|147.1|ICD9CM|Malignant neoplasm of posterior wall of nasopharynx|Malignant neoplasm of posterior wall of nasopharynx
C0153395|T191|AB|147.2|ICD9CM|Mal neo lat nasopharynx|Mal neo lat nasopharynx
C0153395|T191|PT|147.2|ICD9CM|Malignant neoplasm of lateral wall of nasopharynx|Malignant neoplasm of lateral wall of nasopharynx
C0153396|T191|AB|147.3|ICD9CM|Mal neo ant nasopharynx|Mal neo ant nasopharynx
C0153396|T191|PT|147.3|ICD9CM|Malignant neoplasm of anterior wall of nasopharynx|Malignant neoplasm of anterior wall of nasopharynx
C0153397|T191|AB|147.8|ICD9CM|Mal neo nasopharynx NEC|Mal neo nasopharynx NEC
C0153397|T191|PT|147.8|ICD9CM|Malignant neoplasm of other specified sites of nasopharynx|Malignant neoplasm of other specified sites of nasopharynx
C0153392|T191|AB|147.9|ICD9CM|Mal neo nasopharynx NOS|Mal neo nasopharynx NOS
C0153392|T191|PT|147.9|ICD9CM|Malignant neoplasm of nasopharynx, unspecified site|Malignant neoplasm of nasopharynx, unspecified site
C0153398|T191|HT|148|ICD9CM|Malignant neoplasm of hypopharynx|Malignant neoplasm of hypopharynx
C0496769|T191|AB|148.0|ICD9CM|Mal neo postcricoid|Mal neo postcricoid
C0496769|T191|PT|148.0|ICD9CM|Malignant neoplasm of postcricoid region of hypopharynx|Malignant neoplasm of postcricoid region of hypopharynx
C0153400|T191|AB|148.1|ICD9CM|Mal neo pyriform sinus|Mal neo pyriform sinus
C0153400|T191|PT|148.1|ICD9CM|Malignant neoplasm of pyriform sinus|Malignant neoplasm of pyriform sinus
C0153401|T191|AB|148.2|ICD9CM|Mal neo aryepiglott fold|Mal neo aryepiglott fold
C0153401|T191|PT|148.2|ICD9CM|Malignant neoplasm of aryepiglottic fold, hypopharyngeal aspect|Malignant neoplasm of aryepiglottic fold, hypopharyngeal aspect
C0496770|T191|AB|148.3|ICD9CM|Mal neo post hypopharynx|Mal neo post hypopharynx
C0496770|T191|PT|148.3|ICD9CM|Malignant neoplasm of posterior hypopharyngeal wall|Malignant neoplasm of posterior hypopharyngeal wall
C0153403|T191|AB|148.8|ICD9CM|Mal neo hypopharynx NEC|Mal neo hypopharynx NEC
C0153403|T191|PT|148.8|ICD9CM|Malignant neoplasm of other specified sites of hypopharynx|Malignant neoplasm of other specified sites of hypopharynx
C0153398|T191|AB|148.9|ICD9CM|Mal neo hypopharynx NOS|Mal neo hypopharynx NOS
C0153398|T191|PT|148.9|ICD9CM|Malignant neoplasm of hypopharynx, unspecified site|Malignant neoplasm of hypopharynx, unspecified site
C0153404|T191|HT|149|ICD9CM|Malignant neoplasm of other and ill-defined sites within the lip, oral cavity, and pharynx|Malignant neoplasm of other and ill-defined sites within the lip, oral cavity, and pharynx
C0153405|T191|AB|149.0|ICD9CM|Mal neo pharynx NOS|Mal neo pharynx NOS
C0153405|T191|PT|149.0|ICD9CM|Malignant neoplasm of pharynx, unspecified|Malignant neoplasm of pharynx, unspecified
C0153406|T191|AB|149.1|ICD9CM|Mal neo waldeyer's ring|Mal neo waldeyer's ring
C0153406|T191|PT|149.1|ICD9CM|Malignant neoplasm of waldeyer's ring|Malignant neoplasm of waldeyer's ring
C0153407|T191|AB|149.8|ICD9CM|Mal neo oral/pharynx NEC|Mal neo oral/pharynx NEC
C0153407|T191|PT|149.8|ICD9CM|Malignant neoplasm of other sites within the lip and oral cavity|Malignant neoplasm of other sites within the lip and oral cavity
C0153408|T191|AB|149.9|ICD9CM|Mal neo orophryn ill-def|Mal neo orophryn ill-def
C0153408|T191|PT|149.9|ICD9CM|Malignant neoplasm of ill-defined sites within the lip and oral cavity|Malignant neoplasm of ill-defined sites within the lip and oral cavity
C0546837|T191|HT|150|ICD9CM|Malignant neoplasm of esophagus|Malignant neoplasm of esophagus
C0555264|T191|HT|150-159.99|ICD9CM|MALIGNANT NEOPLASM OF DIGESTIVE ORGANS AND PERITONEUM|MALIGNANT NEOPLASM OF DIGESTIVE ORGANS AND PERITONEUM
C0496773|T191|AB|150.0|ICD9CM|Mal neo cervical esophag|Mal neo cervical esophag
C0496773|T191|PT|150.0|ICD9CM|Malignant neoplasm of cervical esophagus|Malignant neoplasm of cervical esophagus
C0153411|T191|AB|150.1|ICD9CM|Mal neo thoracic esophag|Mal neo thoracic esophag
C0153411|T191|PT|150.1|ICD9CM|Malignant neoplasm of thoracic esophagus|Malignant neoplasm of thoracic esophagus
C0496775|T191|AB|150.2|ICD9CM|Mal neo abdomin esophag|Mal neo abdomin esophag
C0496775|T191|PT|150.2|ICD9CM|Malignant neoplasm of abdominal esophagus|Malignant neoplasm of abdominal esophagus
C0153413|T191|AB|150.3|ICD9CM|Mal neo upper 3rd esoph|Mal neo upper 3rd esoph
C0153413|T191|PT|150.3|ICD9CM|Malignant neoplasm of upper third of esophagus|Malignant neoplasm of upper third of esophagus
C0153414|T191|AB|150.4|ICD9CM|Mal neo middle 3rd esoph|Mal neo middle 3rd esoph
C0153414|T191|PT|150.4|ICD9CM|Malignant neoplasm of middle third of esophagus|Malignant neoplasm of middle third of esophagus
C0153415|T191|AB|150.5|ICD9CM|Mal neo lower 3rd esoph|Mal neo lower 3rd esoph
C0153415|T191|PT|150.5|ICD9CM|Malignant neoplasm of lower third of esophagus|Malignant neoplasm of lower third of esophagus
C0153416|T191|AB|150.8|ICD9CM|Mal neo esophagus NEC|Mal neo esophagus NEC
C0153416|T191|PT|150.8|ICD9CM|Malignant neoplasm of other specified part of esophagus|Malignant neoplasm of other specified part of esophagus
C0546837|T191|AB|150.9|ICD9CM|Mal neo esophagus NOS|Mal neo esophagus NOS
C0546837|T191|PT|150.9|ICD9CM|Malignant neoplasm of esophagus, unspecified site|Malignant neoplasm of esophagus, unspecified site
C0024623|T191|HT|151|ICD9CM|Malignant neoplasm of stomach|Malignant neoplasm of stomach
C0153417|T191|AB|151.0|ICD9CM|Mal neo stomach cardia|Mal neo stomach cardia
C0153417|T191|PT|151.0|ICD9CM|Malignant neoplasm of cardia|Malignant neoplasm of cardia
C0153418|T191|AB|151.1|ICD9CM|Malignant neo pylorus|Malignant neo pylorus
C0153418|T191|PT|151.1|ICD9CM|Malignant neoplasm of pylorus|Malignant neoplasm of pylorus
C0153419|T191|AB|151.2|ICD9CM|Mal neo pyloric antrum|Mal neo pyloric antrum
C0153419|T191|PT|151.2|ICD9CM|Malignant neoplasm of pyloric antrum|Malignant neoplasm of pyloric antrum
C0153420|T191|AB|151.3|ICD9CM|Mal neo stomach fundus|Mal neo stomach fundus
C0153420|T191|PT|151.3|ICD9CM|Malignant neoplasm of fundus of stomach|Malignant neoplasm of fundus of stomach
C0153421|T191|AB|151.4|ICD9CM|Mal neo stomach body|Mal neo stomach body
C0153421|T191|PT|151.4|ICD9CM|Malignant neoplasm of body of stomach|Malignant neoplasm of body of stomach
C0153422|T191|AB|151.5|ICD9CM|Mal neo stom lesser curv|Mal neo stom lesser curv
C0153422|T191|PT|151.5|ICD9CM|Malignant neoplasm of lesser curvature of stomach, unspecified|Malignant neoplasm of lesser curvature of stomach, unspecified
C0153423|T191|AB|151.6|ICD9CM|Mal neo stom great curv|Mal neo stom great curv
C0153423|T191|PT|151.6|ICD9CM|Malignant neoplasm of greater curvature of stomach, unspecified|Malignant neoplasm of greater curvature of stomach, unspecified
C0153424|T191|AB|151.8|ICD9CM|Malig neopl stomach NEC|Malig neopl stomach NEC
C0153424|T191|PT|151.8|ICD9CM|Malignant neoplasm of other specified sites of stomach|Malignant neoplasm of other specified sites of stomach
C0024623|T191|AB|151.9|ICD9CM|Malig neopl stomach NOS|Malig neopl stomach NOS
C0024623|T191|PT|151.9|ICD9CM|Malignant neoplasm of stomach, unspecified site|Malignant neoplasm of stomach, unspecified site
C1112753|T191|HT|152|ICD9CM|Malignant neoplasm of small intestine, including duodenum|Malignant neoplasm of small intestine, including duodenum
C0153426|T191|AB|152.0|ICD9CM|Malignant neopl duodenum|Malignant neopl duodenum
C0153426|T191|PT|152.0|ICD9CM|Malignant neoplasm of duodenum|Malignant neoplasm of duodenum
C0153427|T191|AB|152.1|ICD9CM|Malignant neopl jejunum|Malignant neopl jejunum
C0153427|T191|PT|152.1|ICD9CM|Malignant neoplasm of jejunum|Malignant neoplasm of jejunum
C0153428|T191|AB|152.2|ICD9CM|Malignant neoplasm ileum|Malignant neoplasm ileum
C0153428|T191|PT|152.2|ICD9CM|Malignant neoplasm of ileum|Malignant neoplasm of ileum
C0153429|T191|AB|152.3|ICD9CM|Mal neo meckel's divert|Mal neo meckel's divert
C0153429|T191|PT|152.3|ICD9CM|Malignant neoplasm of Meckel's diverticulum|Malignant neoplasm of Meckel's diverticulum
C0153430|T191|AB|152.8|ICD9CM|Mal neo small bowel NEC|Mal neo small bowel NEC
C0153430|T191|PT|152.8|ICD9CM|Malignant neoplasm of other specified sites of small intestine|Malignant neoplasm of other specified sites of small intestine
C0153425|T191|AB|152.9|ICD9CM|Mal neo small bowel NOS|Mal neo small bowel NOS
C0153425|T191|PT|152.9|ICD9CM|Malignant neoplasm of small intestine, unspecified site|Malignant neoplasm of small intestine, unspecified site
C0007102|T191|HT|153|ICD9CM|Malignant neoplasm of colon|Malignant neoplasm of colon
C0153433|T191|AB|153.0|ICD9CM|Mal neo hepatic flexure|Mal neo hepatic flexure
C0153433|T191|PT|153.0|ICD9CM|Malignant neoplasm of hepatic flexure|Malignant neoplasm of hepatic flexure
C0153434|T191|AB|153.1|ICD9CM|Mal neo transverse colon|Mal neo transverse colon
C0153434|T191|PT|153.1|ICD9CM|Malignant neoplasm of transverse colon|Malignant neoplasm of transverse colon
C0153435|T191|AB|153.2|ICD9CM|Mal neo descend colon|Mal neo descend colon
C0153435|T191|PT|153.2|ICD9CM|Malignant neoplasm of descending colon|Malignant neoplasm of descending colon
C0153436|T191|AB|153.3|ICD9CM|Mal neo sigmoid colon|Mal neo sigmoid colon
C0153436|T191|PT|153.3|ICD9CM|Malignant neoplasm of sigmoid colon|Malignant neoplasm of sigmoid colon
C0153437|T191|AB|153.4|ICD9CM|Malignant neoplasm cecum|Malignant neoplasm cecum
C0153437|T191|PT|153.4|ICD9CM|Malignant neoplasm of cecum|Malignant neoplasm of cecum
C0496779|T191|AB|153.5|ICD9CM|Malignant neo appendix|Malignant neo appendix
C0496779|T191|PT|153.5|ICD9CM|Malignant neoplasm of appendix vermiformis|Malignant neoplasm of appendix vermiformis
C0153439|T191|AB|153.6|ICD9CM|Malig neo ascend colon|Malig neo ascend colon
C0153439|T191|PT|153.6|ICD9CM|Malignant neoplasm of ascending colon|Malignant neoplasm of ascending colon
C0153440|T191|AB|153.7|ICD9CM|Mal neo splenic flexure|Mal neo splenic flexure
C0153440|T191|PT|153.7|ICD9CM|Malignant neoplasm of splenic flexure|Malignant neoplasm of splenic flexure
C0153441|T191|AB|153.8|ICD9CM|Malignant neo colon NEC|Malignant neo colon NEC
C0153441|T191|PT|153.8|ICD9CM|Malignant neoplasm of other specified sites of large intestine|Malignant neoplasm of other specified sites of large intestine
C0007102|T191|AB|153.9|ICD9CM|Malignant neo colon NOS|Malignant neo colon NOS
C0007102|T191|PT|153.9|ICD9CM|Malignant neoplasm of colon, unspecified site|Malignant neoplasm of colon, unspecified site
C0153442|T191|HT|154|ICD9CM|Malignant neoplasm of rectum, rectosigmoid junction, and anus|Malignant neoplasm of rectum, rectosigmoid junction, and anus
C0153443|T191|AB|154.0|ICD9CM|Mal neo rectosigmoid jct|Mal neo rectosigmoid jct
C0153443|T191|PT|154.0|ICD9CM|Malignant neoplasm of rectosigmoid junction|Malignant neoplasm of rectosigmoid junction
C0949022|T191|AB|154.1|ICD9CM|Malignant neopl rectum|Malignant neopl rectum
C0949022|T191|PT|154.1|ICD9CM|Malignant neoplasm of rectum|Malignant neoplasm of rectum
C0153445|T191|AB|154.2|ICD9CM|Malig neopl anal canal|Malig neopl anal canal
C0153445|T191|PT|154.2|ICD9CM|Malignant neoplasm of anal canal|Malignant neoplasm of anal canal
C0153446|T191|AB|154.3|ICD9CM|Malignant neo anus NOS|Malignant neo anus NOS
C0153446|T191|PT|154.3|ICD9CM|Malignant neoplasm of anus, unspecified site|Malignant neoplasm of anus, unspecified site
C0153447|T191|AB|154.8|ICD9CM|Mal neo rectum/anus NEC|Mal neo rectum/anus NEC
C0153447|T191|PT|154.8|ICD9CM|Malignant neoplasm of other sites of rectum, rectosigmoid junction, and anus|Malignant neoplasm of other sites of rectum, rectosigmoid junction, and anus
C0153448|T191|HT|155|ICD9CM|Malignant neoplasm of liver and intrahepatic bile ducts|Malignant neoplasm of liver and intrahepatic bile ducts
C0024620|T191|AB|155.0|ICD9CM|Mal neo liver, primary|Mal neo liver, primary
C0024620|T191|PT|155.0|ICD9CM|Malignant neoplasm of liver, primary|Malignant neoplasm of liver, primary
C0546835|T191|AB|155.1|ICD9CM|Mal neo intrahepat ducts|Mal neo intrahepat ducts
C0546835|T191|PT|155.1|ICD9CM|Malignant neoplasm of intrahepatic bile ducts|Malignant neoplasm of intrahepatic bile ducts
C0345904|T191|AB|155.2|ICD9CM|Malignant neo liver NOS|Malignant neo liver NOS
C0345904|T191|PT|155.2|ICD9CM|Malignant neoplasm of liver, not specified as primary or secondary|Malignant neoplasm of liver, not specified as primary or secondary
C1306605|T191|HT|156|ICD9CM|Malignant neoplasm of gallbladder and extrahepatic bile ducts|Malignant neoplasm of gallbladder and extrahepatic bile ducts
C0153452|T191|AB|156.0|ICD9CM|Malig neo gallbladder|Malig neo gallbladder
C0153452|T191|PT|156.0|ICD9CM|Malignant neoplasm of gallbladder|Malignant neoplasm of gallbladder
C0153453|T191|AB|156.1|ICD9CM|Mal neo extrahepat ducts|Mal neo extrahepat ducts
C0153453|T191|PT|156.1|ICD9CM|Malignant neoplasm of extrahepatic bile ducts|Malignant neoplasm of extrahepatic bile ducts
C0153454|T191|AB|156.2|ICD9CM|Mal neo ampulla of vater|Mal neo ampulla of vater
C0153454|T191|PT|156.2|ICD9CM|Malignant neoplasm of ampulla of vater|Malignant neoplasm of ampulla of vater
C0153455|T191|AB|156.8|ICD9CM|Malig neo biliary NEC|Malig neo biliary NEC
C0153455|T191|PT|156.8|ICD9CM|Malignant neoplasm of other specified sites of gallbladder and extrahepatic bile ducts|Malignant neoplasm of other specified sites of gallbladder and extrahepatic bile ducts
C0750952|T191|AB|156.9|ICD9CM|Malig neo biliary NOS|Malig neo biliary NOS
C0750952|T191|PT|156.9|ICD9CM|Malignant neoplasm of biliary tract, part unspecified site|Malignant neoplasm of biliary tract, part unspecified site
C0346647|T191|HT|157|ICD9CM|Malignant neoplasm of pancreas|Malignant neoplasm of pancreas
C0153458|T191|AB|157.0|ICD9CM|Mal neo pancreas head|Mal neo pancreas head
C0153458|T191|PT|157.0|ICD9CM|Malignant neoplasm of head of pancreas|Malignant neoplasm of head of pancreas
C0153459|T191|AB|157.1|ICD9CM|Mal neo pancreas body|Mal neo pancreas body
C0153459|T191|PT|157.1|ICD9CM|Malignant neoplasm of body of pancreas|Malignant neoplasm of body of pancreas
C0153460|T191|AB|157.2|ICD9CM|Mal neo pancreas tail|Mal neo pancreas tail
C0153460|T191|PT|157.2|ICD9CM|Malignant neoplasm of tail of pancreas|Malignant neoplasm of tail of pancreas
C0153461|T191|AB|157.3|ICD9CM|Mal neo pancreatic duct|Mal neo pancreatic duct
C0153461|T191|PT|157.3|ICD9CM|Malignant neoplasm of pancreatic duct|Malignant neoplasm of pancreatic duct
C1328479|T191|AB|157.4|ICD9CM|Mal neo islet langerhans|Mal neo islet langerhans
C1328479|T191|PT|157.4|ICD9CM|Malignant neoplasm of islets of langerhans|Malignant neoplasm of islets of langerhans
C0153463|T191|AB|157.8|ICD9CM|Malig neo pancreas NEC|Malig neo pancreas NEC
C0153463|T191|PT|157.8|ICD9CM|Malignant neoplasm of other specified sites of pancreas|Malignant neoplasm of other specified sites of pancreas
C0346647|T191|AB|157.9|ICD9CM|Malig neo pancreas NOS|Malig neo pancreas NOS
C0346647|T191|PT|157.9|ICD9CM|Malignant neoplasm of pancreas, part unspecified|Malignant neoplasm of pancreas, part unspecified
C0153464|T191|HT|158|ICD9CM|Malignant neoplasm of retroperitoneum and peritoneum|Malignant neoplasm of retroperitoneum and peritoneum
C0153465|T191|AB|158.0|ICD9CM|Mal neo retroperitoneum|Mal neo retroperitoneum
C0153465|T191|PT|158.0|ICD9CM|Malignant neoplasm of retroperitoneum|Malignant neoplasm of retroperitoneum
C0153466|T191|AB|158.8|ICD9CM|Mal neo peritoneum NEC|Mal neo peritoneum NEC
C0153466|T191|PT|158.8|ICD9CM|Malignant neoplasm of specified parts of peritoneum|Malignant neoplasm of specified parts of peritoneum
C0153467|T191|AB|158.9|ICD9CM|Mal neo peritoneum NOS|Mal neo peritoneum NOS
C0153467|T191|PT|158.9|ICD9CM|Malignant neoplasm of peritoneum, unspecified|Malignant neoplasm of peritoneum, unspecified
C0153468|T191|HT|159|ICD9CM|Malignant neoplasm of other and ill-defined sites within the digestive organs and peritoneum|Malignant neoplasm of other and ill-defined sites within the digestive organs and peritoneum
C0346627|T191|AB|159.0|ICD9CM|Malig neo intestine NOS|Malig neo intestine NOS
C0346627|T191|PT|159.0|ICD9CM|Malignant neoplasm of intestinal tract, part unspecified|Malignant neoplasm of intestinal tract, part unspecified
C0869278|T191|AB|159.1|ICD9CM|Malignant neo spleen NEC|Malignant neo spleen NEC
C0869278|T191|PT|159.1|ICD9CM|Malignant neoplasm of spleen, not elsewhere classified|Malignant neoplasm of spleen, not elsewhere classified
C0153471|T191|AB|159.8|ICD9CM|Mal neo gi/intra-abd NEC|Mal neo gi/intra-abd NEC
C0153471|T191|PT|159.8|ICD9CM|Malignant neoplasm of other sites of digestive system and intra-abdominal organs|Malignant neoplasm of other sites of digestive system and intra-abdominal organs
C0153472|T191|AB|159.9|ICD9CM|Mal neo GI tract ill-def|Mal neo GI tract ill-def
C0153472|T191|PT|159.9|ICD9CM|Malignant neoplasm of ill-defined sites within the digestive organs and peritoneum|Malignant neoplasm of ill-defined sites within the digestive organs and peritoneum
C0153473|T191|HT|160|ICD9CM|Malignant neoplasm of nasal cavities, middle ear, and accessory sinuses|Malignant neoplasm of nasal cavities, middle ear, and accessory sinuses
C0178249|T191|HT|160-165.99|ICD9CM|MALIGNANT NEOPLASM OF RESPIRATORY AND INTRATHORACIC ORGANS|MALIGNANT NEOPLASM OF RESPIRATORY AND INTRATHORACIC ORGANS
C0728864|T191|AB|160.0|ICD9CM|Mal neo nasal cavities|Mal neo nasal cavities
C0728864|T191|PT|160.0|ICD9CM|Malignant neoplasm of nasal cavities|Malignant neoplasm of nasal cavities
C0153475|T191|AB|160.1|ICD9CM|Malig neo middle ear|Malig neo middle ear
C0153475|T191|PT|160.1|ICD9CM|Malignant neoplasm of auditory tube, middle ear, and mastoid air cells|Malignant neoplasm of auditory tube, middle ear, and mastoid air cells
C0153476|T191|AB|160.2|ICD9CM|Mal neo maxillary sinus|Mal neo maxillary sinus
C0153476|T191|PT|160.2|ICD9CM|Malignant neoplasm of maxillary sinus|Malignant neoplasm of maxillary sinus
C0153477|T191|AB|160.3|ICD9CM|Mal neo ethmoidal sinus|Mal neo ethmoidal sinus
C0153477|T191|PT|160.3|ICD9CM|Malignant neoplasm of ethmoidal sinus|Malignant neoplasm of ethmoidal sinus
C0153478|T191|AB|160.4|ICD9CM|Malig neo frontal sinus|Malig neo frontal sinus
C0153478|T191|PT|160.4|ICD9CM|Malignant neoplasm of frontal sinus|Malignant neoplasm of frontal sinus
C0153479|T191|AB|160.5|ICD9CM|Mal neo sphenoid sinus|Mal neo sphenoid sinus
C0153479|T191|PT|160.5|ICD9CM|Malignant neoplasm of sphenoidal sinus|Malignant neoplasm of sphenoidal sinus
C0153480|T191|AB|160.8|ICD9CM|Mal neo access sinus NEC|Mal neo access sinus NEC
C0153480|T191|PT|160.8|ICD9CM|Malignant neoplasm of other accessory sinuses|Malignant neoplasm of other accessory sinuses
C0153474|T191|AB|160.9|ICD9CM|Mal neo access sinus NOS|Mal neo access sinus NOS
C0153474|T191|PT|160.9|ICD9CM|Malignant neoplasm of accessory sinus, unspecified|Malignant neoplasm of accessory sinus, unspecified
C0007107|T191|HT|161|ICD9CM|Malignant neoplasm of larynx|Malignant neoplasm of larynx
C0153483|T191|AB|161.0|ICD9CM|Malignant neo glottis|Malignant neo glottis
C0153483|T191|PT|161.0|ICD9CM|Malignant neoplasm of glottis|Malignant neoplasm of glottis
C0153484|T191|AB|161.1|ICD9CM|Malig neo supraglottis|Malig neo supraglottis
C0153484|T191|PT|161.1|ICD9CM|Malignant neoplasm of supraglottis|Malignant neoplasm of supraglottis
C0153485|T191|AB|161.2|ICD9CM|Malig neo subglottis|Malig neo subglottis
C0153485|T191|PT|161.2|ICD9CM|Malignant neoplasm of subglottis|Malignant neoplasm of subglottis
C0153486|T191|AB|161.3|ICD9CM|Mal neo cartilage larynx|Mal neo cartilage larynx
C0153486|T191|PT|161.3|ICD9CM|Malignant neoplasm of laryngeal cartilages|Malignant neoplasm of laryngeal cartilages
C0153487|T191|AB|161.8|ICD9CM|Malignant neo larynx NEC|Malignant neo larynx NEC
C0153487|T191|PT|161.8|ICD9CM|Malignant neoplasm of other specified sites of larynx|Malignant neoplasm of other specified sites of larynx
C0007107|T191|AB|161.9|ICD9CM|Malignant neo larynx NOS|Malignant neo larynx NOS
C0007107|T191|PT|161.9|ICD9CM|Malignant neoplasm of larynx, unspecified|Malignant neoplasm of larynx, unspecified
C0153488|T191|HT|162|ICD9CM|Malignant neoplasm of trachea, bronchus, and lung|Malignant neoplasm of trachea, bronchus, and lung
C0153489|T191|AB|162.0|ICD9CM|Malignant neo trachea|Malignant neo trachea
C0153489|T191|PT|162.0|ICD9CM|Malignant neoplasm of trachea|Malignant neoplasm of trachea
C0153490|T191|AB|162.2|ICD9CM|Malig neo main bronchus|Malig neo main bronchus
C0153490|T191|PT|162.2|ICD9CM|Malignant neoplasm of main bronchus|Malignant neoplasm of main bronchus
C0024624|T191|AB|162.3|ICD9CM|Mal neo upper lobe lung|Mal neo upper lobe lung
C0024624|T191|PT|162.3|ICD9CM|Malignant neoplasm of upper lobe, bronchus or lung|Malignant neoplasm of upper lobe, bronchus or lung
C0153491|T191|AB|162.4|ICD9CM|Mal neo middle lobe lung|Mal neo middle lobe lung
C0153491|T191|PT|162.4|ICD9CM|Malignant neoplasm of middle lobe, bronchus or lung|Malignant neoplasm of middle lobe, bronchus or lung
C0153492|T191|AB|162.5|ICD9CM|Mal neo lower lobe lung|Mal neo lower lobe lung
C0153492|T191|PT|162.5|ICD9CM|Malignant neoplasm of lower lobe, bronchus or lung|Malignant neoplasm of lower lobe, bronchus or lung
C0153493|T191|AB|162.8|ICD9CM|Mal neo bronch/lung NEC|Mal neo bronch/lung NEC
C0153493|T191|PT|162.8|ICD9CM|Malignant neoplasm of other parts of bronchus or lung|Malignant neoplasm of other parts of bronchus or lung
C0348343|T191|AB|162.9|ICD9CM|Mal neo bronch/lung NOS|Mal neo bronch/lung NOS
C0348343|T191|PT|162.9|ICD9CM|Malignant neoplasm of bronchus and lung, unspecified|Malignant neoplasm of bronchus and lung, unspecified
C0153494|T191|HT|163|ICD9CM|Malignant neoplasm of pleura|Malignant neoplasm of pleura
C2004481|T191|AB|163.0|ICD9CM|Mal neo parietal pleura|Mal neo parietal pleura
C2004481|T191|PT|163.0|ICD9CM|Malignant neoplasm of parietal pleura|Malignant neoplasm of parietal pleura
C2607950|T191|AB|163.1|ICD9CM|Mal neo visceral pleura|Mal neo visceral pleura
C2607950|T191|PT|163.1|ICD9CM|Malignant neoplasm of visceral pleura|Malignant neoplasm of visceral pleura
C0153497|T191|AB|163.8|ICD9CM|Malig neopl pleura NEC|Malig neopl pleura NEC
C0153497|T191|PT|163.8|ICD9CM|Malignant neoplasm of other specified sites of pleura|Malignant neoplasm of other specified sites of pleura
C0153494|T191|AB|163.9|ICD9CM|Malig neopl pleura NOS|Malig neopl pleura NOS
C0153494|T191|PT|163.9|ICD9CM|Malignant neoplasm of pleura, unspecified|Malignant neoplasm of pleura, unspecified
C0153498|T191|HT|164|ICD9CM|Malignant neoplasm of thymus, heart, and mediastinum|Malignant neoplasm of thymus, heart, and mediastinum
C0751552|T191|AB|164.0|ICD9CM|Malignant neopl thymus|Malignant neopl thymus
C0751552|T191|PT|164.0|ICD9CM|Malignant neoplasm of thymus|Malignant neoplasm of thymus
C0153500|T191|AB|164.1|ICD9CM|Malignant neopl heart|Malignant neopl heart
C0153500|T191|PT|164.1|ICD9CM|Malignant neoplasm of heart|Malignant neoplasm of heart
C0153501|T191|AB|164.2|ICD9CM|Mal neo ant mediastinum|Mal neo ant mediastinum
C0153501|T191|PT|164.2|ICD9CM|Malignant neoplasm of anterior mediastinum|Malignant neoplasm of anterior mediastinum
C0153502|T191|AB|164.3|ICD9CM|Mal neo post mediastinum|Mal neo post mediastinum
C0153502|T191|PT|164.3|ICD9CM|Malignant neoplasm of posterior mediastinum|Malignant neoplasm of posterior mediastinum
C0153503|T191|AB|164.8|ICD9CM|Mal neo mediastinum NEC|Mal neo mediastinum NEC
C0153503|T191|PT|164.8|ICD9CM|Malignant neoplasm of other parts of mediastinum|Malignant neoplasm of other parts of mediastinum
C0153504|T191|AB|164.9|ICD9CM|Mal neo mediastinum NOS|Mal neo mediastinum NOS
C0153504|T191|PT|164.9|ICD9CM|Malignant neoplasm of mediastinum, part unspecified|Malignant neoplasm of mediastinum, part unspecified
C0153506|T191|AB|165.0|ICD9CM|Mal neo upper resp NOS|Mal neo upper resp NOS
C0153506|T191|PT|165.0|ICD9CM|Malignant neoplasm of upper respiratory tract, part unspecified|Malignant neoplasm of upper respiratory tract, part unspecified
C0153507|T191|AB|165.8|ICD9CM|Mal neo thorax/resp NEC|Mal neo thorax/resp NEC
C0153507|T191|PT|165.8|ICD9CM|Malignant neoplasm of other sites within the respiratory system and intrathoracic organs|Malignant neoplasm of other sites within the respiratory system and intrathoracic organs
C0153508|T191|AB|165.9|ICD9CM|Mal neo resp system NOS|Mal neo resp system NOS
C0153508|T191|PT|165.9|ICD9CM|Malignant neoplasm of ill-defined sites within the respiratory system|Malignant neoplasm of ill-defined sites within the respiratory system
C0153509|T191|HT|170|ICD9CM|Malignant neoplasm of bone and articular cartilage|Malignant neoplasm of bone and articular cartilage
C0178250|T191|HT|170-176.99|ICD9CM|MALIGNANT NEOPLASM OF BONE, CONNECTIVE TISSUE, SKIN, AND BREAST|MALIGNANT NEOPLASM OF BONE, CONNECTIVE TISSUE, SKIN, AND BREAST
C0153510|T191|AB|170.0|ICD9CM|Mal neo skull/face bone|Mal neo skull/face bone
C0153510|T191|PT|170.0|ICD9CM|Malignant neoplasm of bones of skull and face, except mandible|Malignant neoplasm of bones of skull and face, except mandible
C0153511|T191|AB|170.1|ICD9CM|Malignant neo mandible|Malignant neo mandible
C0153511|T191|PT|170.1|ICD9CM|Malignant neoplasm of mandible|Malignant neoplasm of mandible
C0153512|T191|AB|170.2|ICD9CM|Malig neo vertebrae|Malig neo vertebrae
C0153512|T191|PT|170.2|ICD9CM|Malignant neoplasm of vertebral column, excluding sacrum and coccyx|Malignant neoplasm of vertebral column, excluding sacrum and coccyx
C0153513|T191|AB|170.3|ICD9CM|Mal neo ribs/stern/clav|Mal neo ribs/stern/clav
C0153513|T191|PT|170.3|ICD9CM|Malignant neoplasm of ribs, sternum, and clavicle|Malignant neoplasm of ribs, sternum, and clavicle
C0153514|T191|AB|170.4|ICD9CM|Mal neo long bones arm|Mal neo long bones arm
C0153514|T191|PT|170.4|ICD9CM|Malignant neoplasm of scapula and long bones of upper limb|Malignant neoplasm of scapula and long bones of upper limb
C0153515|T191|AB|170.5|ICD9CM|Mal neo bones wrist/hand|Mal neo bones wrist/hand
C0153515|T191|PT|170.5|ICD9CM|Malignant neoplasm of short bones of upper limb|Malignant neoplasm of short bones of upper limb
C0153516|T191|AB|170.6|ICD9CM|Mal neo pelvic girdle|Mal neo pelvic girdle
C0153516|T191|PT|170.6|ICD9CM|Malignant neoplasm of pelvic bones, sacrum, and coccyx|Malignant neoplasm of pelvic bones, sacrum, and coccyx
C0153517|T191|AB|170.7|ICD9CM|Mal neo long bones leg|Mal neo long bones leg
C0153517|T191|PT|170.7|ICD9CM|Malignant neoplasm of long bones of lower limb|Malignant neoplasm of long bones of lower limb
C0153518|T191|AB|170.8|ICD9CM|Mal neo bones ankle/foot|Mal neo bones ankle/foot
C0153518|T191|PT|170.8|ICD9CM|Malignant neoplasm of short bones of lower limb|Malignant neoplasm of short bones of lower limb
C0153509|T191|AB|170.9|ICD9CM|Malig neopl bone NOS|Malig neopl bone NOS
C0153509|T191|PT|170.9|ICD9CM|Malignant neoplasm of bone and articular cartilage, site unspecified|Malignant neoplasm of bone and articular cartilage, site unspecified
C0153519|T191|HT|171|ICD9CM|Malignant neoplasm of connective and other soft tissue|Malignant neoplasm of connective and other soft tissue
C0153520|T191|AB|171.0|ICD9CM|Mal neo soft tissue head|Mal neo soft tissue head
C0153520|T191|PT|171.0|ICD9CM|Malignant neoplasm of connective and other soft tissue of head, face, and neck|Malignant neoplasm of connective and other soft tissue of head, face, and neck
C0153521|T191|AB|171.2|ICD9CM|Mal neo soft tissue arm|Mal neo soft tissue arm
C0153521|T191|PT|171.2|ICD9CM|Malignant neoplasm of connective and other soft tissue of upper limb, including shoulder|Malignant neoplasm of connective and other soft tissue of upper limb, including shoulder
C0153522|T191|AB|171.3|ICD9CM|Mal neo soft tissue leg|Mal neo soft tissue leg
C0153522|T191|PT|171.3|ICD9CM|Malignant neoplasm of connective and other soft tissue of lower limb, including hip|Malignant neoplasm of connective and other soft tissue of lower limb, including hip
C0153523|T191|AB|171.4|ICD9CM|Mal neo soft tis thorax|Mal neo soft tis thorax
C0153523|T191|PT|171.4|ICD9CM|Malignant neoplasm of connective and other soft tissue of thorax|Malignant neoplasm of connective and other soft tissue of thorax
C0153524|T191|AB|171.5|ICD9CM|Mal neo soft tis abdomen|Mal neo soft tis abdomen
C0153524|T191|PT|171.5|ICD9CM|Malignant neoplasm of connective and other soft tissue of abdomen|Malignant neoplasm of connective and other soft tissue of abdomen
C0153525|T191|AB|171.6|ICD9CM|Mal neo soft tis pelvis|Mal neo soft tis pelvis
C0153525|T191|PT|171.6|ICD9CM|Malignant neoplasm of connective and other soft tissue of pelvis|Malignant neoplasm of connective and other soft tissue of pelvis
C0375065|T191|AB|171.7|ICD9CM|Mal neopl trunk NOS|Mal neopl trunk NOS
C0375065|T191|PT|171.7|ICD9CM|Malignant neoplasm of connective and other soft tissue of trunk, unspecified|Malignant neoplasm of connective and other soft tissue of trunk, unspecified
C0153527|T191|AB|171.8|ICD9CM|Mal neo soft tissue NEC|Mal neo soft tissue NEC
C0153527|T191|PT|171.8|ICD9CM|Malignant neoplasm of other specified sites of connective and other soft tissue|Malignant neoplasm of other specified sites of connective and other soft tissue
C0153519|T191|AB|171.9|ICD9CM|Mal neo soft tissue NOS|Mal neo soft tissue NOS
C0153519|T191|PT|171.9|ICD9CM|Malignant neoplasm of connective and other soft tissue, site unspecified|Malignant neoplasm of connective and other soft tissue, site unspecified
C0151779|T191|HT|172|ICD9CM|Malignant melanoma of skin|Malignant melanoma of skin
C0153529|T191|AB|172.0|ICD9CM|Malig melanoma lip|Malig melanoma lip
C0153529|T191|PT|172.0|ICD9CM|Malignant melanoma of skin of lip|Malignant melanoma of skin of lip
C3665588|T191|AB|172.1|ICD9CM|Malig melanoma eyelid|Malig melanoma eyelid
C3665588|T191|PT|172.1|ICD9CM|Malignant melanoma of skin of eyelid, including canthus|Malignant melanoma of skin of eyelid, including canthus
C0346773|T191|AB|172.2|ICD9CM|Malig melanoma ear|Malig melanoma ear
C0346773|T191|PT|172.2|ICD9CM|Malignant melanoma of skin of ear and external auditory canal|Malignant melanoma of skin of ear and external auditory canal
C0153532|T191|AB|172.3|ICD9CM|Mal melanom face NEC/NOS|Mal melanom face NEC/NOS
C0153532|T191|PT|172.3|ICD9CM|Malignant melanoma of skin of other and unspecified parts of face|Malignant melanoma of skin of other and unspecified parts of face
C0346782|T191|AB|172.4|ICD9CM|Mal melanoma scalp/neck|Mal melanoma scalp/neck
C0346782|T191|PT|172.4|ICD9CM|Malignant melanoma of skin of scalp and neck|Malignant melanoma of skin of scalp and neck
C1112782|T191|AB|172.5|ICD9CM|Malig melanoma trunk|Malig melanoma trunk
C1112782|T191|PT|172.5|ICD9CM|Malignant melanoma of skin of trunk, except scrotum|Malignant melanoma of skin of trunk, except scrotum
C1112533|T191|AB|172.6|ICD9CM|Malig melanoma arm|Malig melanoma arm
C1112533|T191|PT|172.6|ICD9CM|Malignant melanoma of skin of upper limb, including shoulder|Malignant melanoma of skin of upper limb, including shoulder
C1112532|T191|AB|172.7|ICD9CM|Malig melanoma leg|Malig melanoma leg
C1112532|T191|PT|172.7|ICD9CM|Malignant melanoma of skin of lower limb, including hip|Malignant melanoma of skin of lower limb, including hip
C0153537|T191|AB|172.8|ICD9CM|Malig melanoma skin NEC|Malig melanoma skin NEC
C0153537|T191|PT|172.8|ICD9CM|Malignant melanoma of other specified sites of skin|Malignant melanoma of other specified sites of skin
C0151779|T191|AB|172.9|ICD9CM|Malig melanoma skin NOS|Malig melanoma skin NOS
C0151779|T191|PT|172.9|ICD9CM|Melanoma of skin, site unspecified|Melanoma of skin, site unspecified
C3161362|T191|HT|173|ICD9CM|Other and unspecified malignant neoplasm of skin|Other and unspecified malignant neoplasm of skin
C0153539|T191|HT|173.0|ICD9CM|Other malignant neoplasm of skin of lip|Other malignant neoplasm of skin of lip
C3161037|T191|AB|173.00|ICD9CM|Malig neopl skin lip NOS|Malig neopl skin lip NOS
C3161037|T191|PT|173.00|ICD9CM|Unspecified malignant neoplasm of skin of lip|Unspecified malignant neoplasm of skin of lip
C1274259|T191|AB|173.01|ICD9CM|Basal cell ca skin lip|Basal cell ca skin lip
C1274259|T191|PT|173.01|ICD9CM|Basal cell carcinoma of skin of lip|Basal cell carcinoma of skin of lip
C3161038|T191|AB|173.02|ICD9CM|Squamous cell ca skn lip|Squamous cell ca skn lip
C3161038|T191|PT|173.02|ICD9CM|Squamous cell carcinoma of skin of lip|Squamous cell carcinoma of skin of lip
C3161039|T191|AB|173.09|ICD9CM|Malig neo skin lip NEC|Malig neo skin lip NEC
C3161039|T191|PT|173.09|ICD9CM|Other specified malignant neoplasm of skin of lip|Other specified malignant neoplasm of skin of lip
C3161363|T191|HT|173.1|ICD9CM|Other and unspecified malignant neoplasm of skin of eyelid, including canthus|Other and unspecified malignant neoplasm of skin of eyelid, including canthus
C3161040|T191|AB|173.10|ICD9CM|Mal neo eyelid/canth NOS|Mal neo eyelid/canth NOS
C3161040|T191|PT|173.10|ICD9CM|Unspecified malignant neoplasm of eyelid, including canthus|Unspecified malignant neoplasm of eyelid, including canthus
C3161041|T191|AB|173.11|ICD9CM|Basal cell ca lid/canth|Basal cell ca lid/canth
C3161041|T191|PT|173.11|ICD9CM|Basal cell carcinoma of eyelid, including canthus|Basal cell carcinoma of eyelid, including canthus
C3161042|T191|AB|173.12|ICD9CM|Squam cell ca lid/canth|Squam cell ca lid/canth
C3161042|T191|PT|173.12|ICD9CM|Squamous cell carcinoma of eyelid, including canthus|Squamous cell carcinoma of eyelid, including canthus
C3161043|T191|AB|173.19|ICD9CM|Mal neo eyelid/canth NEC|Mal neo eyelid/canth NEC
C3161043|T191|PT|173.19|ICD9CM|Other specified malignant neoplasm of eyelid, including canthus|Other specified malignant neoplasm of eyelid, including canthus
C3161364|T191|HT|173.2|ICD9CM|Other and unspecified malignant neoplasm of skin of ear and external auditory canal|Other and unspecified malignant neoplasm of skin of ear and external auditory canal
C3161044|T191|AB|173.20|ICD9CM|Malig neo skin ear NOS|Malig neo skin ear NOS
C3161044|T191|PT|173.20|ICD9CM|Unspecified malignant neoplasm of skin of ear and external auditory canal|Unspecified malignant neoplasm of skin of ear and external auditory canal
C3161045|T191|AB|173.21|ICD9CM|Basal cell ca skin ear|Basal cell ca skin ear
C3161045|T191|PT|173.21|ICD9CM|Basal cell carcinoma of skin of ear and external auditory canal|Basal cell carcinoma of skin of ear and external auditory canal
C3161046|T191|AB|173.22|ICD9CM|Squam cell ca skin ear|Squam cell ca skin ear
C3161046|T191|PT|173.22|ICD9CM|Squamous cell carcinoma of skin of ear and external auditory canal|Squamous cell carcinoma of skin of ear and external auditory canal
C3161047|T191|AB|173.29|ICD9CM|Neo skin ear/ex canl NEC|Neo skin ear/ex canl NEC
C3161047|T191|PT|173.29|ICD9CM|Other specified malignant neoplasm of skin of ear and external auditory canal|Other specified malignant neoplasm of skin of ear and external auditory canal
C3161365|T191|HT|173.3|ICD9CM|Other and unspecified malignant neoplasm of skin of other and unspecified parts of face|Other and unspecified malignant neoplasm of skin of other and unspecified parts of face
C3161048|T047|AB|173.30|ICD9CM|Mal neo skn face NEC/NOS|Mal neo skn face NEC/NOS
C3161048|T047|PT|173.30|ICD9CM|Unspecified malignant neoplasm of skin of other and unspecified parts of face|Unspecified malignant neoplasm of skin of other and unspecified parts of face
C3161049|T191|PT|173.31|ICD9CM|Basal cell carcinoma of skin of other and unspecified parts of face|Basal cell carcinoma of skin of other and unspecified parts of face
C3161049|T191|AB|173.31|ICD9CM|Bsl cel skn face NEC/NOS|Bsl cel skn face NEC/NOS
C3161050|T191|AB|173.32|ICD9CM|Sqm cel skn face NEC/NOS|Sqm cel skn face NEC/NOS
C3161050|T191|PT|173.32|ICD9CM|Squamous cell carcinoma of skin of other and unspecified parts of face|Squamous cell carcinoma of skin of other and unspecified parts of face
C3161048|T047|AB|173.39|ICD9CM|Mal neo skn face NEC/NOS|Mal neo skn face NEC/NOS
C3161048|T047|PT|173.39|ICD9CM|Other specified malignant neoplasm of skin of other and unspecified parts of face|Other specified malignant neoplasm of skin of other and unspecified parts of face
C3161366|T191|HT|173.4|ICD9CM|Other and unspecified malignant neoplasm of scalp and skin of neck|Other and unspecified malignant neoplasm of scalp and skin of neck
C3161051|T191|AB|173.40|ICD9CM|Mal neo sclp/skn nck NOS|Mal neo sclp/skn nck NOS
C3161051|T191|PT|173.40|ICD9CM|Unspecified malignant neoplasm of scalp and skin of neck|Unspecified malignant neoplasm of scalp and skin of neck
C3161052|T191|PT|173.41|ICD9CM|Basal cell carcinoma of scalp and skin of neck|Basal cell carcinoma of scalp and skin of neck
C3161052|T191|AB|173.41|ICD9CM|Bsl cell ca scalp/skn nk|Bsl cell ca scalp/skn nk
C3161053|T191|AB|173.42|ICD9CM|Sqam cell ca sclp/skn nk|Sqam cell ca sclp/skn nk
C3161053|T191|PT|173.42|ICD9CM|Squamous cell carcinoma of scalp and skin of neck|Squamous cell carcinoma of scalp and skin of neck
C3161054|T191|AB|173.49|ICD9CM|Mal neo sclp/skn nck NEC|Mal neo sclp/skn nck NEC
C3161054|T191|PT|173.49|ICD9CM|Other specified malignant neoplasm of scalp and skin of neck|Other specified malignant neoplasm of scalp and skin of neck
C3161367|T191|HT|173.5|ICD9CM|Other and unspecified malignant neoplasm of skin of trunk, except scrotum|Other and unspecified malignant neoplasm of skin of trunk, except scrotum
C3161055|T191|AB|173.50|ICD9CM|Malig neo skin trunk NOS|Malig neo skin trunk NOS
C3161055|T191|PT|173.50|ICD9CM|Unspecified malignant neoplasm of skin of trunk, except scrotum|Unspecified malignant neoplasm of skin of trunk, except scrotum
C3161056|T191|AB|173.51|ICD9CM|Basal cell ca skin trunk|Basal cell ca skin trunk
C3161056|T191|PT|173.51|ICD9CM|Basal cell carcinoma of skin of trunk, except scrotum|Basal cell carcinoma of skin of trunk, except scrotum
C3161057|T191|AB|173.52|ICD9CM|Squam cell ca skin trunk|Squam cell ca skin trunk
C3161057|T191|PT|173.52|ICD9CM|Squamous cell carcinoma of skin of trunk, except scrotum|Squamous cell carcinoma of skin of trunk, except scrotum
C3161058|T191|AB|173.59|ICD9CM|Malig neo skin trunk NEC|Malig neo skin trunk NEC
C3161058|T191|PT|173.59|ICD9CM|Other specified malignant neoplasm of skin of trunk, except scrotum|Other specified malignant neoplasm of skin of trunk, except scrotum
C3161368|T191|HT|173.6|ICD9CM|Other and unspecified malignant neoplasm of skin of upper limb, including shoulder|Other and unspecified malignant neoplasm of skin of upper limb, including shoulder
C2838014|T191|AB|173.60|ICD9CM|Mal neo skin up limb NOS|Mal neo skin up limb NOS
C2838014|T191|PT|173.60|ICD9CM|Unspecified malignant neoplasm of skin of upper limb, including shoulder|Unspecified malignant neoplasm of skin of upper limb, including shoulder
C3161059|T191|AB|173.61|ICD9CM|Basal cell ca skn up lmb|Basal cell ca skn up lmb
C3161059|T191|PT|173.61|ICD9CM|Basal cell carcinoma of skin of upper limb, including shoulder|Basal cell carcinoma of skin of upper limb, including shoulder
C3161060|T191|AB|173.62|ICD9CM|Squam cell ca skn up lmb|Squam cell ca skn up lmb
C3161060|T191|PT|173.62|ICD9CM|Squamous cell carcinoma of skin of upper limb, including shoulder|Squamous cell carcinoma of skin of upper limb, including shoulder
C3161061|T191|AB|173.69|ICD9CM|Malig neo skn up lmb NEC|Malig neo skn up lmb NEC
C3161061|T191|PT|173.69|ICD9CM|Other specified malignant neoplasm of skin of upper limb, including shoulder|Other specified malignant neoplasm of skin of upper limb, including shoulder
C3161369|T191|HT|173.7|ICD9CM|Other and unspecified malignant neoplasm of skin of lower limb, including hip|Other and unspecified malignant neoplasm of skin of lower limb, including hip
C2838017|T191|AB|173.70|ICD9CM|Mal neo skn low limb NOS|Mal neo skn low limb NOS
C2838017|T191|PT|173.70|ICD9CM|Unspecified malignant neoplasm of skin of lower limb, including hip|Unspecified malignant neoplasm of skin of lower limb, including hip
C3161062|T191|PT|173.71|ICD9CM|Basal cell carcinoma of skin of lower limb, including hip|Basal cell carcinoma of skin of lower limb, including hip
C3161062|T191|AB|173.71|ICD9CM|Basl cell ca skn low lmb|Basl cell ca skn low lmb
C3161063|T191|AB|173.72|ICD9CM|Sqam cell ca skn low lmb|Sqam cell ca skn low lmb
C3161063|T191|PT|173.72|ICD9CM|Squamous cell carcinoma of skin of lower limb, including hip|Squamous cell carcinoma of skin of lower limb, including hip
C3161064|T191|AB|173.79|ICD9CM|Mal neo skin low lmb NEC|Mal neo skin low lmb NEC
C3161064|T191|PT|173.79|ICD9CM|Other specified malignant neoplasm of skin of lower limb, including hip|Other specified malignant neoplasm of skin of lower limb, including hip
C3161370|T191|HT|173.8|ICD9CM|Other and unspecified malignant neoplasm of other specified sites of skin|Other and unspecified malignant neoplasm of other specified sites of skin
C3161065|T047|AB|173.80|ICD9CM|Mal neo skn site NEC/NOS|Mal neo skn site NEC/NOS
C3161065|T047|PT|173.80|ICD9CM|Unspecified malignant neoplasm of other specified sites of skin|Unspecified malignant neoplasm of other specified sites of skin
C3161066|T191|PT|173.81|ICD9CM|Basal cell carcinoma of other specified sites of skin|Basal cell carcinoma of other specified sites of skin
C3161066|T191|AB|173.81|ICD9CM|Bsl cell ca skn site NEC|Bsl cell ca skn site NEC
C3161067|T191|AB|173.82|ICD9CM|Sqm cell ca skn site NEC|Sqm cell ca skn site NEC
C3161067|T191|PT|173.82|ICD9CM|Squamous cell carcinoma of other specified sites of skin|Squamous cell carcinoma of other specified sites of skin
C3161068|T191|AB|173.89|ICD9CM|Oth mal neo skn site NEC|Oth mal neo skn site NEC
C3161068|T191|PT|173.89|ICD9CM|Other specified malignant neoplasm of other specified sites of skin|Other specified malignant neoplasm of other specified sites of skin
C3161371|T191|HT|173.9|ICD9CM|Other and unspecified malignant neoplasm of skin, site unspecified|Other and unspecified malignant neoplasm of skin, site unspecified
C3161069|T191|AB|173.90|ICD9CM|Malig neo skin site NOS|Malig neo skin site NOS
C3161069|T191|PT|173.90|ICD9CM|Unspecified malignant neoplasm of skin, site unspecified|Unspecified malignant neoplasm of skin, site unspecified
C3161070|T191|AB|173.91|ICD9CM|Basal cell ca skin NOS|Basal cell ca skin NOS
C3161070|T191|PT|173.91|ICD9CM|Basal cell carcinoma of skin, site unspecified|Basal cell carcinoma of skin, site unspecified
C3161071|T191|AB|173.92|ICD9CM|Squam cell ca skin NOS|Squam cell ca skin NOS
C3161071|T191|PT|173.92|ICD9CM|Squamous cell carcinoma of skin, site unspecified|Squamous cell carcinoma of skin, site unspecified
C3161065|T047|AB|173.99|ICD9CM|Oth mal neo skn site NOS|Oth mal neo skn site NOS
C3161065|T047|PT|173.99|ICD9CM|Other specified malignant neoplasm of skin, site unspecified|Other specified malignant neoplasm of skin, site unspecified
C0235653|T191|HT|174|ICD9CM|Malignant neoplasm of female breast|Malignant neoplasm of female breast
C0024621|T191|AB|174.0|ICD9CM|Malig neo nipple|Malig neo nipple
C0024621|T191|PT|174.0|ICD9CM|Malignant neoplasm of nipple and areola of female breast|Malignant neoplasm of nipple and areola of female breast
C0153549|T191|AB|174.1|ICD9CM|Mal neo breast-central|Mal neo breast-central
C0153549|T191|PT|174.1|ICD9CM|Malignant neoplasm of central portion of female breast|Malignant neoplasm of central portion of female breast
C0153550|T191|AB|174.2|ICD9CM|Mal neo breast up-inner|Mal neo breast up-inner
C0153550|T191|PT|174.2|ICD9CM|Malignant neoplasm of upper-inner quadrant of female breast|Malignant neoplasm of upper-inner quadrant of female breast
C0153551|T191|AB|174.3|ICD9CM|Mal neo breast low-inner|Mal neo breast low-inner
C0153551|T191|PT|174.3|ICD9CM|Malignant neoplasm of lower-inner quadrant of female breast|Malignant neoplasm of lower-inner quadrant of female breast
C0153552|T191|AB|174.4|ICD9CM|Mal neo breast up-outer|Mal neo breast up-outer
C0153552|T191|PT|174.4|ICD9CM|Malignant neoplasm of upper-outer quadrant of female breast|Malignant neoplasm of upper-outer quadrant of female breast
C0153553|T191|AB|174.5|ICD9CM|Mal neo breast low-outer|Mal neo breast low-outer
C0153553|T191|PT|174.5|ICD9CM|Malignant neoplasm of lower-outer quadrant of female breast|Malignant neoplasm of lower-outer quadrant of female breast
C0153554|T191|AB|174.6|ICD9CM|Mal neo breast-axillary|Mal neo breast-axillary
C0153554|T191|PT|174.6|ICD9CM|Malignant neoplasm of axillary tail of female breast|Malignant neoplasm of axillary tail of female breast
C0153555|T191|AB|174.8|ICD9CM|Malign neopl breast NEC|Malign neopl breast NEC
C0153555|T191|PT|174.8|ICD9CM|Malignant neoplasm of other specified sites of female breast|Malignant neoplasm of other specified sites of female breast
C0235653|T191|AB|174.9|ICD9CM|Malign neopl breast NOS|Malign neopl breast NOS
C0235653|T191|PT|174.9|ICD9CM|Malignant neoplasm of breast (female), unspecified|Malignant neoplasm of breast (female), unspecified
C0242787|T191|HT|175|ICD9CM|Malignant neoplasm of male breast|Malignant neoplasm of male breast
C0153558|T191|AB|175.0|ICD9CM|Mal neo male nipple|Mal neo male nipple
C0153558|T191|PT|175.0|ICD9CM|Malignant neoplasm of nipple and areola of male breast|Malignant neoplasm of nipple and areola of male breast
C0153559|T191|AB|175.9|ICD9CM|Mal neo male breast NEC|Mal neo male breast NEC
C0153559|T191|PT|175.9|ICD9CM|Malignant neoplasm of other and unspecified sites of male breast|Malignant neoplasm of other and unspecified sites of male breast
C0036220|T191|HT|176|ICD9CM|Kaposi's sarcoma|Kaposi's sarcoma
C0153560|T191|PT|176.0|ICD9CM|Kaposi's sarcoma, skin|Kaposi's sarcoma, skin
C0153560|T191|AB|176.0|ICD9CM|Skin - kaposi's sarcoma|Skin - kaposi's sarcoma
C0153561|T191|PT|176.1|ICD9CM|Kaposi's sarcoma, soft tissue|Kaposi's sarcoma, soft tissue
C0153561|T191|AB|176.1|ICD9CM|Sft tisue - kpsi's srcma|Sft tisue - kpsi's srcma
C0153562|T191|PT|176.2|ICD9CM|Kaposi's sarcoma, palate|Kaposi's sarcoma, palate
C0153562|T191|AB|176.2|ICD9CM|Palate - kpsi's sarcoma|Palate - kpsi's sarcoma
C0153563|T191|AB|176.3|ICD9CM|GI sites - kpsi's srcoma|GI sites - kpsi's srcoma
C0153563|T191|PT|176.3|ICD9CM|Kaposi's sarcoma, gastrointestinal sites|Kaposi's sarcoma, gastrointestinal sites
C0153564|T191|PT|176.4|ICD9CM|Kaposi's sarcoma, lung|Kaposi's sarcoma, lung
C0153564|T191|AB|176.4|ICD9CM|Lung - kaposi's sarcoma|Lung - kaposi's sarcoma
C0153565|T191|PT|176.5|ICD9CM|Kaposi's sarcoma, lymph nodes|Kaposi's sarcoma, lymph nodes
C0153565|T191|AB|176.5|ICD9CM|Lym nds - kpsi's sarcoma|Lym nds - kpsi's sarcoma
C0153566|T191|PT|176.8|ICD9CM|Kaposi's sarcoma, other specified sites|Kaposi's sarcoma, other specified sites
C0153566|T191|AB|176.8|ICD9CM|Spf sts - kpsi's sarcoma|Spf sts - kpsi's sarcoma
C0036220|T191|AB|176.9|ICD9CM|Kaposi's sarcoma NOS|Kaposi's sarcoma NOS
C0036220|T191|PT|176.9|ICD9CM|Kaposi's sarcoma, unspecified site|Kaposi's sarcoma, unspecified site
C0153567|T191|AB|179|ICD9CM|Malig neopl uterus NOS|Malig neopl uterus NOS
C0153567|T191|PT|179|ICD9CM|Malignant neoplasm of uterus, part unspecified|Malignant neoplasm of uterus, part unspecified
C0178251|T191|HT|179-189.99|ICD9CM|MALIGNANT NEOPLASM OF GENITOURINARY ORGANS|MALIGNANT NEOPLASM OF GENITOURINARY ORGANS
C0007847|T191|HT|180|ICD9CM|Malignant neoplasm of cervix uteri|Malignant neoplasm of cervix uteri
C0153569|T191|AB|180.0|ICD9CM|Malig neo endocervix|Malig neo endocervix
C0153569|T191|PT|180.0|ICD9CM|Malignant neoplasm of endocervix|Malignant neoplasm of endocervix
C0153570|T191|AB|180.1|ICD9CM|Malig neo exocervix|Malig neo exocervix
C0153570|T191|PT|180.1|ICD9CM|Malignant neoplasm of exocervix|Malignant neoplasm of exocervix
C0153571|T191|AB|180.8|ICD9CM|Malig neo cervix NEC|Malig neo cervix NEC
C0153571|T191|PT|180.8|ICD9CM|Malignant neoplasm of other specified sites of cervix|Malignant neoplasm of other specified sites of cervix
C0007847|T191|AB|180.9|ICD9CM|Mal neo cervix uteri NOS|Mal neo cervix uteri NOS
C0007847|T191|PT|180.9|ICD9CM|Malignant neoplasm of cervix uteri, unspecified site|Malignant neoplasm of cervix uteri, unspecified site
C0153572|T191|AB|181|ICD9CM|Malignant neopl placenta|Malignant neopl placenta
C0153572|T191|PT|181|ICD9CM|Malignant neoplasm of placenta|Malignant neoplasm of placenta
C0153574|T191|HT|182|ICD9CM|Malignant neoplasm of body of uterus|Malignant neoplasm of body of uterus
C1279258|T191|AB|182.0|ICD9CM|Malig neo corpus uteri|Malig neo corpus uteri
C1279258|T191|PT|182.0|ICD9CM|Malignant neoplasm of corpus uteri, except isthmus|Malignant neoplasm of corpus uteri, except isthmus
C0153575|T191|AB|182.1|ICD9CM|Mal neo uterine isthmus|Mal neo uterine isthmus
C0153575|T191|PT|182.1|ICD9CM|Malignant neoplasm of isthmus|Malignant neoplasm of isthmus
C0153576|T191|AB|182.8|ICD9CM|Mal neo body uterus NEC|Mal neo body uterus NEC
C0153576|T191|PT|182.8|ICD9CM|Malignant neoplasm of other specified sites of body of uterus|Malignant neoplasm of other specified sites of body of uterus
C0153577|T191|HT|183|ICD9CM|Malignant neoplasm of ovary and other uterine adnexa|Malignant neoplasm of ovary and other uterine adnexa
C1140680|T191|AB|183.0|ICD9CM|Malign neopl ovary|Malign neopl ovary
C1140680|T191|PT|183.0|ICD9CM|Malignant neoplasm of ovary|Malignant neoplasm of ovary
C0153579|T191|AB|183.2|ICD9CM|Mal neo fallopian tube|Mal neo fallopian tube
C0153579|T191|PT|183.2|ICD9CM|Malignant neoplasm of fallopian tube|Malignant neoplasm of fallopian tube
C0346866|T191|AB|183.3|ICD9CM|Mal neo broad ligament|Mal neo broad ligament
C0346866|T191|PT|183.3|ICD9CM|Malignant neoplasm of broad ligament of uterus|Malignant neoplasm of broad ligament of uterus
C0153581|T191|AB|183.4|ICD9CM|Malig neo parametrium|Malig neo parametrium
C0153581|T191|PT|183.4|ICD9CM|Malignant neoplasm of parametrium|Malignant neoplasm of parametrium
C0346867|T191|AB|183.5|ICD9CM|Mal neo round ligament|Mal neo round ligament
C0346867|T191|PT|183.5|ICD9CM|Malignant neoplasm of round ligament of uterus|Malignant neoplasm of round ligament of uterus
C0153583|T191|AB|183.8|ICD9CM|Mal neo adnexa NEC|Mal neo adnexa NEC
C0153583|T191|PT|183.8|ICD9CM|Malignant neoplasm of other specified sites of uterine adnexa|Malignant neoplasm of other specified sites of uterine adnexa
C0153584|T191|AB|183.9|ICD9CM|Mal neo adnexa NOS|Mal neo adnexa NOS
C0153584|T191|PT|183.9|ICD9CM|Malignant neoplasm of uterine adnexa, unspecified site|Malignant neoplasm of uterine adnexa, unspecified site
C0153585|T191|HT|184|ICD9CM|Malignant neoplasm of other and unspecified female genital organs|Malignant neoplasm of other and unspecified female genital organs
C0042237|T191|AB|184.0|ICD9CM|Malign neopl vagina|Malign neopl vagina
C0042237|T191|PT|184.0|ICD9CM|Malignant neoplasm of vagina|Malignant neoplasm of vagina
C0496814|T191|AB|184.1|ICD9CM|Mal neo labia majora|Mal neo labia majora
C0496814|T191|PT|184.1|ICD9CM|Malignant neoplasm of labia majora|Malignant neoplasm of labia majora
C0496815|T191|AB|184.2|ICD9CM|Mal neo labia minora|Mal neo labia minora
C0496815|T191|PT|184.2|ICD9CM|Malignant neoplasm of labia minora|Malignant neoplasm of labia minora
C0153589|T191|AB|184.3|ICD9CM|Malign neopl clitoris|Malign neopl clitoris
C0153589|T191|PT|184.3|ICD9CM|Malignant neoplasm of clitoris|Malignant neoplasm of clitoris
C0375071|T191|AB|184.4|ICD9CM|Malign neopl vulva NOS|Malign neopl vulva NOS
C0375071|T191|PT|184.4|ICD9CM|Malignant neoplasm of vulva, unspecified site|Malignant neoplasm of vulva, unspecified site
C0153591|T191|AB|184.8|ICD9CM|Mal neo female genit NEC|Mal neo female genit NEC
C0153591|T191|PT|184.8|ICD9CM|Malignant neoplasm of other specified sites of female genital organs|Malignant neoplasm of other specified sites of female genital organs
C0153592|T191|AB|184.9|ICD9CM|Mal neo female genit NOS|Mal neo female genit NOS
C0153592|T191|PT|184.9|ICD9CM|Malignant neoplasm of female genital organ, site unspecified|Malignant neoplasm of female genital organ, site unspecified
C0376358|T191|AB|185|ICD9CM|Malign neopl prostate|Malign neopl prostate
C0376358|T191|PT|185|ICD9CM|Malignant neoplasm of prostate|Malignant neoplasm of prostate
C0153594|T191|HT|186|ICD9CM|Malignant neoplasm of testis|Malignant neoplasm of testis
C0153595|T191|AB|186.0|ICD9CM|Mal neo undescend testis|Mal neo undescend testis
C0153595|T191|PT|186.0|ICD9CM|Malignant neoplasm of undescended testis|Malignant neoplasm of undescended testis
C0153596|T191|AB|186.9|ICD9CM|Malig neo testis NEC|Malig neo testis NEC
C0153596|T191|PT|186.9|ICD9CM|Malignant neoplasm of other and unspecified testis|Malignant neoplasm of other and unspecified testis
C0153597|T191|HT|187|ICD9CM|Malignant neoplasm of penis and other male genital organs|Malignant neoplasm of penis and other male genital organs
C0153598|T191|AB|187.1|ICD9CM|Malign neopl prepuce|Malign neopl prepuce
C0153598|T191|PT|187.1|ICD9CM|Malignant neoplasm of prepuce|Malignant neoplasm of prepuce
C0153599|T191|AB|187.2|ICD9CM|Malig neo glans penis|Malig neo glans penis
C0153599|T191|PT|187.2|ICD9CM|Malignant neoplasm of glans penis|Malignant neoplasm of glans penis
C0153600|T191|AB|187.3|ICD9CM|Malig neo penis body|Malig neo penis body
C0153600|T191|PT|187.3|ICD9CM|Malignant neoplasm of body of penis|Malignant neoplasm of body of penis
C0153601|T191|AB|187.4|ICD9CM|Malig neo penis NOS|Malig neo penis NOS
C0153601|T191|PT|187.4|ICD9CM|Malignant neoplasm of penis, part unspecified|Malignant neoplasm of penis, part unspecified
C0153602|T191|AB|187.5|ICD9CM|Malig neo epididymis|Malig neo epididymis
C0153602|T191|PT|187.5|ICD9CM|Malignant neoplasm of epididymis|Malignant neoplasm of epididymis
C0153603|T191|AB|187.6|ICD9CM|Mal neo spermatic cord|Mal neo spermatic cord
C0153603|T191|PT|187.6|ICD9CM|Malignant neoplasm of spermatic cord|Malignant neoplasm of spermatic cord
C0153604|T191|AB|187.7|ICD9CM|Malign neopl scrotum|Malign neopl scrotum
C0153604|T191|PT|187.7|ICD9CM|Malignant neoplasm of scrotum|Malignant neoplasm of scrotum
C0153605|T191|AB|187.8|ICD9CM|Mal neo male genital NEC|Mal neo male genital NEC
C0153605|T191|PT|187.8|ICD9CM|Malignant neoplasm of other specified sites of male genital organs|Malignant neoplasm of other specified sites of male genital organs
C0153606|T191|AB|187.9|ICD9CM|Mal neo male genital NOS|Mal neo male genital NOS
C0153606|T191|PT|187.9|ICD9CM|Malignant neoplasm of male genital organ, site unspecified|Malignant neoplasm of male genital organ, site unspecified
C0005684|T191|HT|188|ICD9CM|Malignant neoplasm of bladder|Malignant neoplasm of bladder
C0496826|T191|AB|188.0|ICD9CM|Mal neo bladder-trigone|Mal neo bladder-trigone
C0496826|T191|PT|188.0|ICD9CM|Malignant neoplasm of trigone of urinary bladder|Malignant neoplasm of trigone of urinary bladder
C0496827|T191|AB|188.1|ICD9CM|Mal neo bladder-dome|Mal neo bladder-dome
C0496827|T191|PT|188.1|ICD9CM|Malignant neoplasm of dome of urinary bladder|Malignant neoplasm of dome of urinary bladder
C0496828|T191|AB|188.2|ICD9CM|Mal neo bladder-lateral|Mal neo bladder-lateral
C0496828|T191|PT|188.2|ICD9CM|Malignant neoplasm of lateral wall of urinary bladder|Malignant neoplasm of lateral wall of urinary bladder
C0153611|T191|AB|188.3|ICD9CM|Mal neo bladder-anterior|Mal neo bladder-anterior
C0153611|T191|PT|188.3|ICD9CM|Malignant neoplasm of anterior wall of urinary bladder|Malignant neoplasm of anterior wall of urinary bladder
C0153612|T191|AB|188.4|ICD9CM|Mal neo bladder-post|Mal neo bladder-post
C0153612|T191|PT|188.4|ICD9CM|Malignant neoplasm of posterior wall of urinary bladder|Malignant neoplasm of posterior wall of urinary bladder
C0153613|T191|AB|188.5|ICD9CM|Mal neo bladder neck|Mal neo bladder neck
C0153613|T191|PT|188.5|ICD9CM|Malignant neoplasm of bladder neck|Malignant neoplasm of bladder neck
C0153614|T191|AB|188.6|ICD9CM|Mal neo ureteric orifice|Mal neo ureteric orifice
C0153614|T191|PT|188.6|ICD9CM|Malignant neoplasm of ureteric orifice|Malignant neoplasm of ureteric orifice
C0153615|T191|AB|188.7|ICD9CM|Malig neo urachus|Malig neo urachus
C0153615|T191|PT|188.7|ICD9CM|Malignant neoplasm of urachus|Malignant neoplasm of urachus
C0153616|T191|AB|188.8|ICD9CM|Malig neo bladder NEC|Malig neo bladder NEC
C0153616|T191|PT|188.8|ICD9CM|Malignant neoplasm of other specified sites of bladder|Malignant neoplasm of other specified sites of bladder
C0005684|T191|AB|188.9|ICD9CM|Malig neo bladder NOS|Malig neo bladder NOS
C0005684|T191|PT|188.9|ICD9CM|Malignant neoplasm of bladder, part unspecified|Malignant neoplasm of bladder, part unspecified
C0153617|T191|HT|189|ICD9CM|Malignant neoplasm of kidney and other and unspecified urinary organs|Malignant neoplasm of kidney and other and unspecified urinary organs
C0494158|T191|AB|189.0|ICD9CM|Malig neopl kidney|Malig neopl kidney
C0494158|T191|PT|189.0|ICD9CM|Malignant neoplasm of kidney, except pelvis|Malignant neoplasm of kidney, except pelvis
C0153618|T191|AB|189.1|ICD9CM|Malig neo renal pelvis|Malig neo renal pelvis
C0153618|T191|PT|189.1|ICD9CM|Malignant neoplasm of renal pelvis|Malignant neoplasm of renal pelvis
C0153619|T191|AB|189.2|ICD9CM|Malign neopl ureter|Malign neopl ureter
C0153619|T191|PT|189.2|ICD9CM|Malignant neoplasm of ureter|Malignant neoplasm of ureter
C0153620|T191|AB|189.3|ICD9CM|Malign neopl urethra|Malign neopl urethra
C0153620|T191|PT|189.3|ICD9CM|Malignant neoplasm of urethra|Malignant neoplasm of urethra
C0153621|T191|AB|189.4|ICD9CM|Mal neo paraurethral|Mal neo paraurethral
C0153621|T191|PT|189.4|ICD9CM|Malignant neoplasm of paraurethral glands|Malignant neoplasm of paraurethral glands
C0153622|T191|AB|189.8|ICD9CM|Mal neo urinary NEC|Mal neo urinary NEC
C0153622|T191|PT|189.8|ICD9CM|Malignant neoplasm of other specified sites of urinary organs|Malignant neoplasm of other specified sites of urinary organs
C0348371|T191|AB|189.9|ICD9CM|Mal neo urinary NOS|Mal neo urinary NOS
C0348371|T191|PT|189.9|ICD9CM|Malignant neoplasm of urinary organ, site unspecified|Malignant neoplasm of urinary organ, site unspecified
C0496836|T191|HT|190|ICD9CM|Malignant neoplasm of eye|Malignant neoplasm of eye
C0347071|T191|HT|190-199.99|ICD9CM|MALIGNANT NEOPLASM OF OTHER AND UNSPECIFIED SITES|MALIGNANT NEOPLASM OF OTHER AND UNSPECIFIED SITES
C0153625|T191|AB|190.0|ICD9CM|Malign neopl eyeball|Malign neopl eyeball
C0153625|T191|PT|190.0|ICD9CM|Malignant neoplasm of eyeball, except conjunctiva, cornea, retina, and choroid|Malignant neoplasm of eyeball, except conjunctiva, cornea, retina, and choroid
C0153626|T191|AB|190.1|ICD9CM|Malign neopl orbit|Malign neopl orbit
C0153626|T191|PT|190.1|ICD9CM|Malignant neoplasm of orbit|Malignant neoplasm of orbit
C0153627|T191|AB|190.2|ICD9CM|Mal neo lacrimal gland|Mal neo lacrimal gland
C0153627|T191|PT|190.2|ICD9CM|Malignant neoplasm of lacrimal gland|Malignant neoplasm of lacrimal gland
C0153628|T191|AB|190.3|ICD9CM|Mal neo conjunctiva|Mal neo conjunctiva
C0153628|T191|PT|190.3|ICD9CM|Malignant neoplasm of conjunctiva|Malignant neoplasm of conjunctiva
C0153629|T191|AB|190.4|ICD9CM|Malign neopl cornea|Malign neopl cornea
C0153629|T191|PT|190.4|ICD9CM|Malignant neoplasm of cornea|Malignant neoplasm of cornea
C0024622|T191|AB|190.5|ICD9CM|Malign neopl retina|Malign neopl retina
C0024622|T191|PT|190.5|ICD9CM|Malignant neoplasm of retina|Malignant neoplasm of retina
C0153630|T191|AB|190.6|ICD9CM|Malign neopl choroid|Malign neopl choroid
C0153630|T191|PT|190.6|ICD9CM|Malignant neoplasm of choroid|Malignant neoplasm of choroid
C0153631|T191|AB|190.7|ICD9CM|Mal neo lacrimal duct|Mal neo lacrimal duct
C0153631|T191|PT|190.7|ICD9CM|Malignant neoplasm of lacrimal duct|Malignant neoplasm of lacrimal duct
C0153632|T191|AB|190.8|ICD9CM|Malign neopl eye NEC|Malign neopl eye NEC
C0153632|T191|PT|190.8|ICD9CM|Malignant neoplasm of other specified sites of eye|Malignant neoplasm of other specified sites of eye
C0496836|T191|AB|190.9|ICD9CM|Malign neopl eye NOS|Malign neopl eye NOS
C0496836|T191|PT|190.9|ICD9CM|Malignant neoplasm of eye, part unspecified|Malignant neoplasm of eye, part unspecified
C0153633|T191|HT|191|ICD9CM|Malignant neoplasm of brain|Malignant neoplasm of brain
C0153634|T191|AB|191.0|ICD9CM|Malign neopl cerebrum|Malign neopl cerebrum
C0153634|T191|PT|191.0|ICD9CM|Malignant neoplasm of cerebrum, except lobes and ventricles|Malignant neoplasm of cerebrum, except lobes and ventricles
C0153635|T191|AB|191.1|ICD9CM|Malig neo frontal lobe|Malig neo frontal lobe
C0153635|T191|PT|191.1|ICD9CM|Malignant neoplasm of frontal lobe|Malignant neoplasm of frontal lobe
C0153636|T191|AB|191.2|ICD9CM|Mal neo temporal lobe|Mal neo temporal lobe
C0153636|T191|PT|191.2|ICD9CM|Malignant neoplasm of temporal lobe|Malignant neoplasm of temporal lobe
C0153637|T191|AB|191.3|ICD9CM|Mal neo parietal lobe|Mal neo parietal lobe
C0153637|T191|PT|191.3|ICD9CM|Malignant neoplasm of parietal lobe|Malignant neoplasm of parietal lobe
C0153638|T191|AB|191.4|ICD9CM|Mal neo occipital lobe|Mal neo occipital lobe
C0153638|T191|PT|191.4|ICD9CM|Malignant neoplasm of occipital lobe|Malignant neoplasm of occipital lobe
C0346906|T191|AB|191.5|ICD9CM|Mal neo cereb ventricle|Mal neo cereb ventricle
C0346906|T191|PT|191.5|ICD9CM|Malignant neoplasm of ventricles|Malignant neoplasm of ventricles
C0153640|T191|AB|191.6|ICD9CM|Mal neo cerebellum NOS|Mal neo cerebellum NOS
C0153640|T191|PT|191.6|ICD9CM|Malignant neoplasm of cerebellum nos|Malignant neoplasm of cerebellum nos
C0153641|T191|AB|191.7|ICD9CM|Mal neo brain stem|Mal neo brain stem
C0153641|T191|PT|191.7|ICD9CM|Malignant neoplasm of brain stem|Malignant neoplasm of brain stem
C0153642|T191|AB|191.8|ICD9CM|Malig neo brain NEC|Malig neo brain NEC
C0153642|T191|PT|191.8|ICD9CM|Malignant neoplasm of other parts of brain|Malignant neoplasm of other parts of brain
C0153633|T191|AB|191.9|ICD9CM|Malig neo brain NOS|Malig neo brain NOS
C0153633|T191|PT|191.9|ICD9CM|Malignant neoplasm of brain, unspecified|Malignant neoplasm of brain, unspecified
C0153643|T191|HT|192|ICD9CM|Malignant neoplasm of other and unspecified parts of nervous system|Malignant neoplasm of other and unspecified parts of nervous system
C0153644|T191|AB|192.0|ICD9CM|Mal neo cranial nerves|Mal neo cranial nerves
C0153644|T191|PT|192.0|ICD9CM|Malignant neoplasm of cranial nerves|Malignant neoplasm of cranial nerves
C0153645|T191|AB|192.1|ICD9CM|Mal neo cerebral mening|Mal neo cerebral mening
C0153645|T191|PT|192.1|ICD9CM|Malignant neoplasm of cerebral meninges|Malignant neoplasm of cerebral meninges
C0153646|T191|AB|192.2|ICD9CM|Mal neo spinal cord|Mal neo spinal cord
C0153646|T191|PT|192.2|ICD9CM|Malignant neoplasm of spinal cord|Malignant neoplasm of spinal cord
C0153647|T191|AB|192.3|ICD9CM|Mal neo spinal meninges|Mal neo spinal meninges
C0153647|T191|PT|192.3|ICD9CM|Malignant neoplasm of spinal meninges|Malignant neoplasm of spinal meninges
C0153648|T191|AB|192.8|ICD9CM|Mal neo nervous syst NEC|Mal neo nervous syst NEC
C0153648|T191|PT|192.8|ICD9CM|Malignant neoplasm of other specified sites of nervous system|Malignant neoplasm of other specified sites of nervous system
C0153643|T191|AB|192.9|ICD9CM|Mal neo nervous syst NOS|Mal neo nervous syst NOS
C0153643|T191|PT|192.9|ICD9CM|Malignant neoplasm of nervous system, part unspecified|Malignant neoplasm of nervous system, part unspecified
C0007115|T191|AB|193|ICD9CM|Malign neopl thyroid|Malign neopl thyroid
C0007115|T191|PT|193|ICD9CM|Malignant neoplasm of thyroid gland|Malignant neoplasm of thyroid gland
C0153651|T191|HT|194|ICD9CM|Malignant neoplasm of other endocrine glands and related structures|Malignant neoplasm of other endocrine glands and related structures
C0750887|T191|AB|194.0|ICD9CM|Malign neopl adrenal|Malign neopl adrenal
C0750887|T191|PT|194.0|ICD9CM|Malignant neoplasm of adrenal gland|Malignant neoplasm of adrenal gland
C0153653|T191|AB|194.1|ICD9CM|Malig neo parathyroid|Malig neo parathyroid
C0153653|T191|PT|194.1|ICD9CM|Malignant neoplasm of parathyroid gland|Malignant neoplasm of parathyroid gland
C0153654|T191|AB|194.3|ICD9CM|Malig neo pituitary|Malig neo pituitary
C0153654|T191|PT|194.3|ICD9CM|Malignant neoplasm of pituitary gland and craniopharyngeal duct|Malignant neoplasm of pituitary gland and craniopharyngeal duct
C0153655|T191|AB|194.4|ICD9CM|Malign neo pineal gland|Malign neo pineal gland
C0153655|T191|PT|194.4|ICD9CM|Malignant neoplasm of pineal gland|Malignant neoplasm of pineal gland
C0153656|T191|AB|194.5|ICD9CM|Mal neo carotid body|Mal neo carotid body
C0153656|T191|PT|194.5|ICD9CM|Malignant neoplasm of carotid body|Malignant neoplasm of carotid body
C0438413|T191|AB|194.6|ICD9CM|Mal neo paraganglia NEC|Mal neo paraganglia NEC
C0438413|T191|PT|194.6|ICD9CM|Malignant neoplasm of aortic body and other paraganglia|Malignant neoplasm of aortic body and other paraganglia
C0153651|T191|AB|194.8|ICD9CM|Mal neo endocrine NEC|Mal neo endocrine NEC
C0153651|T191|PT|194.8|ICD9CM|Malignant neoplasm of other endocrine glands and related structures|Malignant neoplasm of other endocrine glands and related structures
C0153658|T191|AB|194.9|ICD9CM|Mal neo endocrine NOS|Mal neo endocrine NOS
C0153658|T191|PT|194.9|ICD9CM|Malignant neoplasm of endocrine gland, site unspecified|Malignant neoplasm of endocrine gland, site unspecified
C0153659|T191|HT|195|ICD9CM|Malignant neoplasm of other and ill-defined sites|Malignant neoplasm of other and ill-defined sites
C0153660|T191|AB|195.0|ICD9CM|Mal neo head/face/neck|Mal neo head/face/neck
C0153660|T191|PT|195.0|ICD9CM|Malignant neoplasm of head, face, and neck|Malignant neoplasm of head, face, and neck
C0153661|T191|AB|195.1|ICD9CM|Malign neopl thorax|Malign neopl thorax
C0153661|T191|PT|195.1|ICD9CM|Malignant neoplasm of thorax|Malignant neoplasm of thorax
C0153662|T191|AB|195.2|ICD9CM|Malig neo abdomen|Malig neo abdomen
C0153662|T191|PT|195.2|ICD9CM|Malignant neoplasm of abdomen|Malignant neoplasm of abdomen
C0153663|T191|AB|195.3|ICD9CM|Malign neopl pelvis|Malign neopl pelvis
C0153663|T191|PT|195.3|ICD9CM|Malignant neoplasm of pelvis|Malignant neoplasm of pelvis
C0153664|T191|AB|195.4|ICD9CM|Malign neopl arm|Malign neopl arm
C0153664|T191|PT|195.4|ICD9CM|Malignant neoplasm of upper limb|Malignant neoplasm of upper limb
C0153665|T191|AB|195.5|ICD9CM|Malign neopl leg|Malign neopl leg
C0153665|T191|PT|195.5|ICD9CM|Malignant neoplasm of lower limb|Malignant neoplasm of lower limb
C0153666|T191|AB|195.8|ICD9CM|Malig neo site NEC|Malig neo site NEC
C0153666|T191|PT|195.8|ICD9CM|Malignant neoplasm of other specified sites|Malignant neoplasm of other specified sites
C0686619|T191|HT|196|ICD9CM|Secondary and unspecified malignant neoplasm of lymph nodes|Secondary and unspecified malignant neoplasm of lymph nodes
C0153668|T191|AB|196.0|ICD9CM|Mal neo lymph-head/neck|Mal neo lymph-head/neck
C0153668|T191|PT|196.0|ICD9CM|Secondary and unspecified malignant neoplasm of lymph nodes of head, face, and neck|Secondary and unspecified malignant neoplasm of lymph nodes of head, face, and neck
C0686645|T191|AB|196.1|ICD9CM|Mal neo lymph-intrathor|Mal neo lymph-intrathor
C0686645|T191|PT|196.1|ICD9CM|Secondary and unspecified malignant neoplasm of intrathoracic lymph nodes|Secondary and unspecified malignant neoplasm of intrathoracic lymph nodes
C0686655|T191|AB|196.2|ICD9CM|Mal neo lymph intra-abd|Mal neo lymph intra-abd
C0686655|T191|PT|196.2|ICD9CM|Secondary and unspecified malignant neoplasm of intra-abdominal lymph nodes|Secondary and unspecified malignant neoplasm of intra-abdominal lymph nodes
C0153671|T191|AB|196.3|ICD9CM|Mal neo lymph-axilla/arm|Mal neo lymph-axilla/arm
C0153671|T191|PT|196.3|ICD9CM|Secondary and unspecified malignant neoplasm of lymph nodes of axilla and upper limb|Secondary and unspecified malignant neoplasm of lymph nodes of axilla and upper limb
C0347055|T191|AB|196.5|ICD9CM|Mal neo lymph-inguin/leg|Mal neo lymph-inguin/leg
C0347055|T191|PT|196.5|ICD9CM|Secondary and unspecified malignant neoplasm of lymph nodes of inguinal region and lower limb|Secondary and unspecified malignant neoplasm of lymph nodes of inguinal region and lower limb
C0686689|T191|AB|196.6|ICD9CM|Mal neo lymph-intrapelv|Mal neo lymph-intrapelv
C0686689|T191|PT|196.6|ICD9CM|Secondary and unspecified malignant neoplasm of intrapelvic lymph nodes|Secondary and unspecified malignant neoplasm of intrapelvic lymph nodes
C0348382|T191|AB|196.8|ICD9CM|Mal neo lymph node-mult|Mal neo lymph node-mult
C0348382|T191|PT|196.8|ICD9CM|Secondary and unspecified malignant neoplasm of lymph nodes of multiple sites|Secondary and unspecified malignant neoplasm of lymph nodes of multiple sites
C0686619|T191|AB|196.9|ICD9CM|Mal neo lymph node NOS|Mal neo lymph node NOS
C0686619|T191|PT|196.9|ICD9CM|Secondary and unspecified malignant neoplasm of lymph nodes, site unspecified|Secondary and unspecified malignant neoplasm of lymph nodes, site unspecified
C0153675|T191|HT|197|ICD9CM|Secondary malignant neoplasm of respiratory and digestive systems|Secondary malignant neoplasm of respiratory and digestive systems
C0153676|T191|AB|197.0|ICD9CM|Secondary malig neo lung|Secondary malig neo lung
C0153676|T191|PT|197.0|ICD9CM|Secondary malignant neoplasm of lung|Secondary malignant neoplasm of lung
C0153677|T191|AB|197.1|ICD9CM|Sec mal neo mediastinum|Sec mal neo mediastinum
C0153677|T191|PT|197.1|ICD9CM|Secondary malignant neoplasm of mediastinum|Secondary malignant neoplasm of mediastinum
C0153678|T191|AB|197.2|ICD9CM|Second malig neo pleura|Second malig neo pleura
C0153678|T191|PT|197.2|ICD9CM|Secondary malignant neoplasm of pleura|Secondary malignant neoplasm of pleura
C2745961|T191|AB|197.3|ICD9CM|Sec malig neo resp NEC|Sec malig neo resp NEC
C2745961|T191|PT|197.3|ICD9CM|Secondary malignant neoplasm of other respiratory organs|Secondary malignant neoplasm of other respiratory organs
C0494164|T191|AB|197.4|ICD9CM|Sec malig neo sm bowel|Sec malig neo sm bowel
C0494164|T191|PT|197.4|ICD9CM|Secondary malignant neoplasm of small intestine including duodenum|Secondary malignant neoplasm of small intestine including duodenum
C0153681|T191|AB|197.5|ICD9CM|Sec malig neo lg bowel|Sec malig neo lg bowel
C0153681|T191|PT|197.5|ICD9CM|Secondary malignant neoplasm of large intestine and rectum|Secondary malignant neoplasm of large intestine and rectum
C0036528|T191|AB|197.6|ICD9CM|Sec mal neo peritoneum|Sec mal neo peritoneum
C0036528|T191|PT|197.6|ICD9CM|Secondary malignant neoplasm of retroperitoneum and peritoneum|Secondary malignant neoplasm of retroperitoneum and peritoneum
C0494165|T191|PT|197.7|ICD9CM|Malignant neoplasm of liver, secondary|Malignant neoplasm of liver, secondary
C0494165|T191|AB|197.7|ICD9CM|Second malig neo liver|Second malig neo liver
C0153683|T191|AB|197.8|ICD9CM|Sec mal neo GI NEC|Sec mal neo GI NEC
C0153683|T191|PT|197.8|ICD9CM|Secondary malignant neoplasm of other digestive organs and spleen|Secondary malignant neoplasm of other digestive organs and spleen
C0153684|T191|HT|198|ICD9CM|Secondary malignant neoplasm of other specified sites|Secondary malignant neoplasm of other specified sites
C0153685|T191|AB|198.0|ICD9CM|Second malig neo kidney|Second malig neo kidney
C0153685|T191|PT|198.0|ICD9CM|Secondary malignant neoplasm of kidney|Secondary malignant neoplasm of kidney
C2845968|T191|AB|198.1|ICD9CM|Sec malig neo urin NEC|Sec malig neo urin NEC
C2845968|T191|PT|198.1|ICD9CM|Secondary malignant neoplasm of other urinary organs|Secondary malignant neoplasm of other urinary organs
C0153687|T191|AB|198.2|ICD9CM|Secondary malig neo skin|Secondary malig neo skin
C0153687|T191|PT|198.2|ICD9CM|Secondary malignant neoplasm of skin|Secondary malignant neoplasm of skin
C0153688|T191|AB|198.3|ICD9CM|Sec mal neo brain/spine|Sec mal neo brain/spine
C0153688|T191|PT|198.3|ICD9CM|Secondary malignant neoplasm of brain and spinal cord|Secondary malignant neoplasm of brain and spinal cord
C0153689|T191|AB|198.4|ICD9CM|Sec malig neo nerve NEC|Sec malig neo nerve NEC
C0153689|T191|PT|198.4|ICD9CM|Secondary malignant neoplasm of other parts of nervous system|Secondary malignant neoplasm of other parts of nervous system
C0153690|T191|AB|198.5|ICD9CM|Secondary malig neo bone|Secondary malig neo bone
C0153690|T191|PT|198.5|ICD9CM|Secondary malignant neoplasm of bone and bone marrow|Secondary malignant neoplasm of bone and bone marrow
C3647143|T191|AB|198.6|ICD9CM|Second malig neo ovary|Second malig neo ovary
C3647143|T191|PT|198.6|ICD9CM|Secondary malignant neoplasm of ovary|Secondary malignant neoplasm of ovary
C0153691|T191|AB|198.7|ICD9CM|Second malig neo adrenal|Second malig neo adrenal
C0153691|T191|PT|198.7|ICD9CM|Secondary malignant neoplasm of adrenal gland|Secondary malignant neoplasm of adrenal gland
C0153684|T191|HT|198.8|ICD9CM|Secondary malignant neoplasm of other specified sites|Secondary malignant neoplasm of other specified sites
C0346993|T191|AB|198.81|ICD9CM|Second malig neo breast|Second malig neo breast
C0346993|T191|PT|198.81|ICD9CM|Secondary malignant neoplasm of breast|Secondary malignant neoplasm of breast
C0153693|T191|AB|198.82|ICD9CM|Second malig neo genital|Second malig neo genital
C0153693|T191|PT|198.82|ICD9CM|Secondary malignant neoplasm of genital organs|Secondary malignant neoplasm of genital organs
C0153684|T191|AB|198.89|ICD9CM|Secondary malig neo NEC|Secondary malig neo NEC
C0153684|T191|PT|198.89|ICD9CM|Secondary malignant neoplasm of other specified sites|Secondary malignant neoplasm of other specified sites
C0006826|T191|HT|199|ICD9CM|Malignant neoplasm without specification of site|Malignant neoplasm without specification of site
C0346957|T191|PT|199.0|ICD9CM|Disseminated malignant neoplasm without specification of site|Disseminated malignant neoplasm without specification of site
C0346957|T191|AB|199.0|ICD9CM|Malig neo disseminated|Malig neo disseminated
C0347071|T191|AB|199.1|ICD9CM|Malignant neoplasm NOS|Malignant neoplasm NOS
C0347071|T191|PT|199.1|ICD9CM|Other malignant neoplasm without specification of site|Other malignant neoplasm without specification of site
C2349259|T191|AB|199.2|ICD9CM|Malig neopl-transp organ|Malig neopl-transp organ
C2349259|T191|PT|199.2|ICD9CM|Malignant neoplasm associated with transplant organ|Malignant neoplasm associated with transplant organ
C1955727|T191|HT|200|ICD9CM|Lymphosarcoma and reticulosarcoma and other specified malignant tumors of lymphatic tissue|Lymphosarcoma and reticulosarcoma and other specified malignant tumors of lymphatic tissue
C0348393|T191|HT|200-208.99|ICD9CM|MALIGNANT NEOPLASM OF LYMPHATIC AND HEMATOPOIETIC TISSUE|MALIGNANT NEOPLASM OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0024302|T191|HT|200.0|ICD9CM|Reticulosarcoma|Reticulosarcoma
C0375075|T191|AB|200.00|ICD9CM|Retclsrc unsp xtrndl org|Retclsrc unsp xtrndl org
C0375075|T191|PT|200.00|ICD9CM|Reticulosarcoma, unspecified site, extranodal and solid organ sites|Reticulosarcoma, unspecified site, extranodal and solid organ sites
C0153696|T191|AB|200.01|ICD9CM|Reticulosarcoma head|Reticulosarcoma head
C0153696|T191|PT|200.01|ICD9CM|Reticulosarcoma, lymph nodes of head, face, and neck|Reticulosarcoma, lymph nodes of head, face, and neck
C0153697|T191|AB|200.02|ICD9CM|Reticulosarcoma thorax|Reticulosarcoma thorax
C0153697|T191|PT|200.02|ICD9CM|Reticulosarcoma, intrathoracic lymph nodes|Reticulosarcoma, intrathoracic lymph nodes
C0153698|T191|AB|200.03|ICD9CM|Reticulosarcoma abdom|Reticulosarcoma abdom
C0153698|T191|PT|200.03|ICD9CM|Reticulosarcoma, intra-abdominal lymph nodes|Reticulosarcoma, intra-abdominal lymph nodes
C0153699|T191|AB|200.04|ICD9CM|Reticulosarcoma axilla|Reticulosarcoma axilla
C0153699|T191|PT|200.04|ICD9CM|Reticulosarcoma, lymph nodes of axilla and upper limb|Reticulosarcoma, lymph nodes of axilla and upper limb
C0153700|T191|AB|200.05|ICD9CM|Reticulosarcoma inguin|Reticulosarcoma inguin
C0153700|T191|PT|200.05|ICD9CM|Reticulosarcoma, lymph nodes of inguinal region and lower limb|Reticulosarcoma, lymph nodes of inguinal region and lower limb
C0153701|T191|AB|200.06|ICD9CM|Reticulosarcoma pelvic|Reticulosarcoma pelvic
C0153701|T191|PT|200.06|ICD9CM|Reticulosarcoma, intrapelvic lymph nodes|Reticulosarcoma, intrapelvic lymph nodes
C0153702|T191|AB|200.07|ICD9CM|Reticulosarcoma spleen|Reticulosarcoma spleen
C0153702|T191|PT|200.07|ICD9CM|Reticulosarcoma, spleen|Reticulosarcoma, spleen
C0153703|T191|AB|200.08|ICD9CM|Reticulosarcoma mult|Reticulosarcoma mult
C0153703|T191|PT|200.08|ICD9CM|Reticulosarcoma, lymph nodes of multiple sites|Reticulosarcoma, lymph nodes of multiple sites
C3714542|T191|HT|200.1|ICD9CM|Lymphosarcoma|Lymphosarcoma
C0375076|T191|PT|200.10|ICD9CM|Lymphosarcoma, unspecified site, extranodal and solid organ sites|Lymphosarcoma, unspecified site, extranodal and solid organ sites
C0375076|T191|AB|200.10|ICD9CM|Lymphsrc unsp xtrndl org|Lymphsrc unsp xtrndl org
C0153704|T191|AB|200.11|ICD9CM|Lymphosarcoma head|Lymphosarcoma head
C0153704|T191|PT|200.11|ICD9CM|Lymphosarcoma, lymph nodes of head, face, and neck|Lymphosarcoma, lymph nodes of head, face, and neck
C0153705|T191|AB|200.12|ICD9CM|Lymphosarcoma thorax|Lymphosarcoma thorax
C0153705|T191|PT|200.12|ICD9CM|Lymphosarcoma, intrathoracic lymph nodes|Lymphosarcoma, intrathoracic lymph nodes
C0153706|T191|AB|200.13|ICD9CM|Lymphosarcoma abdom|Lymphosarcoma abdom
C0153706|T191|PT|200.13|ICD9CM|Lymphosarcoma, intra-abdominal lymph nodes|Lymphosarcoma, intra-abdominal lymph nodes
C0153707|T191|AB|200.14|ICD9CM|Lymphosarcoma axilla|Lymphosarcoma axilla
C0153707|T191|PT|200.14|ICD9CM|Lymphosarcoma, lymph nodes of axilla and upper limb|Lymphosarcoma, lymph nodes of axilla and upper limb
C0153708|T191|AB|200.15|ICD9CM|Lymphosarcoma inguin|Lymphosarcoma inguin
C0153708|T191|PT|200.15|ICD9CM|Lymphosarcoma, lymph nodes of inguinal region and lower limb|Lymphosarcoma, lymph nodes of inguinal region and lower limb
C0153709|T191|AB|200.16|ICD9CM|Lymphosarcoma pelvic|Lymphosarcoma pelvic
C0153709|T191|PT|200.16|ICD9CM|Lymphosarcoma, intrapelvic lymph nodes|Lymphosarcoma, intrapelvic lymph nodes
C0153710|T191|AB|200.17|ICD9CM|Lymphosarcoma spleen|Lymphosarcoma spleen
C0153710|T191|PT|200.17|ICD9CM|Lymphosarcoma, spleen|Lymphosarcoma, spleen
C0153711|T191|AB|200.18|ICD9CM|Lymphosarcoma mult|Lymphosarcoma mult
C0153711|T191|PT|200.18|ICD9CM|Lymphosarcoma, lymph nodes of multiple sites|Lymphosarcoma, lymph nodes of multiple sites
C0006413|T191|HT|200.2|ICD9CM|Burkitt's tumor or lymphoma|Burkitt's tumor or lymphoma
C0375077|T191|AB|200.20|ICD9CM|Brkt tmr unsp xtrndl org|Brkt tmr unsp xtrndl org
C0375077|T191|PT|200.20|ICD9CM|Burkitt's tumor or lymphoma, unspecified site, extranodal and solid organ sites|Burkitt's tumor or lymphoma, unspecified site, extranodal and solid organ sites
C0153712|T191|AB|200.21|ICD9CM|Burkitt's tumor head|Burkitt's tumor head
C0153712|T191|PT|200.21|ICD9CM|Burkitt's tumor or lymphoma, lymph nodes of head, face, and neck|Burkitt's tumor or lymphoma, lymph nodes of head, face, and neck
C0153713|T191|PT|200.22|ICD9CM|Burkitt's tumor or lymphoma, intrathoracic lymph nodes|Burkitt's tumor or lymphoma, intrathoracic lymph nodes
C0153713|T191|AB|200.22|ICD9CM|Burkitt's tumor thorax|Burkitt's tumor thorax
C0153714|T191|AB|200.23|ICD9CM|Burkitt's tumor abdom|Burkitt's tumor abdom
C0153714|T191|PT|200.23|ICD9CM|Burkitt's tumor or lymphoma, intra-abdominal lymph nodes|Burkitt's tumor or lymphoma, intra-abdominal lymph nodes
C0153715|T191|AB|200.24|ICD9CM|Burkitt's tumor axilla|Burkitt's tumor axilla
C0153715|T191|PT|200.24|ICD9CM|Burkitt's tumor or lymphoma, lymph nodes of axilla and upper limb|Burkitt's tumor or lymphoma, lymph nodes of axilla and upper limb
C0153716|T191|AB|200.25|ICD9CM|Burkitt's tumor inguin|Burkitt's tumor inguin
C0153716|T191|PT|200.25|ICD9CM|Burkitt's tumor or lymphoma, lymph nodes of inguinal region and lower limb|Burkitt's tumor or lymphoma, lymph nodes of inguinal region and lower limb
C0153717|T191|PT|200.26|ICD9CM|Burkitt's tumor or lymphoma, intrapelvic lymph nodes|Burkitt's tumor or lymphoma, intrapelvic lymph nodes
C0153717|T191|AB|200.26|ICD9CM|Burkitt's tumor pelvic|Burkitt's tumor pelvic
C0686546|T191|PT|200.27|ICD9CM|Burkitt's tumor or lymphoma, spleen|Burkitt's tumor or lymphoma, spleen
C0686546|T191|AB|200.27|ICD9CM|Burkitt's tumor spleen|Burkitt's tumor spleen
C0153719|T191|AB|200.28|ICD9CM|Burkitt's tumor mult|Burkitt's tumor mult
C0153719|T191|PT|200.28|ICD9CM|Burkitt's tumor or lymphoma, lymph nodes of multiple sites|Burkitt's tumor or lymphoma, lymph nodes of multiple sites
C1367654|T191|HT|200.3|ICD9CM|Marginal zone lymphoma|Marginal zone lymphoma
C1955681|T191|PT|200.30|ICD9CM|Marginal zone lymphoma, unspecified site, extranodal and solid organ sites|Marginal zone lymphoma, unspecified site, extranodal and solid organ sites
C1955681|T191|AB|200.30|ICD9CM|Margnl zone lym xtrndl|Margnl zone lym xtrndl
C1955682|T191|AB|200.31|ICD9CM|Margin zone lym head|Margin zone lym head
C1955682|T191|PT|200.31|ICD9CM|Marginal zone lymphoma, lymph nodes of head, face, and neck|Marginal zone lymphoma, lymph nodes of head, face, and neck
C1955683|T191|AB|200.32|ICD9CM|Margin zone lym thorax|Margin zone lym thorax
C1955683|T191|PT|200.32|ICD9CM|Marginal zone lymphoma, intrathoracic lymph nodes|Marginal zone lymphoma, intrathoracic lymph nodes
C1955684|T191|AB|200.33|ICD9CM|Margin zone lym abdom|Margin zone lym abdom
C1955684|T191|PT|200.33|ICD9CM|Marginal zone lymphoma, intraabdominal lymph nodes|Marginal zone lymphoma, intraabdominal lymph nodes
C1955685|T191|AB|200.34|ICD9CM|Margin zone lym axilla|Margin zone lym axilla
C1955685|T191|PT|200.34|ICD9CM|Marginal zone lymphoma, lymph nodes of axilla and upper limb|Marginal zone lymphoma, lymph nodes of axilla and upper limb
C1955686|T191|AB|200.35|ICD9CM|Margin zone lym inguin|Margin zone lym inguin
C1955686|T191|PT|200.35|ICD9CM|Marginal zone lymphoma, lymph nodes of inguinal region and lower limb|Marginal zone lymphoma, lymph nodes of inguinal region and lower limb
C1955687|T191|AB|200.36|ICD9CM|Margin zone lym pelvic|Margin zone lym pelvic
C1955687|T191|PT|200.36|ICD9CM|Marginal zone lymphoma, intrapelvic lymph nodes|Marginal zone lymphoma, intrapelvic lymph nodes
C0349632|T191|AB|200.37|ICD9CM|Margin zone lymph spleen|Margin zone lymph spleen
C0349632|T191|PT|200.37|ICD9CM|Marginal zone lymphoma, spleen|Marginal zone lymphoma, spleen
C1955689|T191|AB|200.38|ICD9CM|Margin zone lymph multip|Margin zone lymph multip
C1955689|T191|PT|200.38|ICD9CM|Marginal zone lymphoma, lymph nodes of multiple sites|Marginal zone lymphoma, lymph nodes of multiple sites
C4721414|T191|HT|200.4|ICD9CM|Mantle cell lymphoma|Mantle cell lymphoma
C1955691|T191|AB|200.40|ICD9CM|Mantle cell lym xtrrndl|Mantle cell lym xtrrndl
C1955691|T191|PT|200.40|ICD9CM|Mantle cell lymphoma, unspecified site, extranodal and solid organ sites|Mantle cell lymphoma, unspecified site, extranodal and solid organ sites
C2853895|T191|AB|200.41|ICD9CM|Mantle cell lymph head|Mantle cell lymph head
C2853895|T191|PT|200.41|ICD9CM|Mantle cell lymphoma, lymph nodes of head, face, and neck|Mantle cell lymphoma, lymph nodes of head, face, and neck
C2853896|T191|AB|200.42|ICD9CM|Mantle cell lymph thorax|Mantle cell lymph thorax
C2853896|T191|PT|200.42|ICD9CM|Mantle cell lymphoma, intrathoracic lymph nodes|Mantle cell lymphoma, intrathoracic lymph nodes
C2853897|T191|AB|200.43|ICD9CM|Mantle cell lymph abdom|Mantle cell lymph abdom
C2853897|T191|PT|200.43|ICD9CM|Mantle cell lymphoma, intra-abdominal lymph nodes|Mantle cell lymphoma, intra-abdominal lymph nodes
C2853898|T191|AB|200.44|ICD9CM|Mantle cell lymph axilla|Mantle cell lymph axilla
C2853898|T191|PT|200.44|ICD9CM|Mantle cell lymphoma, lymph nodes of axilla and upper limb|Mantle cell lymphoma, lymph nodes of axilla and upper limb
C2853899|T191|AB|200.45|ICD9CM|Mantle cell lymph inguin|Mantle cell lymph inguin
C2853899|T191|PT|200.45|ICD9CM|Mantle cell lymphoma, lymph nodes of inguinal region and lower limb|Mantle cell lymphoma, lymph nodes of inguinal region and lower limb
C2853900|T191|AB|200.46|ICD9CM|Mantle cell lymph pelvic|Mantle cell lymph pelvic
C2853900|T191|PT|200.46|ICD9CM|Mantle cell lymphoma, intrapelvic lymph nodes|Mantle cell lymphoma, intrapelvic lymph nodes
C2018777|T191|AB|200.47|ICD9CM|Mantle cell lymph spleen|Mantle cell lymph spleen
C2018777|T191|PT|200.47|ICD9CM|Mantle cell lymphoma, spleen|Mantle cell lymphoma, spleen
C2853901|T191|AB|200.48|ICD9CM|Mantle cell lymph multip|Mantle cell lymph multip
C2853901|T191|PT|200.48|ICD9CM|Mantle cell lymphoma, lymph nodes of multiple sites|Mantle cell lymphoma, lymph nodes of multiple sites
C0280803|T191|HT|200.5|ICD9CM|Primary central nervous system lymphoma|Primary central nervous system lymphoma
C1955700|T191|PT|200.50|ICD9CM|Primary central nervous system lymphoma, unspecified site, extranodal and solid organ sites|Primary central nervous system lymphoma, unspecified site, extranodal and solid organ sites
C1955700|T191|AB|200.50|ICD9CM|Primary CNS lymph xtrndl|Primary CNS lymph xtrndl
C1955701|T191|PT|200.51|ICD9CM|Primary central nervous system lymphoma, lymph nodes of head, face, and neck|Primary central nervous system lymphoma, lymph nodes of head, face, and neck
C1955701|T191|AB|200.51|ICD9CM|Primary CNS lymph head|Primary CNS lymph head
C1955702|T191|PT|200.52|ICD9CM|Primary central nervous system lymphoma, intrathoracic lymph nodes|Primary central nervous system lymphoma, intrathoracic lymph nodes
C1955702|T191|AB|200.52|ICD9CM|Primary CNS lymph thorax|Primary CNS lymph thorax
C1955703|T191|PT|200.53|ICD9CM|Primary central nervous system lymphoma, intra-abdominal lymph nodes|Primary central nervous system lymphoma, intra-abdominal lymph nodes
C1955703|T191|AB|200.53|ICD9CM|Primary CNS lymph abdom|Primary CNS lymph abdom
C1955704|T191|PT|200.54|ICD9CM|Primary central nervous system lymphoma, lymph nodes of axilla and upper limb|Primary central nervous system lymphoma, lymph nodes of axilla and upper limb
C1955704|T191|AB|200.54|ICD9CM|Primary CNS lymph axilla|Primary CNS lymph axilla
C1955705|T191|PT|200.55|ICD9CM|Primary central nervous system lymphoma, lymph nodes of inguinal region and lower limb|Primary central nervous system lymphoma, lymph nodes of inguinal region and lower limb
C1955705|T191|AB|200.55|ICD9CM|Primary CNS lym inguin|Primary CNS lym inguin
C1955706|T191|PT|200.56|ICD9CM|Primary central nervous system lymphoma, intrapelvic lymph nodes|Primary central nervous system lymphoma, intrapelvic lymph nodes
C1955706|T191|AB|200.56|ICD9CM|Primary CNS lymph pelvic|Primary CNS lymph pelvic
C1955707|T191|PT|200.57|ICD9CM|Primary central nervous system lymphoma, spleen|Primary central nervous system lymphoma, spleen
C1955707|T191|AB|200.57|ICD9CM|Primary CNS lymph spleen|Primary CNS lymph spleen
C1955708|T191|PT|200.58|ICD9CM|Primary central nervous system lymphoma, lymph nodes of multiple sites|Primary central nervous system lymphoma, lymph nodes of multiple sites
C1955708|T191|AB|200.58|ICD9CM|Primary CNS lymph multip|Primary CNS lymph multip
C0206180|T191|HT|200.6|ICD9CM|Anaplastic large cell lymphoma|Anaplastic large cell lymphoma
C1955709|T191|PT|200.60|ICD9CM|Anaplastic large cell lymphoma, unspecified site, extranodal and solid organ sites|Anaplastic large cell lymphoma, unspecified site, extranodal and solid organ sites
C1955709|T191|AB|200.60|ICD9CM|Anaplastic lymph xtrndl|Anaplastic lymph xtrndl
C1955710|T191|PT|200.61|ICD9CM|Anaplastic large cell lymphoma, lymph nodes of head, face, and neck|Anaplastic large cell lymphoma, lymph nodes of head, face, and neck
C1955710|T191|AB|200.61|ICD9CM|Anaplastic lymph head|Anaplastic lymph head
C1955711|T191|PT|200.62|ICD9CM|Anaplastic large cell lymphoma, intrathoracic lymph nodes|Anaplastic large cell lymphoma, intrathoracic lymph nodes
C1955711|T191|AB|200.62|ICD9CM|Anaplastic lymph thorax|Anaplastic lymph thorax
C1955712|T191|PT|200.63|ICD9CM|Anaplastic large cell lymphoma, intra-abdominal lymph nodes|Anaplastic large cell lymphoma, intra-abdominal lymph nodes
C1955712|T191|AB|200.63|ICD9CM|Anaplastic lymph abdom|Anaplastic lymph abdom
C1955713|T191|PT|200.64|ICD9CM|Anaplastic large cell lymphoma, lymph nodes of axilla and upper limb|Anaplastic large cell lymphoma, lymph nodes of axilla and upper limb
C1955713|T191|AB|200.64|ICD9CM|Anaplastic lymph axilla|Anaplastic lymph axilla
C1955714|T191|PT|200.65|ICD9CM|Anaplastic large cell lymphoma, lymph nodes of inguinal region and lower limb|Anaplastic large cell lymphoma, lymph nodes of inguinal region and lower limb
C1955714|T191|AB|200.65|ICD9CM|Anaplastic lymph inguin|Anaplastic lymph inguin
C1955715|T191|PT|200.66|ICD9CM|Anaplastic large cell lymphoma, intrapelvic lymph nodes|Anaplastic large cell lymphoma, intrapelvic lymph nodes
C1955715|T191|AB|200.66|ICD9CM|Anaplastic lymph pelvic|Anaplastic lymph pelvic
C2018768|T191|PT|200.67|ICD9CM|Anaplastic large cell lymphoma, spleen|Anaplastic large cell lymphoma, spleen
C2018768|T191|AB|200.67|ICD9CM|Anaplastic lymph spleen|Anaplastic lymph spleen
C1955717|T191|PT|200.68|ICD9CM|Anaplastic large cell lymphoma, lymph nodes of multiple sites|Anaplastic large cell lymphoma, lymph nodes of multiple sites
C1955717|T191|AB|200.68|ICD9CM|Anaplastic lymph multip|Anaplastic lymph multip
C0024302|T191|HT|200.7|ICD9CM|Large cell lymphoma|Large cell lymphoma
C1955718|T191|AB|200.70|ICD9CM|Large cell lymph xtrndl|Large cell lymph xtrndl
C1955718|T191|PT|200.70|ICD9CM|Large cell lymphoma, unspecified site, extranodal and solid organ sites|Large cell lymphoma, unspecified site, extranodal and solid organ sites
C1955719|T191|AB|200.71|ICD9CM|Large cell lymphoma head|Large cell lymphoma head
C1955719|T191|PT|200.71|ICD9CM|Large cell lymphoma, lymph nodes of head, face, and neck|Large cell lymphoma, lymph nodes of head, face, and neck
C1955720|T191|AB|200.72|ICD9CM|Large cell lymph thorax|Large cell lymph thorax
C1955720|T191|PT|200.72|ICD9CM|Large cell lymphoma, intrathoracic lymph nodes|Large cell lymphoma, intrathoracic lymph nodes
C1955721|T047|AB|200.73|ICD9CM|Large cell lymph abdom|Large cell lymph abdom
C1955721|T047|PT|200.73|ICD9CM|Large cell lymphoma, intra-abdominal lymph nodes|Large cell lymphoma, intra-abdominal lymph nodes
C1955722|T191|AB|200.74|ICD9CM|Large cell lymph axilla|Large cell lymph axilla
C1955722|T191|PT|200.74|ICD9CM|Large cell lymphoma, lymph nodes of axilla and upper limb|Large cell lymphoma, lymph nodes of axilla and upper limb
C1955723|T191|AB|200.75|ICD9CM|Large cell lymph inguin|Large cell lymph inguin
C1955723|T191|PT|200.75|ICD9CM|Large cell lymphoma, lymph nodes of inguinal region and lower limb|Large cell lymphoma, lymph nodes of inguinal region and lower limb
C2711042|T191|AB|200.76|ICD9CM|Large cell lymph pelvic|Large cell lymph pelvic
C2711042|T191|PT|200.76|ICD9CM|Large cell lymphoma, intrapelvic lymph nodes|Large cell lymphoma, intrapelvic lymph nodes
C1955725|T191|AB|200.77|ICD9CM|Large cell lymph spleen|Large cell lymph spleen
C1955725|T191|PT|200.77|ICD9CM|Large cell lymphoma, spleen|Large cell lymphoma, spleen
C1955726|T191|AB|200.78|ICD9CM|Large cell lymph multip|Large cell lymph multip
C1955726|T191|PT|200.78|ICD9CM|Large cell lymphoma, lymph nodes of multiple sites|Large cell lymphoma, lymph nodes of multiple sites
C0079955|T191|HT|200.8|ICD9CM|Other named variants of lymphosarcoma and reticulosarcoma|Other named variants of lymphosarcoma and reticulosarcoma
C0375078|T191|AB|200.80|ICD9CM|Oth varn unsp xtrndl org|Oth varn unsp xtrndl org
C0153720|T191|AB|200.81|ICD9CM|Mixed lymphosarc head|Mixed lymphosarc head
C0153720|T191|PT|200.81|ICD9CM|Other named variants of lymphosarcoma and reticulosarcoma, lymph nodes of head, face, and neck|Other named variants of lymphosarcoma and reticulosarcoma, lymph nodes of head, face, and neck
C0153721|T191|AB|200.82|ICD9CM|Mixed lymphosarc thorax|Mixed lymphosarc thorax
C0153721|T191|PT|200.82|ICD9CM|Other named variants of lymphosarcoma and reticulosarcoma,intrathoracic lymph nodes|Other named variants of lymphosarcoma and reticulosarcoma,intrathoracic lymph nodes
C0153722|T191|AB|200.83|ICD9CM|Mixed lymphosarc abdom|Mixed lymphosarc abdom
C0153722|T191|PT|200.83|ICD9CM|Other named variants of lymphosarcoma and reticulosarcoma, intra-abdominal lymph nodes|Other named variants of lymphosarcoma and reticulosarcoma, intra-abdominal lymph nodes
C0153723|T191|AB|200.84|ICD9CM|Mixed lymphosarc axilla|Mixed lymphosarc axilla
C0153723|T191|PT|200.84|ICD9CM|Other named variants of lymphosarcoma and reticulosarcoma, lymph nodes of axilla and upper limb|Other named variants of lymphosarcoma and reticulosarcoma, lymph nodes of axilla and upper limb
C0153724|T191|AB|200.85|ICD9CM|Mixed lymphosarc inguin|Mixed lymphosarc inguin
C0153725|T191|AB|200.86|ICD9CM|Mixed lymphosarc pelvic|Mixed lymphosarc pelvic
C0153725|T191|PT|200.86|ICD9CM|Other named variants of lymphosarcoma and reticulosarcoma, intrapelvic lymph nodes|Other named variants of lymphosarcoma and reticulosarcoma, intrapelvic lymph nodes
C0153726|T191|AB|200.87|ICD9CM|Mixed lymphosarc spleen|Mixed lymphosarc spleen
C0153726|T191|PT|200.87|ICD9CM|Other named variants of lymphosarcoma and reticulosarcoma, spleen|Other named variants of lymphosarcoma and reticulosarcoma, spleen
C0153727|T191|AB|200.88|ICD9CM|Mixed lymphosarc mult|Mixed lymphosarc mult
C0153727|T191|PT|200.88|ICD9CM|Other named variants of lymphosarcoma and reticulosarcoma, lymph nodes of multiple sites|Other named variants of lymphosarcoma and reticulosarcoma, lymph nodes of multiple sites
C0019829|T191|HT|201|ICD9CM|Hodgkin's disease|Hodgkin's disease
C0019829|T191|HT|201.0|ICD9CM|Hodgkin's paragranuloma|Hodgkin's paragranuloma
C0686560|T191|AB|201.00|ICD9CM|Hdgk prg unsp xtrndl org|Hdgk prg unsp xtrndl org
C0686560|T191|PT|201.00|ICD9CM|Hodgkin's paragranuloma, unspecified site, extranodal and solid organ sites|Hodgkin's paragranuloma, unspecified site, extranodal and solid organ sites
C0153728|T191|PT|201.01|ICD9CM|Hodgkin's paragranuloma, lymph nodes of head, face, and neck|Hodgkin's paragranuloma, lymph nodes of head, face, and neck
C0153728|T191|AB|201.01|ICD9CM|Hodgkins paragran head|Hodgkins paragran head
C0153729|T191|PT|201.02|ICD9CM|Hodgkin's paragranuloma, intrathoracic lymph nodes|Hodgkin's paragranuloma, intrathoracic lymph nodes
C0153729|T191|AB|201.02|ICD9CM|Hodgkins paragran thorax|Hodgkins paragran thorax
C0153730|T191|PT|201.03|ICD9CM|Hodgkin's paragranuloma, intra-abdominal lymph nodes|Hodgkin's paragranuloma, intra-abdominal lymph nodes
C0153730|T191|AB|201.03|ICD9CM|Hodgkins paragran abdom|Hodgkins paragran abdom
C0153731|T191|PT|201.04|ICD9CM|Hodgkin's paragranuloma, lymph nodes of axilla and upper limb|Hodgkin's paragranuloma, lymph nodes of axilla and upper limb
C0153731|T191|AB|201.04|ICD9CM|Hodgkins paragran axilla|Hodgkins paragran axilla
C0153732|T191|PT|201.05|ICD9CM|Hodgkin's paragranuloma, lymph nodes of inguinal region and lower limb|Hodgkin's paragranuloma, lymph nodes of inguinal region and lower limb
C0153732|T191|AB|201.05|ICD9CM|Hodgkins paragran inguin|Hodgkins paragran inguin
C0153733|T191|PT|201.06|ICD9CM|Hodgkin's paragranuloma, intrapelvic lymph nodes|Hodgkin's paragranuloma, intrapelvic lymph nodes
C0153733|T191|AB|201.06|ICD9CM|Hodgkins paragran pelvic|Hodgkins paragran pelvic
C0153734|T191|PT|201.07|ICD9CM|Hodgkin's paragranuloma, spleen|Hodgkin's paragranuloma, spleen
C0153734|T191|AB|201.07|ICD9CM|Hodgkins paragran spleen|Hodgkins paragran spleen
C0432534|T191|PT|201.08|ICD9CM|Hodgkin's paragranuloma, lymph nodes of multiple sites|Hodgkin's paragranuloma, lymph nodes of multiple sites
C0432534|T191|AB|201.08|ICD9CM|Hodgkins paragran mult|Hodgkins paragran mult
C0019829|T191|HT|201.1|ICD9CM|Hodgkin's granuloma|Hodgkin's granuloma
C0375080|T191|AB|201.10|ICD9CM|Hdgk grn unsp xtrndl org|Hdgk grn unsp xtrndl org
C0375080|T191|PT|201.10|ICD9CM|Hodgkin's granuloma, unspecified site, extranodal and solid organ sites|Hodgkin's granuloma, unspecified site, extranodal and solid organ sites
C0153736|T191|PT|201.11|ICD9CM|Hodgkin's granuloma, lymph nodes of head, face, and neck|Hodgkin's granuloma, lymph nodes of head, face, and neck
C0153736|T191|AB|201.11|ICD9CM|Hodgkins granulom head|Hodgkins granulom head
C0153737|T191|PT|201.12|ICD9CM|Hodgkin's granuloma, intrathoracic lymph nodes|Hodgkin's granuloma, intrathoracic lymph nodes
C0153737|T191|AB|201.12|ICD9CM|Hodgkins granulom thorax|Hodgkins granulom thorax
C0153738|T191|PT|201.13|ICD9CM|Hodgkin's granuloma, intra-abdominal lymph nodes|Hodgkin's granuloma, intra-abdominal lymph nodes
C0153738|T191|AB|201.13|ICD9CM|Hodgkins granulom abdom|Hodgkins granulom abdom
C0153739|T191|PT|201.14|ICD9CM|Hodgkin's granuloma, lymph nodes of axilla and upper limb|Hodgkin's granuloma, lymph nodes of axilla and upper limb
C0153739|T191|AB|201.14|ICD9CM|Hodgkins granulom axilla|Hodgkins granulom axilla
C0153740|T191|PT|201.15|ICD9CM|Hodgkin's granuloma, lymph nodes of inguinal region and lower limb|Hodgkin's granuloma, lymph nodes of inguinal region and lower limb
C0153740|T191|AB|201.15|ICD9CM|Hodgkins granulom inguin|Hodgkins granulom inguin
C0153741|T191|PT|201.16|ICD9CM|Hodgkin's granuloma, intrapelvic lymph nodes|Hodgkin's granuloma, intrapelvic lymph nodes
C0153741|T191|AB|201.16|ICD9CM|Hodgkins granulom pelvic|Hodgkins granulom pelvic
C0700143|T191|PT|201.17|ICD9CM|Hodgkin's granuloma, spleen|Hodgkin's granuloma, spleen
C0700143|T191|AB|201.17|ICD9CM|Hodgkins granulom spleen|Hodgkins granulom spleen
C0153742|T191|PT|201.18|ICD9CM|Hodgkin's granuloma, lymph nodes of multiple sites|Hodgkin's granuloma, lymph nodes of multiple sites
C0153742|T191|AB|201.18|ICD9CM|Hodgkins granulom mult|Hodgkins granulom mult
C0019829|T191|HT|201.2|ICD9CM|Hodgkin's sarcoma|Hodgkin's sarcoma
C0375081|T191|AB|201.20|ICD9CM|Hdgk src unsp xtrndl org|Hdgk src unsp xtrndl org
C0375081|T191|PT|201.20|ICD9CM|Hodgkin's sarcoma, unspecified site, extranodal and solid organ sites|Hodgkin's sarcoma, unspecified site, extranodal and solid organ sites
C0153744|T191|PT|201.21|ICD9CM|Hodgkin's sarcoma, lymph nodes of head, face, and neck|Hodgkin's sarcoma, lymph nodes of head, face, and neck
C0153744|T191|AB|201.21|ICD9CM|Hodgkins sarcoma head|Hodgkins sarcoma head
C0153745|T191|PT|201.22|ICD9CM|Hodgkin's sarcoma, intrathoracic lymph nodes|Hodgkin's sarcoma, intrathoracic lymph nodes
C0153745|T191|AB|201.22|ICD9CM|Hodgkins sarcoma thorax|Hodgkins sarcoma thorax
C0153746|T191|PT|201.23|ICD9CM|Hodgkin's sarcoma, intra-abdominal lymph nodes|Hodgkin's sarcoma, intra-abdominal lymph nodes
C0153746|T191|AB|201.23|ICD9CM|Hodgkins sarcoma abdom|Hodgkins sarcoma abdom
C0153747|T191|PT|201.24|ICD9CM|Hodgkin's sarcoma, lymph nodes of axilla and upper limb|Hodgkin's sarcoma, lymph nodes of axilla and upper limb
C0153747|T191|AB|201.24|ICD9CM|Hodgkins sarcoma axilla|Hodgkins sarcoma axilla
C0153748|T191|PT|201.25|ICD9CM|Hodgkin's sarcoma, lymph nodes of inguinal region and lower limb|Hodgkin's sarcoma, lymph nodes of inguinal region and lower limb
C0153748|T191|AB|201.25|ICD9CM|Hodgkins sarcoma inguin|Hodgkins sarcoma inguin
C0153749|T191|PT|201.26|ICD9CM|Hodgkin's sarcoma, intrapelvic lymph nodes|Hodgkin's sarcoma, intrapelvic lymph nodes
C0153749|T191|AB|201.26|ICD9CM|Hodgkins sarcoma pelvic|Hodgkins sarcoma pelvic
C0153750|T191|PT|201.27|ICD9CM|Hodgkin's sarcoma, spleen|Hodgkin's sarcoma, spleen
C0153750|T191|AB|201.27|ICD9CM|Hodgkins sarcoma spleen|Hodgkins sarcoma spleen
C0153751|T191|PT|201.28|ICD9CM|Hodgkin's sarcoma, lymph nodes of multiple sites|Hodgkin's sarcoma, lymph nodes of multiple sites
C0153751|T191|AB|201.28|ICD9CM|Hodgkins sarcoma mult|Hodgkins sarcoma mult
C1266194|T191|HT|201.4|ICD9CM|Hodgkin's disease, lymphocytic-histiocytic predominance|Hodgkin's disease, lymphocytic-histiocytic predominance
C0375082|T191|AB|201.40|ICD9CM|Lym-hst unsp xtrndl orgn|Lym-hst unsp xtrndl orgn
C0153752|T191|AB|201.41|ICD9CM|Hodg lymph-histio head|Hodg lymph-histio head
C0153752|T191|PT|201.41|ICD9CM|Hodgkin's disease, lymphocytic-histiocytic predominance, lymph nodes of head, face, and neck|Hodgkin's disease, lymphocytic-histiocytic predominance, lymph nodes of head, face, and neck
C0153753|T191|AB|201.42|ICD9CM|Hodg lymph-histio thorax|Hodg lymph-histio thorax
C0153753|T191|PT|201.42|ICD9CM|Hodgkin's disease, lymphocytic-histiocytic predominance, intrathoracic lymph nodes|Hodgkin's disease, lymphocytic-histiocytic predominance, intrathoracic lymph nodes
C0153754|T191|AB|201.43|ICD9CM|Hodg lymph-histio abdom|Hodg lymph-histio abdom
C0153754|T191|PT|201.43|ICD9CM|Hodgkin's disease, lymphocytic-histiocytic predominance, intra-abdominal lymph nodes|Hodgkin's disease, lymphocytic-histiocytic predominance, intra-abdominal lymph nodes
C0153755|T191|AB|201.44|ICD9CM|Hodg lymph-histio axilla|Hodg lymph-histio axilla
C0153755|T191|PT|201.44|ICD9CM|Hodgkin's disease, lymphocytic-histiocytic predominance, lymph nodes of axilla and upper limb|Hodgkin's disease, lymphocytic-histiocytic predominance, lymph nodes of axilla and upper limb
C0153756|T191|AB|201.45|ICD9CM|Hodg lymph-histio inguin|Hodg lymph-histio inguin
C0153757|T191|AB|201.46|ICD9CM|Hodg lymph-histio pelvic|Hodg lymph-histio pelvic
C0153757|T191|PT|201.46|ICD9CM|Hodgkin's disease, lymphocytic-histiocytic predominance, intrapelvic lymph nodes|Hodgkin's disease, lymphocytic-histiocytic predominance, intrapelvic lymph nodes
C0153758|T191|AB|201.47|ICD9CM|Hodg lymph-histio spleen|Hodg lymph-histio spleen
C0153758|T191|PT|201.47|ICD9CM|Hodgkin's disease, lymphocytic-histiocytic predominance, spleen|Hodgkin's disease, lymphocytic-histiocytic predominance, spleen
C0153759|T191|AB|201.48|ICD9CM|Hodg lymph-histio mult|Hodg lymph-histio mult
C0153759|T191|PT|201.48|ICD9CM|Hodgkin's disease, lymphocytic-histiocytic predominance, lymph nodes of multiple sites|Hodgkin's disease, lymphocytic-histiocytic predominance, lymph nodes of multiple sites
C0152268|T191|HT|201.5|ICD9CM|Hodgkin's disease, nodular sclerosis|Hodgkin's disease, nodular sclerosis
C0375083|T191|PT|201.50|ICD9CM|Hodgkin's disease, nodular sclerosis, unspecified site, extranodal and solid organ sites|Hodgkin's disease, nodular sclerosis, unspecified site, extranodal and solid organ sites
C0375083|T191|AB|201.50|ICD9CM|Ndr sclr unsp xtrndl org|Ndr sclr unsp xtrndl org
C0153760|T191|AB|201.51|ICD9CM|Hodg nodul sclero head|Hodg nodul sclero head
C0153760|T191|PT|201.51|ICD9CM|Hodgkin's disease, nodular sclerosis, lymph nodes of head, face, and neck|Hodgkin's disease, nodular sclerosis, lymph nodes of head, face, and neck
C0153761|T191|AB|201.52|ICD9CM|Hodg nodul sclero thorax|Hodg nodul sclero thorax
C0153761|T191|PT|201.52|ICD9CM|Hodgkin's disease, nodular sclerosis, intrathoracic lymph nodes|Hodgkin's disease, nodular sclerosis, intrathoracic lymph nodes
C0153762|T191|AB|201.53|ICD9CM|Hodg nodul sclero abdom|Hodg nodul sclero abdom
C0153762|T191|PT|201.53|ICD9CM|Hodgkin's disease, nodular sclerosis, intra-abdominal lymph nodes|Hodgkin's disease, nodular sclerosis, intra-abdominal lymph nodes
C0153763|T191|AB|201.54|ICD9CM|Hodg nodul sclero axilla|Hodg nodul sclero axilla
C0153763|T191|PT|201.54|ICD9CM|Hodgkin's disease, nodular sclerosis, lymph nodes of axilla and upper limb|Hodgkin's disease, nodular sclerosis, lymph nodes of axilla and upper limb
C0153764|T191|AB|201.55|ICD9CM|Hodg nodul sclero inguin|Hodg nodul sclero inguin
C0153764|T191|PT|201.55|ICD9CM|Hodgkin's disease, nodular sclerosis, lymph nodes of inguinal region and lower limb|Hodgkin's disease, nodular sclerosis, lymph nodes of inguinal region and lower limb
C0153765|T191|AB|201.56|ICD9CM|Hodg nodul sclero pelvic|Hodg nodul sclero pelvic
C0153765|T191|PT|201.56|ICD9CM|Hodgkin's disease, nodular sclerosis, intrapelvic lymph nodes|Hodgkin's disease, nodular sclerosis, intrapelvic lymph nodes
C0153766|T191|AB|201.57|ICD9CM|Hodg nodul sclero spleen|Hodg nodul sclero spleen
C0153766|T191|PT|201.57|ICD9CM|Hodgkin's disease, nodular sclerosis, spleen|Hodgkin's disease, nodular sclerosis, spleen
C0153767|T191|AB|201.58|ICD9CM|Hodg nodul sclero mult|Hodg nodul sclero mult
C0153767|T191|PT|201.58|ICD9CM|Hodgkin's disease, nodular sclerosis, lymph nodes of multiple sites|Hodgkin's disease, nodular sclerosis, lymph nodes of multiple sites
C0152266|T191|HT|201.6|ICD9CM|Hodgkin's disease, mixed cellularity|Hodgkin's disease, mixed cellularity
C0375084|T191|PT|201.60|ICD9CM|Hodgkin's disease, mixed cellularity, unspecified site, extranodal and solid organ sites|Hodgkin's disease, mixed cellularity, unspecified site, extranodal and solid organ sites
C0375084|T191|AB|201.60|ICD9CM|Mxd celr unsp xtrndl org|Mxd celr unsp xtrndl org
C0153768|T191|PT|201.61|ICD9CM|Hodgkin's disease, mixed cellularity, lymph nodes of head, face, and neck|Hodgkin's disease, mixed cellularity, lymph nodes of head, face, and neck
C0153768|T191|AB|201.61|ICD9CM|Hodgkins mix cell head|Hodgkins mix cell head
C0153769|T191|PT|201.62|ICD9CM|Hodgkin's disease, mixed cellularity, intrathoracic lymph nodes|Hodgkin's disease, mixed cellularity, intrathoracic lymph nodes
C0153769|T191|AB|201.62|ICD9CM|Hodgkins mix cell thorax|Hodgkins mix cell thorax
C0153770|T191|PT|201.63|ICD9CM|Hodgkin's disease, mixed cellularity, intra-abdominal lymph nodes|Hodgkin's disease, mixed cellularity, intra-abdominal lymph nodes
C0153770|T191|AB|201.63|ICD9CM|Hodgkins mix cell abdom|Hodgkins mix cell abdom
C0153771|T191|PT|201.64|ICD9CM|Hodgkin's disease, mixed cellularity, lymph nodes of axilla and upper limb|Hodgkin's disease, mixed cellularity, lymph nodes of axilla and upper limb
C0153771|T191|AB|201.64|ICD9CM|Hodgkins mix cell axilla|Hodgkins mix cell axilla
C0153772|T191|PT|201.65|ICD9CM|Hodgkin's disease, mixed cellularity, lymph nodes of inguinal region and lower limb|Hodgkin's disease, mixed cellularity, lymph nodes of inguinal region and lower limb
C0153772|T191|AB|201.65|ICD9CM|Hodgkins mix cell inguin|Hodgkins mix cell inguin
C0153773|T191|PT|201.66|ICD9CM|Hodgkin's disease, mixed cellularity, intrapelvic lymph nodes|Hodgkin's disease, mixed cellularity, intrapelvic lymph nodes
C0153773|T191|AB|201.66|ICD9CM|Hodgkins mix cell pelvic|Hodgkins mix cell pelvic
C0153774|T191|PT|201.67|ICD9CM|Hodgkin's disease, mixed cellularity, spleen|Hodgkin's disease, mixed cellularity, spleen
C0153774|T191|AB|201.67|ICD9CM|Hodgkins mix cell spleen|Hodgkins mix cell spleen
C0153775|T191|PT|201.68|ICD9CM|Hodgkin's disease, mixed cellularity, lymph nodes of multiple sites|Hodgkin's disease, mixed cellularity, lymph nodes of multiple sites
C0153775|T191|AB|201.68|ICD9CM|Hodgkins mix cell mult|Hodgkins mix cell mult
C0152267|T191|HT|201.7|ICD9CM|Hodgkin's disease, lymphocytic depletion|Hodgkin's disease, lymphocytic depletion
C0375085|T191|PT|201.70|ICD9CM|Hodgkin's disease, lymphocytic depletion, unspecified site, extranodal and solid organ sites|Hodgkin's disease, lymphocytic depletion, unspecified site, extranodal and solid organ sites
C0375085|T191|AB|201.70|ICD9CM|Lym dplt unsp xtrndl org|Lym dplt unsp xtrndl org
C0153776|T191|AB|201.71|ICD9CM|Hodg lymph deplet head|Hodg lymph deplet head
C0153776|T191|PT|201.71|ICD9CM|Hodgkin's disease, lymphocytic depletion, lymph nodes of head, face, and neck|Hodgkin's disease, lymphocytic depletion, lymph nodes of head, face, and neck
C0153777|T191|AB|201.72|ICD9CM|Hodg lymph deplet thorax|Hodg lymph deplet thorax
C0153777|T191|PT|201.72|ICD9CM|Hodgkin's disease, lymphocytic depletion, intrathoracic lymph nodes|Hodgkin's disease, lymphocytic depletion, intrathoracic lymph nodes
C0153778|T191|AB|201.73|ICD9CM|Hodg lymph deplet abdom|Hodg lymph deplet abdom
C0153778|T191|PT|201.73|ICD9CM|Hodgkin's disease, lymphocytic depletion, intra-abdominal lymph nodes|Hodgkin's disease, lymphocytic depletion, intra-abdominal lymph nodes
C0153779|T191|AB|201.74|ICD9CM|Hodg lymph deplet axilla|Hodg lymph deplet axilla
C0153779|T191|PT|201.74|ICD9CM|Hodgkin's disease, lymphocytic depletion, lymph nodes of axilla and upper limb|Hodgkin's disease, lymphocytic depletion, lymph nodes of axilla and upper limb
C0153780|T191|AB|201.75|ICD9CM|Hodg lymph deplet inguin|Hodg lymph deplet inguin
C0153780|T191|PT|201.75|ICD9CM|Hodgkin's disease, lymphocytic depletion, lymph nodes of inguinal region and lower limb|Hodgkin's disease, lymphocytic depletion, lymph nodes of inguinal region and lower limb
C0153781|T191|AB|201.76|ICD9CM|Hodg lymph deplet pelvic|Hodg lymph deplet pelvic
C0153781|T191|PT|201.76|ICD9CM|Hodgkin's disease, lymphocytic depletion, intrapelvic lymph nodes|Hodgkin's disease, lymphocytic depletion, intrapelvic lymph nodes
C0153782|T191|AB|201.77|ICD9CM|Hodg lymph deplet spleen|Hodg lymph deplet spleen
C0153782|T191|PT|201.77|ICD9CM|Hodgkin's disease, lymphocytic depletion, spleen|Hodgkin's disease, lymphocytic depletion, spleen
C0153783|T191|AB|201.78|ICD9CM|Hodg lymph deplet mult|Hodg lymph deplet mult
C0153783|T191|PT|201.78|ICD9CM|Hodgkin's disease, lymphocytic depletion, lymph nodes of multiple sites|Hodgkin's disease, lymphocytic depletion, lymph nodes of multiple sites
C0019829|T191|HT|201.9|ICD9CM|Hodgkin's disease, unspecified type|Hodgkin's disease, unspecified type
C0375086|T191|AB|201.90|ICD9CM|Hdgk dis unsp xtrndl org|Hdgk dis unsp xtrndl org
C0375086|T191|PT|201.90|ICD9CM|Hodgkin's disease, unspecified type, unspecified site, extranodal and solid organ sites|Hodgkin's disease, unspecified type, unspecified site, extranodal and solid organ sites
C0153785|T191|PT|201.91|ICD9CM|Hodgkin's disease, unspecified type, lymph nodes of head, face, and neck|Hodgkin's disease, unspecified type, lymph nodes of head, face, and neck
C0153785|T191|AB|201.91|ICD9CM|Hodgkins dis NOS head|Hodgkins dis NOS head
C0153786|T191|PT|201.92|ICD9CM|Hodgkin's disease, unspecified type, intrathoracic lymph nodes|Hodgkin's disease, unspecified type, intrathoracic lymph nodes
C0153786|T191|AB|201.92|ICD9CM|Hodgkins dis NOS thorax|Hodgkins dis NOS thorax
C1306638|T191|PT|201.93|ICD9CM|Hodgkin's disease, unspecified type, intra-abdominal lymph nodes|Hodgkin's disease, unspecified type, intra-abdominal lymph nodes
C1306638|T191|AB|201.93|ICD9CM|Hodgkins dis NOS abdom|Hodgkins dis NOS abdom
C0153788|T191|PT|201.94|ICD9CM|Hodgkin's disease, unspecified type, lymph nodes of axilla and upper limb|Hodgkin's disease, unspecified type, lymph nodes of axilla and upper limb
C0153788|T191|AB|201.94|ICD9CM|Hodgkins dis NOS axilla|Hodgkins dis NOS axilla
C0153789|T191|PT|201.95|ICD9CM|Hodgkin's disease, unspecified type, lymph nodes of inguinal region and lower limb|Hodgkin's disease, unspecified type, lymph nodes of inguinal region and lower limb
C0153789|T191|AB|201.95|ICD9CM|Hodgkins dis NOS inguin|Hodgkins dis NOS inguin
C0153790|T191|PT|201.96|ICD9CM|Hodgkin's disease, unspecified type, intrapelvic lymph nodes|Hodgkin's disease, unspecified type, intrapelvic lymph nodes
C0153790|T191|AB|201.96|ICD9CM|Hodgkins dis NOS pelvic|Hodgkins dis NOS pelvic
C0153791|T191|PT|201.97|ICD9CM|Hodgkin's disease, unspecified type, spleen|Hodgkin's disease, unspecified type, spleen
C0153791|T191|AB|201.97|ICD9CM|Hodgkins dis NOS spleen|Hodgkins dis NOS spleen
C0153792|T191|PT|201.98|ICD9CM|Hodgkin's disease, unspecified type, lymph nodes of multiple sites|Hodgkin's disease, unspecified type, lymph nodes of multiple sites
C0153792|T191|AB|201.98|ICD9CM|Hodgkins dis NOS mult|Hodgkins dis NOS mult
C0153793|T191|HT|202|ICD9CM|Other malignant neoplasms of lymphoid and histiocytic tissue|Other malignant neoplasms of lymphoid and histiocytic tissue
C0024301|T191|HT|202.0|ICD9CM|Nodular lymphoma|Nodular lymphoma
C0375087|T191|AB|202.00|ICD9CM|Ndlr lym unsp xtrndl org|Ndlr lym unsp xtrndl org
C0375087|T191|PT|202.00|ICD9CM|Nodular lymphoma, unspecified site, extranodal and solid organ sites|Nodular lymphoma, unspecified site, extranodal and solid organ sites
C0153794|T191|AB|202.01|ICD9CM|Nodular lymphoma head|Nodular lymphoma head
C0153794|T191|PT|202.01|ICD9CM|Nodular lymphoma, lymph nodes of head, face, and neck|Nodular lymphoma, lymph nodes of head, face, and neck
C0153795|T191|AB|202.02|ICD9CM|Nodular lymphoma thorax|Nodular lymphoma thorax
C0153795|T191|PT|202.02|ICD9CM|Nodular lymphoma, intrathoracic lymph nodes|Nodular lymphoma, intrathoracic lymph nodes
C0153796|T191|AB|202.03|ICD9CM|Nodular lymphoma abdom|Nodular lymphoma abdom
C0153796|T191|PT|202.03|ICD9CM|Nodular lymphoma, intra-abdominal lymph nodes|Nodular lymphoma, intra-abdominal lymph nodes
C0153797|T191|AB|202.04|ICD9CM|Nodular lymphoma axilla|Nodular lymphoma axilla
C0153797|T191|PT|202.04|ICD9CM|Nodular lymphoma, lymph nodes of axilla and upper limb|Nodular lymphoma, lymph nodes of axilla and upper limb
C0153798|T191|AB|202.05|ICD9CM|Nodular lymphoma inguin|Nodular lymphoma inguin
C0153798|T191|PT|202.05|ICD9CM|Nodular lymphoma, lymph nodes of inguinal region and lower limb|Nodular lymphoma, lymph nodes of inguinal region and lower limb
C0153799|T191|AB|202.06|ICD9CM|Nodular lymphoma pelvic|Nodular lymphoma pelvic
C0153799|T191|PT|202.06|ICD9CM|Nodular lymphoma, intrapelvic lymph nodes|Nodular lymphoma, intrapelvic lymph nodes
C0153800|T191|AB|202.07|ICD9CM|Nodular lymphoma spleen|Nodular lymphoma spleen
C0153800|T191|PT|202.07|ICD9CM|Nodular lymphoma, spleen|Nodular lymphoma, spleen
C0153801|T191|AB|202.08|ICD9CM|Nodular lymphoma mult|Nodular lymphoma mult
C0153801|T191|PT|202.08|ICD9CM|Nodular lymphoma, lymph nodes of multiple sites|Nodular lymphoma, lymph nodes of multiple sites
C0026948|T191|HT|202.1|ICD9CM|Mycosis fungoides|Mycosis fungoides
C0375088|T191|PT|202.10|ICD9CM|Mycosis fungoides, unspecified site, extranodal and solid organ sites|Mycosis fungoides, unspecified site, extranodal and solid organ sites
C0375088|T191|AB|202.10|ICD9CM|Mycs fng unsp xtrndl org|Mycs fng unsp xtrndl org
C0153802|T191|AB|202.11|ICD9CM|Mycosis fungoides head|Mycosis fungoides head
C0153802|T191|PT|202.11|ICD9CM|Mycosis fungoides, lymph nodes of head, face, and neck|Mycosis fungoides, lymph nodes of head, face, and neck
C0153803|T191|AB|202.12|ICD9CM|Mycosis fungoides thorax|Mycosis fungoides thorax
C0153803|T191|PT|202.12|ICD9CM|Mycosis fungoides, intrathoracic lymph nodes|Mycosis fungoides, intrathoracic lymph nodes
C0153804|T191|AB|202.13|ICD9CM|Mycosis fungoides abdom|Mycosis fungoides abdom
C0153804|T191|PT|202.13|ICD9CM|Mycosis fungoides, intra-abdominal lymph nodes|Mycosis fungoides, intra-abdominal lymph nodes
C0153805|T191|AB|202.14|ICD9CM|Mycosis fungoides axilla|Mycosis fungoides axilla
C0153805|T191|PT|202.14|ICD9CM|Mycosis fungoides, lymph nodes of axilla and upper limb|Mycosis fungoides, lymph nodes of axilla and upper limb
C0153806|T191|AB|202.15|ICD9CM|Mycosis fungoides inguin|Mycosis fungoides inguin
C0153806|T191|PT|202.15|ICD9CM|Mycosis fungoides, lymph nodes of inguinal region and lower limb|Mycosis fungoides, lymph nodes of inguinal region and lower limb
C0153807|T191|AB|202.16|ICD9CM|Mycosis fungoides pelvic|Mycosis fungoides pelvic
C0153807|T191|PT|202.16|ICD9CM|Mycosis fungoides, intrapelvic lymph nodes|Mycosis fungoides, intrapelvic lymph nodes
C0153808|T191|AB|202.17|ICD9CM|Mycosis fungoides spleen|Mycosis fungoides spleen
C0153808|T191|PT|202.17|ICD9CM|Mycosis fungoides, spleen|Mycosis fungoides, spleen
C0153809|T191|AB|202.18|ICD9CM|Mycosis fungoides mult|Mycosis fungoides mult
C0153809|T191|PT|202.18|ICD9CM|Mycosis fungoides, lymph nodes of multiple sites|Mycosis fungoides, lymph nodes of multiple sites
C0036920|T191|HT|202.2|ICD9CM|Sezary's disease|Sezary's disease
C0375089|T191|PT|202.20|ICD9CM|Sezary's disease, unspecified site, extranodal and solid organ sites|Sezary's disease, unspecified site, extranodal and solid organ sites
C0375089|T191|AB|202.20|ICD9CM|Szry dis unsp xtrndl org|Szry dis unsp xtrndl org
C0153810|T191|AB|202.21|ICD9CM|Sezary's disease head|Sezary's disease head
C0153810|T191|PT|202.21|ICD9CM|Sezary's disease, lymph nodes of head, face, and neck|Sezary's disease, lymph nodes of head, face, and neck
C0153811|T191|AB|202.22|ICD9CM|Sezary's disease thorax|Sezary's disease thorax
C0153811|T191|PT|202.22|ICD9CM|Sezary's disease, intrathoracic lymph nodes|Sezary's disease, intrathoracic lymph nodes
C0153812|T191|AB|202.23|ICD9CM|Sezary's disease abdom|Sezary's disease abdom
C0153812|T191|PT|202.23|ICD9CM|Sezary's disease, intra-abdominal lymph nodes|Sezary's disease, intra-abdominal lymph nodes
C0153813|T191|AB|202.24|ICD9CM|Sezary's disease axilla|Sezary's disease axilla
C0153813|T191|PT|202.24|ICD9CM|Sezary's disease, lymph nodes of axilla and upper limb|Sezary's disease, lymph nodes of axilla and upper limb
C0153814|T191|AB|202.25|ICD9CM|Sezary's disease inguin|Sezary's disease inguin
C0153814|T191|PT|202.25|ICD9CM|Sezary's disease, lymph nodes of inguinal region and lower limb|Sezary's disease, lymph nodes of inguinal region and lower limb
C0153815|T191|AB|202.26|ICD9CM|Sezary's disease pelvic|Sezary's disease pelvic
C0153815|T191|PT|202.26|ICD9CM|Sezary's disease, intrapelvic lymph nodes|Sezary's disease, intrapelvic lymph nodes
C0153816|T191|AB|202.27|ICD9CM|Sezary's disease spleen|Sezary's disease spleen
C0153816|T191|PT|202.27|ICD9CM|Sezary's disease, spleen|Sezary's disease, spleen
C0153817|T191|AB|202.28|ICD9CM|Sezary's disease mult|Sezary's disease mult
C0153817|T191|PT|202.28|ICD9CM|Sezary's disease, lymph nodes of multiple sites|Sezary's disease, lymph nodes of multiple sites
C0019623|T191|HT|202.3|ICD9CM|Malignant histiocytosis|Malignant histiocytosis
C0375090|T191|PT|202.30|ICD9CM|Malignant histiocytosis, unspecified site, extranodal and solid organ sites|Malignant histiocytosis, unspecified site, extranodal and solid organ sites
C0375090|T191|AB|202.30|ICD9CM|Mlg hist unsp xtrndl org|Mlg hist unsp xtrndl org
C0432538|T191|AB|202.31|ICD9CM|Mal histiocytosis head|Mal histiocytosis head
C0432538|T191|PT|202.31|ICD9CM|Malignant histiocytosis, lymph nodes of head, face, and neck|Malignant histiocytosis, lymph nodes of head, face, and neck
C0432539|T191|AB|202.32|ICD9CM|Mal histiocytosis thorax|Mal histiocytosis thorax
C0432539|T191|PT|202.32|ICD9CM|Malignant histiocytosis, intrathoracic lymph nodes|Malignant histiocytosis, intrathoracic lymph nodes
C0432540|T191|AB|202.33|ICD9CM|Mal histiocytosis abdom|Mal histiocytosis abdom
C0432540|T191|PT|202.33|ICD9CM|Malignant histiocytosis, intra-abdominal lymph nodes|Malignant histiocytosis, intra-abdominal lymph nodes
C0432541|T191|AB|202.34|ICD9CM|Mal histiocytosis axilla|Mal histiocytosis axilla
C0432541|T191|PT|202.34|ICD9CM|Malignant histiocytosis, lymph nodes of axilla and upper limb|Malignant histiocytosis, lymph nodes of axilla and upper limb
C0432542|T191|AB|202.35|ICD9CM|Mal histiocytosis inguin|Mal histiocytosis inguin
C0432542|T191|PT|202.35|ICD9CM|Malignant histiocytosis, lymph nodes of inguinal region and lower limb|Malignant histiocytosis, lymph nodes of inguinal region and lower limb
C0432543|T191|AB|202.36|ICD9CM|Mal histiocytosis pelvic|Mal histiocytosis pelvic
C0432543|T191|PT|202.36|ICD9CM|Malignant histiocytosis, intrapelvic lymph nodes|Malignant histiocytosis, intrapelvic lymph nodes
C0432544|T191|AB|202.37|ICD9CM|Mal histiocytosis spleen|Mal histiocytosis spleen
C0432544|T191|PT|202.37|ICD9CM|Malignant histiocytosis, spleen|Malignant histiocytosis, spleen
C0432545|T191|AB|202.38|ICD9CM|Mal histiocytosis mult|Mal histiocytosis mult
C0432545|T191|PT|202.38|ICD9CM|Malignant histiocytosis, lymph nodes of multiple sites|Malignant histiocytosis, lymph nodes of multiple sites
C0023443|T191|HT|202.4|ICD9CM|Leukemic reticuloendotheliosis|Leukemic reticuloendotheliosis
C0375091|T191|PT|202.40|ICD9CM|Leukemic reticuloendotheliosis, unspecified site, extranodal and solid organ sites|Leukemic reticuloendotheliosis, unspecified site, extranodal and solid organ sites
C0375091|T191|AB|202.40|ICD9CM|Lk rtctl unsp xtrndl org|Lk rtctl unsp xtrndl org
C0153826|T191|AB|202.41|ICD9CM|Hairy-cell leukem head|Hairy-cell leukem head
C0153826|T191|PT|202.41|ICD9CM|Leukemic reticuloendotheliosis, lymph nodes of head, face, and neck|Leukemic reticuloendotheliosis, lymph nodes of head, face, and neck
C0153827|T191|AB|202.42|ICD9CM|Hairy-cell leukem thorax|Hairy-cell leukem thorax
C0153827|T191|PT|202.42|ICD9CM|Leukemic reticuloendotheliosis, intrathoracic lymph nodes|Leukemic reticuloendotheliosis, intrathoracic lymph nodes
C0153828|T191|AB|202.43|ICD9CM|Hairy-cell leukem abdom|Hairy-cell leukem abdom
C0153828|T191|PT|202.43|ICD9CM|Leukemic reticuloendotheliosis, intra-abdominal lymph nodes|Leukemic reticuloendotheliosis, intra-abdominal lymph nodes
C0153829|T191|AB|202.44|ICD9CM|Hairy-cell leukem axilla|Hairy-cell leukem axilla
C0153829|T191|PT|202.44|ICD9CM|Leukemic reticuloendotheliosis, lymph nodes of axilla and upper arm|Leukemic reticuloendotheliosis, lymph nodes of axilla and upper arm
C0153830|T191|AB|202.45|ICD9CM|Hairy-cell leukem inguin|Hairy-cell leukem inguin
C0153830|T191|PT|202.45|ICD9CM|Leukemic reticuloendotheliosis, lymph nodes of inguinal region and lower limb|Leukemic reticuloendotheliosis, lymph nodes of inguinal region and lower limb
C0153831|T191|AB|202.46|ICD9CM|Hairy-cell leukem pelvic|Hairy-cell leukem pelvic
C0153831|T191|PT|202.46|ICD9CM|Leukemic reticuloendotheliosis, intrapelvic lymph nodes|Leukemic reticuloendotheliosis, intrapelvic lymph nodes
C0153832|T191|AB|202.47|ICD9CM|Hairy-cell leukem spleen|Hairy-cell leukem spleen
C0153832|T191|PT|202.47|ICD9CM|Leukemic reticuloendotheliosis, spleen|Leukemic reticuloendotheliosis, spleen
C0153833|T191|AB|202.48|ICD9CM|Hairy-cell leukem mult|Hairy-cell leukem mult
C0153833|T191|PT|202.48|ICD9CM|Leukemic reticuloendotheliosis, lymph nodes of multiple sites|Leukemic reticuloendotheliosis, lymph nodes of multiple sites
C0023381|T047|HT|202.5|ICD9CM|Letterer-Siwe disease|Letterer-Siwe disease
C0375092|T191|PT|202.50|ICD9CM|Letterer-siwe disease, unspecified site, extranodal and solid organ sites|Letterer-siwe disease, unspecified site, extranodal and solid organ sites
C0375092|T191|AB|202.50|ICD9CM|Ltr-siwe unsp xtrndl org|Ltr-siwe unsp xtrndl org
C0432547|T191|AB|202.51|ICD9CM|Letterer-siwe dis head|Letterer-siwe dis head
C0432547|T191|PT|202.51|ICD9CM|Letterer-siwe disease, lymph nodes of head, face, and neck|Letterer-siwe disease, lymph nodes of head, face, and neck
C0432548|T191|AB|202.52|ICD9CM|Letterer-siwe dis thorax|Letterer-siwe dis thorax
C0432548|T191|PT|202.52|ICD9CM|Letterer-siwe disease, intrathoracic lymph nodes|Letterer-siwe disease, intrathoracic lymph nodes
C0432549|T191|AB|202.53|ICD9CM|Letterer-siwe dis abdom|Letterer-siwe dis abdom
C0432549|T191|PT|202.53|ICD9CM|Letterer-siwe disease, intra-abdominal lymph nodes|Letterer-siwe disease, intra-abdominal lymph nodes
C0432550|T191|AB|202.54|ICD9CM|Letterer-siwe dis axilla|Letterer-siwe dis axilla
C0432550|T191|PT|202.54|ICD9CM|Letterer-siwe disease, lymph nodes of axilla and upper limb|Letterer-siwe disease, lymph nodes of axilla and upper limb
C0432551|T191|AB|202.55|ICD9CM|Letterer-siwe dis inguin|Letterer-siwe dis inguin
C0432551|T191|PT|202.55|ICD9CM|Letterer-siwe disease, lymph nodes of inguinal region and lower limb|Letterer-siwe disease, lymph nodes of inguinal region and lower limb
C0432552|T191|AB|202.56|ICD9CM|Letterer-siwe dis pelvic|Letterer-siwe dis pelvic
C0432552|T191|PT|202.56|ICD9CM|Letterer-siwe disease, intrapelvic lymph nodes|Letterer-siwe disease, intrapelvic lymph nodes
C0432553|T191|AB|202.57|ICD9CM|Letterer-siwe dis spleen|Letterer-siwe dis spleen
C0432553|T191|PT|202.57|ICD9CM|Letterer-siwe disease, spleen|Letterer-siwe disease, spleen
C0432554|T191|AB|202.58|ICD9CM|Letterer-siwe dis mult|Letterer-siwe dis mult
C0432554|T191|PT|202.58|ICD9CM|Letterer-siwe disease, lymph nodes of multiple sites|Letterer-siwe disease, lymph nodes of multiple sites
C0036221|T191|HT|202.6|ICD9CM|Malignant mast cell tumors|Malignant mast cell tumors
C0375093|T191|PT|202.60|ICD9CM|Malignant mast cell tumors, unspecified site, extranodal and solid organ sites|Malignant mast cell tumors, unspecified site, extranodal and solid organ sites
C0375093|T191|AB|202.60|ICD9CM|Mlg mast unsp xtrndl org|Mlg mast unsp xtrndl org
C0686574|T191|AB|202.61|ICD9CM|Mal mastocytosis head|Mal mastocytosis head
C0686574|T191|PT|202.61|ICD9CM|Malignant mast cell tumors, lymph nodes of head, face, and neck|Malignant mast cell tumors, lymph nodes of head, face, and neck
C0153843|T191|AB|202.62|ICD9CM|Mal mastocytosis thorax|Mal mastocytosis thorax
C0153843|T191|PT|202.62|ICD9CM|Malignant mast cell tumors, intrathoracic lymph nodes|Malignant mast cell tumors, intrathoracic lymph nodes
C0153844|T191|AB|202.63|ICD9CM|Mal mastocytosis abdom|Mal mastocytosis abdom
C0153844|T191|PT|202.63|ICD9CM|Malignant mast cell tumors, intra-abdominal lymph nodes|Malignant mast cell tumors, intra-abdominal lymph nodes
C0153845|T191|AB|202.64|ICD9CM|Mal mastocytosis axilla|Mal mastocytosis axilla
C0153845|T191|PT|202.64|ICD9CM|Malignant mast cell tumors, lymph nodes of axilla and upper limb|Malignant mast cell tumors, lymph nodes of axilla and upper limb
C0153846|T191|AB|202.65|ICD9CM|Mal mastocytosis inguin|Mal mastocytosis inguin
C0153846|T191|PT|202.65|ICD9CM|Malignant mast cell tumors, lymph nodes of inguinal region and lower limb|Malignant mast cell tumors, lymph nodes of inguinal region and lower limb
C0153847|T191|AB|202.66|ICD9CM|Mal mastocytosis pelvic|Mal mastocytosis pelvic
C0153847|T191|PT|202.66|ICD9CM|Malignant mast cell tumors, intrapelvic lymph nodes|Malignant mast cell tumors, intrapelvic lymph nodes
C0153848|T191|AB|202.67|ICD9CM|Mal mastocytosis spleen|Mal mastocytosis spleen
C0153848|T191|PT|202.67|ICD9CM|Malignant mast cell tumors, spleen|Malignant mast cell tumors, spleen
C0153849|T191|AB|202.68|ICD9CM|Mal mastocytosis mult|Mal mastocytosis mult
C0153849|T191|PT|202.68|ICD9CM|Malignant mast cell tumors, lymph nodes of multiple sites|Malignant mast cell tumors, lymph nodes of multiple sites
C0079774|T191|HT|202.7|ICD9CM|Peripheral T-cell lymphoma|Peripheral T-cell lymphoma
C1955728|T191|AB|202.70|ICD9CM|Periph T cell lym xtrndl|Periph T cell lym xtrndl
C1955728|T191|PT|202.70|ICD9CM|Peripheral T cell lymphoma, unspecified site, extranodal and solid organ sites|Peripheral T cell lymphoma, unspecified site, extranodal and solid organ sites
C3648017|T191|AB|202.71|ICD9CM|Periph T cell lymph head|Periph T cell lymph head
C3648017|T191|PT|202.71|ICD9CM|Peripheral T cell lymphoma, lymph nodes of head, face, and neck|Peripheral T cell lymphoma, lymph nodes of head, face, and neck
C1955730|T191|AB|202.72|ICD9CM|Periph T cell lym thorax|Periph T cell lym thorax
C1955730|T191|PT|202.72|ICD9CM|Peripheral T cell lymphoma, intrathoracic lymph nodes|Peripheral T cell lymphoma, intrathoracic lymph nodes
C3648015|T191|AB|202.73|ICD9CM|Periph T cell lym abdom|Periph T cell lym abdom
C3648015|T191|PT|202.73|ICD9CM|Peripheral T cell lymphoma, intra-abdominal lymph nodes|Peripheral T cell lymphoma, intra-abdominal lymph nodes
C3648018|T191|AB|202.74|ICD9CM|Periph T cell lym axilla|Periph T cell lym axilla
C3648018|T191|PT|202.74|ICD9CM|Peripheral T cell lymphoma, lymph nodes of axilla and upper limb|Peripheral T cell lymphoma, lymph nodes of axilla and upper limb
C3648016|T191|AB|202.75|ICD9CM|Periph T cell lym inguin|Periph T cell lym inguin
C3648016|T191|PT|202.75|ICD9CM|Peripheral T cell lymphoma, lymph nodes of inguinal region and lower limb|Peripheral T cell lymphoma, lymph nodes of inguinal region and lower limb
C3648014|T191|AB|202.76|ICD9CM|Periph T cell lym pelvic|Periph T cell lym pelvic
C3648014|T191|PT|202.76|ICD9CM|Peripheral T cell lymphoma, intrapelvic lymph nodes|Peripheral T cell lymphoma, intrapelvic lymph nodes
C1955735|T191|AB|202.77|ICD9CM|Periph T cell lym spleen|Periph T cell lym spleen
C1955735|T191|PT|202.77|ICD9CM|Peripheral T cell lymphoma, spleen|Peripheral T cell lymphoma, spleen
C3648012|T191|AB|202.78|ICD9CM|Periph T cell lym multip|Periph T cell lym multip
C3648012|T191|PT|202.78|ICD9CM|Peripheral T cell lymphoma, lymph nodes of multiple sites|Peripheral T cell lymphoma, lymph nodes of multiple sites
C0029662|T191|HT|202.8|ICD9CM|Other malignant lymphomas|Other malignant lymphomas
C0375094|T191|AB|202.80|ICD9CM|Oth lymp unsp xtrndl org|Oth lymp unsp xtrndl org
C0375094|T191|PT|202.80|ICD9CM|Other malignant lymphomas, unspecified site, extranodal and solid organ sites|Other malignant lymphomas, unspecified site, extranodal and solid organ sites
C0153850|T191|AB|202.81|ICD9CM|Lymphomas NEC head|Lymphomas NEC head
C0153850|T191|PT|202.81|ICD9CM|Other malignant lymphomas, lymph nodes of head, face, and neck|Other malignant lymphomas, lymph nodes of head, face, and neck
C0153851|T191|AB|202.82|ICD9CM|Lymphomas NEC thorax|Lymphomas NEC thorax
C0153851|T191|PT|202.82|ICD9CM|Other malignant lymphomas, intrathoracic lymph nodes|Other malignant lymphomas, intrathoracic lymph nodes
C0153852|T191|AB|202.83|ICD9CM|Lymphomas NEC abdom|Lymphomas NEC abdom
C0153852|T191|PT|202.83|ICD9CM|Other malignant lymphomas, intra-abdominal lymph nodes|Other malignant lymphomas, intra-abdominal lymph nodes
C0153853|T191|AB|202.84|ICD9CM|Lymphomas NEC axilla|Lymphomas NEC axilla
C0153853|T191|PT|202.84|ICD9CM|Other malignant lymphomas, lymph nodes of axilla and upper limb|Other malignant lymphomas, lymph nodes of axilla and upper limb
C0153854|T191|AB|202.85|ICD9CM|Lymphomas NEC inguin|Lymphomas NEC inguin
C0153854|T191|PT|202.85|ICD9CM|Other malignant lymphomas, lymph nodes of inguinal region and lower limb|Other malignant lymphomas, lymph nodes of inguinal region and lower limb
C0153855|T191|AB|202.86|ICD9CM|Lymphomas NEC pelvic|Lymphomas NEC pelvic
C0153855|T191|PT|202.86|ICD9CM|Other malignant lymphomas, intrapelvic lymph nodes|Other malignant lymphomas, intrapelvic lymph nodes
C0153856|T191|AB|202.87|ICD9CM|Lymphomas NEC spleen|Lymphomas NEC spleen
C0153856|T191|PT|202.87|ICD9CM|Other malignant lymphomas, spleen|Other malignant lymphomas, spleen
C0728903|T191|AB|202.88|ICD9CM|Lymphomas NEC mult|Lymphomas NEC mult
C0728903|T191|PT|202.88|ICD9CM|Other malignant lymphomas, lymph nodes of multiple sites|Other malignant lymphomas, lymph nodes of multiple sites
C0153858|T191|HT|202.9|ICD9CM|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue
C0375095|T191|AB|202.90|ICD9CM|Unsp lym unsp xtrndl org|Unsp lym unsp xtrndl org
C0153859|T191|AB|202.91|ICD9CM|Lymphoid mal NEC head|Lymphoid mal NEC head
C0153860|T191|AB|202.92|ICD9CM|Lymphoid mal NEC thorax|Lymphoid mal NEC thorax
C0153861|T191|AB|202.93|ICD9CM|Lymphoid mal NEC abdom|Lymphoid mal NEC abdom
C0153862|T191|AB|202.94|ICD9CM|Lymphoid mal NEC axilla|Lymphoid mal NEC axilla
C0153863|T191|AB|202.95|ICD9CM|Lymphoid mal NEC inguin|Lymphoid mal NEC inguin
C0153864|T191|AB|202.96|ICD9CM|Lymphoid mal NEC pelvic|Lymphoid mal NEC pelvic
C0153865|T191|AB|202.97|ICD9CM|Lymphoid mal NEC spleen|Lymphoid mal NEC spleen
C0153865|T191|PT|202.97|ICD9CM|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue, spleen|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue, spleen
C0153866|T191|AB|202.98|ICD9CM|Lymphoid mal NEC mult|Lymphoid mal NEC mult
C0153867|T191|HT|203|ICD9CM|Multiple myeloma and immunoproliferative neoplasms|Multiple myeloma and immunoproliferative neoplasms
C0026764|T191|HT|203.0|ICD9CM|Multiple myeloma|Multiple myeloma
C2349260|T191|AB|203.00|ICD9CM|Mult mye w/o achv rmson|Mult mye w/o achv rmson
C2349260|T191|PT|203.00|ICD9CM|Multiple myeloma, without mention of having achieved remission|Multiple myeloma, without mention of having achieved remission
C0153869|T191|AB|203.01|ICD9CM|Mult myelm w remission|Mult myelm w remission
C0153869|T191|PT|203.01|ICD9CM|Multiple myeloma, in remission|Multiple myeloma, in remission
C2349261|T191|AB|203.02|ICD9CM|Mult myeloma in relapse|Mult myeloma in relapse
C2349261|T191|PT|203.02|ICD9CM|Multiple myeloma, in relapse|Multiple myeloma, in relapse
C0023484|T191|HT|203.1|ICD9CM|Plasma cell leukemia|Plasma cell leukemia
C2349262|T191|PT|203.10|ICD9CM|Plasma cell leukemia, without mention of having achieved remission|Plasma cell leukemia, without mention of having achieved remission
C2349262|T191|AB|203.10|ICD9CM|Pls cl leu w/o achv rmsn|Pls cl leu w/o achv rmsn
C0153871|T191|PT|203.11|ICD9CM|Plasma cell leukemia, in remission|Plasma cell leukemia, in remission
C0153871|T191|AB|203.11|ICD9CM|Plsm cell leuk w rmson|Plsm cell leuk w rmson
C2349263|T191|PT|203.12|ICD9CM|Plasma cell leukemia, in relapse|Plasma cell leukemia, in relapse
C2349263|T191|AB|203.12|ICD9CM|Plsm cel leuk in relapse|Plsm cel leuk in relapse
C0153872|T191|HT|203.8|ICD9CM|Other immunoproliferative neoplasms|Other immunoproliferative neoplasms
C2349264|T191|AB|203.80|ICD9CM|Oth imno npl wo ach rmsn|Oth imno npl wo ach rmsn
C2349264|T191|PT|203.80|ICD9CM|Other immunoproliferative neoplasms, without mention of having achieved remission|Other immunoproliferative neoplasms, without mention of having achieved remission
C0153874|T191|AB|203.81|ICD9CM|Oth imnprfl npl w rmsn|Oth imnprfl npl w rmsn
C0153874|T191|PT|203.81|ICD9CM|Other immunoproliferative neoplasms, in remission|Other immunoproliferative neoplasms, in remission
C2349265|T191|AB|203.82|ICD9CM|Oth imnprlf neo-relapse|Oth imnprlf neo-relapse
C2349265|T191|PT|203.82|ICD9CM|Other immunoproliferative neoplasms, in relapse|Other immunoproliferative neoplasms, in relapse
C0023448|T191|HT|204|ICD9CM|Lymphoid leukemia|Lymphoid leukemia
C0023449|T191|HT|204.0|ICD9CM|Lymphoid leukemia, acute|Lymphoid leukemia, acute
C2349266|T191|AB|204.00|ICD9CM|Ac lym leuk wo achv rmsn|Ac lym leuk wo achv rmsn
C2349266|T191|PT|204.00|ICD9CM|Acute lymphoid leukemia, without mention of having achieved remission|Acute lymphoid leukemia, without mention of having achieved remission
C0153876|T191|AB|204.01|ICD9CM|Act lym leuk w rmsion|Act lym leuk w rmsion
C0153876|T191|PT|204.01|ICD9CM|Acute lymphoid leukemia, in remission|Acute lymphoid leukemia, in remission
C2349267|T191|AB|204.02|ICD9CM|Act lymp leuk in relapse|Act lymp leuk in relapse
C2349267|T191|PT|204.02|ICD9CM|Acute lymphoid leukemia, in relapse|Acute lymphoid leukemia, in relapse
C0023434|T191|HT|204.1|ICD9CM|Lymphoid leukemia, chronic|Lymphoid leukemia, chronic
C2349268|T191|AB|204.10|ICD9CM|Ch lym leuk wo achv rmsn|Ch lym leuk wo achv rmsn
C2349268|T191|PT|204.10|ICD9CM|Chronic lymphoid leukemia, without mention of having achieved remission|Chronic lymphoid leukemia, without mention of having achieved remission
C0153878|T191|AB|204.11|ICD9CM|Chr lym leuk w rmsion|Chr lym leuk w rmsion
C0153878|T191|PT|204.11|ICD9CM|Chronic lymphoid leukemia, in remission|Chronic lymphoid leukemia, in remission
C0854802|T191|AB|204.12|ICD9CM|Chr lymp leuk in relapse|Chr lymp leuk in relapse
C0854802|T191|PT|204.12|ICD9CM|Chronic lymphoid leukemia, in relapse|Chronic lymphoid leukemia, in relapse
C0152271|T191|HT|204.2|ICD9CM|Lymphoid leukemia, subacute|Lymphoid leukemia, subacute
C2349269|T191|AB|204.20|ICD9CM|Sbac lym leu wo ach rmsn|Sbac lym leu wo ach rmsn
C2349269|T191|PT|204.20|ICD9CM|Subacute lymphoid leukemia, without mention of having achieved remission|Subacute lymphoid leukemia, without mention of having achieved remission
C0153880|T191|AB|204.21|ICD9CM|Sbac lym leuk w rmsion|Sbac lym leuk w rmsion
C0153880|T191|PT|204.21|ICD9CM|Subacute lymphoid leukemia, in remission|Subacute lymphoid leukemia, in remission
C2349270|T191|AB|204.22|ICD9CM|Sbac lym leuk in relapse|Sbac lym leuk in relapse
C2349270|T191|PT|204.22|ICD9CM|Subacute lymphoid leukemia, in relapse|Subacute lymphoid leukemia, in relapse
C0029660|T191|HT|204.8|ICD9CM|Other lymphoid leukemia|Other lymphoid leukemia
C2349271|T191|AB|204.80|ICD9CM|Oth lym leu wo achv rmsn|Oth lym leu wo achv rmsn
C2349271|T191|PT|204.80|ICD9CM|Other lymphoid leukemia, without mention of having achieved remission|Other lymphoid leukemia, without mention of having achieved remission
C0153882|T191|AB|204.81|ICD9CM|Oth lym leuk w rmsion|Oth lym leuk w rmsion
C0153882|T191|PT|204.81|ICD9CM|Other lymphoid leukemia, in remission|Other lymphoid leukemia, in remission
C2349272|T191|AB|204.82|ICD9CM|Oth lym leuk in relapse|Oth lym leuk in relapse
C2349272|T191|PT|204.82|ICD9CM|Other lymphoid leukemia, in relapse|Other lymphoid leukemia, in relapse
C0023448|T191|HT|204.9|ICD9CM|Unspecified lymphoid leukemia|Unspecified lymphoid leukemia
C2349273|T191|AB|204.90|ICD9CM|Uns lym leu wo ach rmsn|Uns lym leu wo ach rmsn
C2349273|T191|PT|204.90|ICD9CM|Unspecified lymphoid leukemia, without mention of having achieved remission|Unspecified lymphoid leukemia, without mention of having achieved remission
C0686597|T191|AB|204.91|ICD9CM|Uns lym leuk w rmsion|Uns lym leuk w rmsion
C0686597|T191|PT|204.91|ICD9CM|Unspecified lymphoid leukemia, in remission|Unspecified lymphoid leukemia, in remission
C2349274|T191|AB|204.92|ICD9CM|Lymp leuk NOS relapse|Lymp leuk NOS relapse
C2349274|T191|PT|204.92|ICD9CM|Unspecified lymphoid leukemia, in relapse|Unspecified lymphoid leukemia, in relapse
C0023470|T191|HT|205|ICD9CM|Myeloid leukemia|Myeloid leukemia
C0023467|T191|HT|205.0|ICD9CM|Myeloid leukemia, acute|Myeloid leukemia, acute
C2349275|T191|AB|205.00|ICD9CM|Ac myl leuk wo achv rmsn|Ac myl leuk wo achv rmsn
C2349275|T191|PT|205.00|ICD9CM|Acute myeloid leukemia, without mention of having achieved remission|Acute myeloid leukemia, without mention of having achieved remission
C0153886|T191|AB|205.01|ICD9CM|Act myl leuk w rmsion|Act myl leuk w rmsion
C0153886|T191|PT|205.01|ICD9CM|Acute myeloid leukemia, in remission|Acute myeloid leukemia, in remission
C2349276|T191|AB|205.02|ICD9CM|Act myel leuk in relapse|Act myel leuk in relapse
C2349276|T191|PT|205.02|ICD9CM|Acute myeloid leukemia, in relapse|Acute myeloid leukemia, in relapse
C0023473|T191|HT|205.1|ICD9CM|Myeloid leukemia, chronic|Myeloid leukemia, chronic
C2349277|T191|AB|205.10|ICD9CM|Ch myl leuk wo achv rmsn|Ch myl leuk wo achv rmsn
C2349277|T191|PT|205.10|ICD9CM|Chronic myeloid leukemia, without mention of having achieved remission|Chronic myeloid leukemia, without mention of having achieved remission
C0153888|T191|AB|205.11|ICD9CM|Chr myl leuk w rmsion|Chr myl leuk w rmsion
C0153888|T191|PT|205.11|ICD9CM|Chronic myeloid leukemia, in remission|Chronic myeloid leukemia, in remission
C1532368|T191|AB|205.12|ICD9CM|Chr myel leuk in relapse|Chr myel leuk in relapse
C1532368|T191|PT|205.12|ICD9CM|Chronic myeloid leukemia, in relapse|Chronic myeloid leukemia, in relapse
C1292772|T191|HT|205.2|ICD9CM|Myeloid leukemia, subacute|Myeloid leukemia, subacute
C2349278|T191|AB|205.20|ICD9CM|Sbac myl leu wo ach rmsn|Sbac myl leu wo ach rmsn
C2349278|T191|PT|205.20|ICD9CM|Subacute myeloid leukemia, without mention of having achieved remission|Subacute myeloid leukemia, without mention of having achieved remission
C0153890|T191|AB|205.21|ICD9CM|Sbac myl leuk w rmsion|Sbac myl leuk w rmsion
C0153890|T191|PT|205.21|ICD9CM|Subacute myeloid leukemia,in remission|Subacute myeloid leukemia,in remission
C2349279|T191|AB|205.22|ICD9CM|Sbac myl leuk in relapse|Sbac myl leuk in relapse
C2349279|T191|PT|205.22|ICD9CM|Subacute myeloid leukemia, in relapse|Subacute myeloid leukemia, in relapse
C4721505|T191|HT|205.3|ICD9CM|Myeloid sarcoma|Myeloid sarcoma
C2349280|T191|PT|205.30|ICD9CM|Myeloid sarcoma, without mention of having achieved remission|Myeloid sarcoma, without mention of having achieved remission
C2349280|T191|AB|205.30|ICD9CM|Myl sarcoma wo achv rmsn|Myl sarcoma wo achv rmsn
C0153892|T191|PT|205.31|ICD9CM|Myeloid sarcoma, in remission|Myeloid sarcoma, in remission
C0153892|T191|AB|205.31|ICD9CM|Myl srcoma w rmsion|Myl srcoma w rmsion
C2349281|T191|AB|205.32|ICD9CM|Myel sarcoma in relapse|Myel sarcoma in relapse
C2349281|T191|PT|205.32|ICD9CM|Myeloid sarcoma, in relapse|Myeloid sarcoma, in relapse
C0029670|T191|HT|205.8|ICD9CM|Other myeloid leukemia|Other myeloid leukemia
C2349282|T191|AB|205.80|ICD9CM|Oth my leuk wo achv rmsn|Oth my leuk wo achv rmsn
C2349282|T191|PT|205.80|ICD9CM|Other myeloid leukemia, without mention of having achieved remission|Other myeloid leukemia, without mention of having achieved remission
C0153894|T191|AB|205.81|ICD9CM|Oth myl leuk w rmsion|Oth myl leuk w rmsion
C0153894|T191|PT|205.81|ICD9CM|Other myeloid leukemia, in remission|Other myeloid leukemia, in remission
C2349283|T191|AB|205.82|ICD9CM|Oth myel leuk in relapse|Oth myel leuk in relapse
C2349283|T191|PT|205.82|ICD9CM|Other myeloid leukemia, in relapse|Other myeloid leukemia, in relapse
C0023470|T191|HT|205.9|ICD9CM|Unspecified myeloid leukemia|Unspecified myeloid leukemia
C2349284|T191|AB|205.90|ICD9CM|Uns my leu wo ach rmsn|Uns my leu wo ach rmsn
C2349284|T191|PT|205.90|ICD9CM|Unspecified myeloid leukemia, without mention of having achieved remission|Unspecified myeloid leukemia, without mention of having achieved remission
C0686593|T191|AB|205.91|ICD9CM|Uns myl leuk w rmsion|Uns myl leuk w rmsion
C0686593|T191|PT|205.91|ICD9CM|Unspecified myeloid leukemia, in remission|Unspecified myeloid leukemia, in remission
C2349285|T191|AB|205.92|ICD9CM|Myel leuk NOS in relapse|Myel leuk NOS in relapse
C2349285|T191|PT|205.92|ICD9CM|Unspecified myeloid leukemia, in relapse|Unspecified myeloid leukemia, in relapse
C0598894|T191|HT|206|ICD9CM|Monocytic leukemia|Monocytic leukemia
C0023465|T191|HT|206.0|ICD9CM|Monocytic leukemia, acute|Monocytic leukemia, acute
C2349286|T191|AB|206.00|ICD9CM|Ac mono leu wo achv rmsn|Ac mono leu wo achv rmsn
C2349286|T191|PT|206.00|ICD9CM|Acute monocytic leukemia, without mention of having achieved remission|Acute monocytic leukemia, without mention of having achieved remission
C0153898|T191|AB|206.01|ICD9CM|Act mono leuk w rmsion|Act mono leuk w rmsion
C0153898|T191|PT|206.01|ICD9CM|Acute monocytic leukemia,in remission|Acute monocytic leukemia,in remission
C2349287|T191|AB|206.02|ICD9CM|Act mono leuk in relapse|Act mono leuk in relapse
C2349287|T191|PT|206.02|ICD9CM|Acute monocytic leukemia, in relapse|Acute monocytic leukemia, in relapse
C0023466|T191|HT|206.1|ICD9CM|Monocytic leukemia, chronic|Monocytic leukemia, chronic
C2349288|T191|AB|206.10|ICD9CM|Ch mono leu wo achv rmsn|Ch mono leu wo achv rmsn
C2349288|T191|PT|206.10|ICD9CM|Chronic monocytic leukemia, without mention of having achieved remission|Chronic monocytic leukemia, without mention of having achieved remission
C0153900|T191|AB|206.11|ICD9CM|Chr mono leuk w rmsion|Chr mono leuk w rmsion
C0153900|T191|PT|206.11|ICD9CM|Chronic monocytic leukemia, in remission|Chronic monocytic leukemia, in remission
C2349289|T191|AB|206.12|ICD9CM|Chr mono leuk in relapse|Chr mono leuk in relapse
C2349289|T191|PT|206.12|ICD9CM|Chronic monocytic leukemia, in relapse|Chronic monocytic leukemia, in relapse
C0152275|T191|HT|206.2|ICD9CM|Monocytic leukemia, subacute|Monocytic leukemia, subacute
C2349290|T191|AB|206.20|ICD9CM|Sbac mno leu wo ach rmsn|Sbac mno leu wo ach rmsn
C2349290|T191|PT|206.20|ICD9CM|Subacute monocytic leukemia, without mention of having achieved remission|Subacute monocytic leukemia, without mention of having achieved remission
C0153902|T191|AB|206.21|ICD9CM|Sbac mono leuk w rmsion|Sbac mono leuk w rmsion
C0153902|T191|PT|206.21|ICD9CM|Subacute monocytic leukemia, in remission|Subacute monocytic leukemia, in remission
C2349291|T191|AB|206.22|ICD9CM|Sbac mono leu in relapse|Sbac mono leu in relapse
C2349291|T191|PT|206.22|ICD9CM|Subacute monocytic leukemia, in relapse|Subacute monocytic leukemia, in relapse
C0153903|T191|HT|206.8|ICD9CM|Other monocytic leukemia|Other monocytic leukemia
C2349292|T191|AB|206.80|ICD9CM|Ot mono leu wo achv rmsn|Ot mono leu wo achv rmsn
C2349292|T191|PT|206.80|ICD9CM|Other monocytic leukemia, without mention of having achieved remission|Other monocytic leukemia, without mention of having achieved remission
C0153905|T191|AB|206.81|ICD9CM|Oth mono leuk w rmsion|Oth mono leuk w rmsion
C0153905|T191|PT|206.81|ICD9CM|Other monocytic leukemia, in remission|Other monocytic leukemia, in remission
C2349293|T191|AB|206.82|ICD9CM|Oth mono leuk in relapse|Oth mono leuk in relapse
C2349293|T191|PT|206.82|ICD9CM|Other monocytic leukemia, in relapse|Other monocytic leukemia, in relapse
C0598894|T191|HT|206.9|ICD9CM|Unspecified monocytic leukemia|Unspecified monocytic leukemia
C2349294|T191|AB|206.90|ICD9CM|Uns mno leu wo ach rmsn|Uns mno leu wo ach rmsn
C2349294|T191|PT|206.90|ICD9CM|Unspecified monocytic leukemia, without mention of having achieved remission|Unspecified monocytic leukemia, without mention of having achieved remission
C0686595|T191|AB|206.91|ICD9CM|Uns mono leuk w rmsion|Uns mono leuk w rmsion
C0686595|T191|PT|206.91|ICD9CM|Unspecified monocytic leukemia, in remission|Unspecified monocytic leukemia, in remission
C2349295|T191|AB|206.92|ICD9CM|Mono leuk NOS relapse|Mono leuk NOS relapse
C2349295|T191|PT|206.92|ICD9CM|Unspecified monocytic leukemia, in relapse|Unspecified monocytic leukemia, in relapse
C0029812|T191|HT|207|ICD9CM|Other specified leukemia|Other specified leukemia
C0001317|T191|HT|207.0|ICD9CM|Acute erythremia and erythroleukemia|Acute erythremia and erythroleukemia
C2349296|T191|AB|207.00|ICD9CM|Ac erth/erlk wo ach rmsn|Ac erth/erlk wo ach rmsn
C2349296|T191|PT|207.00|ICD9CM|Acute erythremia and erythroleukemia, without mention of having achieved remission|Acute erythremia and erythroleukemia, without mention of having achieved remission
C0153910|T191|AB|207.01|ICD9CM|Act erth/erylk w rmson|Act erth/erylk w rmson
C0153910|T191|PT|207.01|ICD9CM|Acute erythremia and erythroleukemia, in remission|Acute erythremia and erythroleukemia, in remission
C2349297|T191|AB|207.02|ICD9CM|Ac erth/erylk in relapse|Ac erth/erylk in relapse
C2349297|T191|PT|207.02|ICD9CM|Acute erythremia and erythroleukemia, in relapse|Acute erythremia and erythroleukemia, in relapse
C0152272|T191|HT|207.1|ICD9CM|Chronic erythremia|Chronic erythremia
C2349298|T191|AB|207.10|ICD9CM|Chr erythrm w/o ach rmsn|Chr erythrm w/o ach rmsn
C2349298|T191|PT|207.10|ICD9CM|Chronic erythremia, without mention of having achieved remission|Chronic erythremia, without mention of having achieved remission
C0153912|T191|AB|207.11|ICD9CM|Chr erythrm w remision|Chr erythrm w remision
C0153912|T191|PT|207.11|ICD9CM|Chronic erythremia, in remission|Chronic erythremia, in remission
C2349299|T191|AB|207.12|ICD9CM|Chr erythrmia in relapse|Chr erythrmia in relapse
C2349299|T191|PT|207.12|ICD9CM|Chronic erythremia, in relapse|Chronic erythremia, in relapse
C0023462|T191|HT|207.2|ICD9CM|Megakaryocytic leukemia|Megakaryocytic leukemia
C2349300|T191|PT|207.20|ICD9CM|Megakaryocytic leukemia, without mention of having achieved remission|Megakaryocytic leukemia, without mention of having achieved remission
C2349300|T191|AB|207.20|ICD9CM|Mgkrcyt leuk wo ach rmsn|Mgkrcyt leuk wo ach rmsn
C0153914|T191|PT|207.21|ICD9CM|Megakaryocytic leukemia, in remission|Megakaryocytic leukemia, in remission
C0153914|T191|AB|207.21|ICD9CM|Mgkrycyt leuk w rmsion|Mgkrycyt leuk w rmsion
C2349301|T191|PT|207.22|ICD9CM|Megakaryocytic leukemia, in relapse|Megakaryocytic leukemia, in relapse
C2349301|T191|AB|207.22|ICD9CM|Mgkrycyt leuk in relapse|Mgkrycyt leuk in relapse
C0029812|T191|HT|207.8|ICD9CM|Other specified leukemia|Other specified leukemia
C2349302|T191|AB|207.80|ICD9CM|Oth leuk w/o achv rmsn|Oth leuk w/o achv rmsn
C2349302|T191|PT|207.80|ICD9CM|Other specified leukemia, without mention of having achieved remission|Other specified leukemia, without mention of having achieved remission
C0153916|T191|AB|207.81|ICD9CM|Oth spf leuk w remsion|Oth spf leuk w remsion
C0153916|T191|PT|207.81|ICD9CM|Other specified leukemia, in remission|Other specified leukemia, in remission
C2349303|T191|AB|207.82|ICD9CM|Oth spf leuk in relapse|Oth spf leuk in relapse
C2349303|T191|PT|207.82|ICD9CM|Other specified leukemia, in relapse|Other specified leukemia, in relapse
C0023418|T191|HT|208|ICD9CM|Leukemia of unspecified cell type|Leukemia of unspecified cell type
C0085669|T191|HT|208.0|ICD9CM|Leukemia of unspecified cell type, acute|Leukemia of unspecified cell type, acute
C2349304|T191|AB|208.00|ICD9CM|Ac leu un cl wo ach rmsn|Ac leu un cl wo ach rmsn
C2349304|T191|PT|208.00|ICD9CM|Acute leukemia of unspecified cell type, without mention of having achieved remission|Acute leukemia of unspecified cell type, without mention of having achieved remission
C0686586|T191|AB|208.01|ICD9CM|Act leuk uns cl w rmson|Act leuk uns cl w rmson
C0686586|T191|PT|208.01|ICD9CM|Acute leukemia of unspecified cell type, in remission|Acute leukemia of unspecified cell type, in remission
C2349305|T191|AB|208.02|ICD9CM|Ac leuk uns cl relapse|Ac leuk uns cl relapse
C2349305|T191|PT|208.02|ICD9CM|Acute leukemia of unspecified cell type, in relapse|Acute leukemia of unspecified cell type, in relapse
C1279296|T191|HT|208.1|ICD9CM|Leukemia of unspecified cell type, chronic|Leukemia of unspecified cell type, chronic
C2349306|T191|AB|208.10|ICD9CM|Ch leu un cl wo ach rmsn|Ch leu un cl wo ach rmsn
C2349306|T191|PT|208.10|ICD9CM|Chronic leukemia of unspecified cell type, without mention of having achieved remission|Chronic leukemia of unspecified cell type, without mention of having achieved remission
C0686589|T191|AB|208.11|ICD9CM|Chr leuk uns cl w rmson|Chr leuk uns cl w rmson
C0686589|T191|PT|208.11|ICD9CM|Chronic leukemia of unspecified cell type, in remission|Chronic leukemia of unspecified cell type, in remission
C2349307|T191|AB|208.12|ICD9CM|Ch leu uns cl in relapse|Ch leu uns cl in relapse
C2349307|T191|PT|208.12|ICD9CM|Chronic leukemia of unspecified cell type, in relapse|Chronic leukemia of unspecified cell type, in relapse
C0153924|T191|HT|208.2|ICD9CM|Leukemia of unspecified cell type, subacute|Leukemia of unspecified cell type, subacute
C2349308|T191|AB|208.20|ICD9CM|Sbc leu un cl wo ah rmsn|Sbc leu un cl wo ah rmsn
C2349308|T191|PT|208.20|ICD9CM|Subacute leukemia of unspecified cell type, without mention of having achieved remission|Subacute leukemia of unspecified cell type, without mention of having achieved remission
C0686591|T191|AB|208.21|ICD9CM|Sbac leuk uns cl w rmson|Sbac leuk uns cl w rmson
C0686591|T191|PT|208.21|ICD9CM|Subacute leukemia of unspecified cell type, in remission|Subacute leukemia of unspecified cell type, in remission
C2349309|T191|AB|208.22|ICD9CM|Sbac leu uns cl-relapse|Sbac leu uns cl-relapse
C2349309|T191|PT|208.22|ICD9CM|Subacute leukemia of unspecified cell type, in relapse|Subacute leukemia of unspecified cell type, in relapse
C0029655|T191|HT|208.8|ICD9CM|Other leukemia of unspecified cell type|Other leukemia of unspecified cell type
C2349310|T191|AB|208.80|ICD9CM|Ot leu un cl wo ach rmsn|Ot leu un cl wo ach rmsn
C2349310|T191|PT|208.80|ICD9CM|Other leukemia of unspecified cell type, without mention of having achieved remission|Other leukemia of unspecified cell type, without mention of having achieved remission
C0153928|T191|AB|208.81|ICD9CM|Oth leuk uns cl w rmson|Oth leuk uns cl w rmson
C0153928|T191|PT|208.81|ICD9CM|Other leukemia of unspecified cell type, in remission|Other leukemia of unspecified cell type, in remission
C2349311|T191|AB|208.82|ICD9CM|Oth leuk uns cl-relapse|Oth leuk uns cl-relapse
C2349311|T191|PT|208.82|ICD9CM|Other leukemia of unspecified cell type, in relapse|Other leukemia of unspecified cell type, in relapse
C0023418|T191|HT|208.9|ICD9CM|Unspecified leukemia|Unspecified leukemia
C2349312|T191|AB|208.90|ICD9CM|Leuk NOS w/o achv rmsn|Leuk NOS w/o achv rmsn
C2349312|T191|PT|208.90|ICD9CM|Unspecified leukemia, without mention of having achieved remission|Unspecified leukemia, without mention of having achieved remission
C0686584|T191|AB|208.91|ICD9CM|Leukemia NOS w remission|Leukemia NOS w remission
C0686584|T191|PT|208.91|ICD9CM|Unspecified leukemia, in remission|Unspecified leukemia, in remission
C0920028|T191|AB|208.92|ICD9CM|Leukemia NOS in relapse|Leukemia NOS in relapse
C0920028|T191|PT|208.92|ICD9CM|Unspecified leukemia, in relapse|Unspecified leukemia, in relapse
C0206754|T191|HT|209|ICD9CM|Neuroendocrine tumors|Neuroendocrine tumors
C0206754|T191|HT|209-209.99|ICD9CM|NEUROENDOCRINE TUMORS|NEUROENDOCRINE TUMORS
C2062527|T191|HT|209.0|ICD9CM|Malignant carcinoid tumors of the small intestine|Malignant carcinoid tumors of the small intestine
C2349313|T191|AB|209.00|ICD9CM|Mal crcnoid sm intst NOS|Mal crcnoid sm intst NOS
C2349313|T191|PT|209.00|ICD9CM|Malignant carcinoid tumor of the small intestine, unspecified portion|Malignant carcinoid tumor of the small intestine, unspecified portion
C2349314|T191|AB|209.01|ICD9CM|Malig carcinoid duodenum|Malig carcinoid duodenum
C2349314|T191|PT|209.01|ICD9CM|Malignant carcinoid tumor of the duodenum|Malignant carcinoid tumor of the duodenum
C2349315|T191|AB|209.02|ICD9CM|Malig carcinoid jejunum|Malig carcinoid jejunum
C2349315|T191|PT|209.02|ICD9CM|Malignant carcinoid tumor of the jejunum|Malignant carcinoid tumor of the jejunum
C2349316|T191|AB|209.03|ICD9CM|Malig carcinoid ileum|Malig carcinoid ileum
C2349316|T191|PT|209.03|ICD9CM|Malignant carcinoid tumor of the ileum|Malignant carcinoid tumor of the ileum
C2349324|T191|HT|209.1|ICD9CM|Malignant carcinoid tumors of the appendix, large intestine, and rectum|Malignant carcinoid tumors of the appendix, large intestine, and rectum
C2349317|T191|AB|209.10|ICD9CM|Mal crcnoid lg intst NOS|Mal crcnoid lg intst NOS
C2349317|T191|PT|209.10|ICD9CM|Malignant carcinoid tumor of the large intestine, unspecified portion|Malignant carcinoid tumor of the large intestine, unspecified portion
C2062529|T191|AB|209.11|ICD9CM|Malig carcinoid appendix|Malig carcinoid appendix
C2062529|T191|PT|209.11|ICD9CM|Malignant carcinoid tumor of the appendix|Malignant carcinoid tumor of the appendix
C2349319|T191|AB|209.12|ICD9CM|Malig carcinoid cecum|Malig carcinoid cecum
C2349319|T191|PT|209.12|ICD9CM|Malignant carcinoid tumor of the cecum|Malignant carcinoid tumor of the cecum
C2349320|T191|AB|209.13|ICD9CM|Mal crcnoid ascend colon|Mal crcnoid ascend colon
C2349320|T191|PT|209.13|ICD9CM|Malignant carcinoid tumor of the ascending colon|Malignant carcinoid tumor of the ascending colon
C2349321|T191|AB|209.14|ICD9CM|Mal crcnoid transv colon|Mal crcnoid transv colon
C2349321|T191|PT|209.14|ICD9CM|Malignant carcinoid tumor of the transverse colon|Malignant carcinoid tumor of the transverse colon
C2349322|T191|AB|209.15|ICD9CM|Mal carcinoid desc colon|Mal carcinoid desc colon
C2349322|T191|PT|209.15|ICD9CM|Malignant carcinoid tumor of the descending colon|Malignant carcinoid tumor of the descending colon
C2349323|T191|AB|209.16|ICD9CM|Mal carcinoid sig colon|Mal carcinoid sig colon
C2349323|T191|PT|209.16|ICD9CM|Malignant carcinoid tumor of the sigmoid colon|Malignant carcinoid tumor of the sigmoid colon
C2205119|T191|AB|209.17|ICD9CM|Malig carcinoid rectum|Malig carcinoid rectum
C2205119|T191|PT|209.17|ICD9CM|Malignant carcinoid tumor of the rectum|Malignant carcinoid tumor of the rectum
C2349332|T191|HT|209.2|ICD9CM|Malignant carcinoid tumors of other and unspecified sites|Malignant carcinoid tumors of other and unspecified sites
C2349325|T191|AB|209.20|ICD9CM|Mal crcnd prim site unkn|Mal crcnd prim site unkn
C2349325|T191|PT|209.20|ICD9CM|Malignant carcinoid tumor of unknown primary site|Malignant carcinoid tumor of unknown primary site
C2349326|T191|AB|209.21|ICD9CM|Mal carcinoid bronc/lung|Mal carcinoid bronc/lung
C2349326|T191|PT|209.21|ICD9CM|Malignant carcinoid tumor of the bronchus and lung|Malignant carcinoid tumor of the bronchus and lung
C1336746|T191|AB|209.22|ICD9CM|Malig carcinoid thymus|Malig carcinoid thymus
C1336746|T191|PT|209.22|ICD9CM|Malignant carcinoid tumor of the thymus|Malignant carcinoid tumor of the thymus
C2062573|T191|AB|209.23|ICD9CM|Malig carcinoid stomach|Malig carcinoid stomach
C2062573|T191|PT|209.23|ICD9CM|Malignant carcinoid tumor of the stomach|Malignant carcinoid tumor of the stomach
C2349327|T191|AB|209.24|ICD9CM|Malig carcinoid kidney|Malig carcinoid kidney
C2349327|T191|PT|209.24|ICD9CM|Malignant carcinoid tumor of the kidney|Malignant carcinoid tumor of the kidney
C2349328|T191|AB|209.25|ICD9CM|Mal carcnoid foregut NOS|Mal carcnoid foregut NOS
C2349328|T191|PT|209.25|ICD9CM|Malignant carcinoid tumor of foregut, not otherwise specified|Malignant carcinoid tumor of foregut, not otherwise specified
C2349329|T191|AB|209.26|ICD9CM|Mal carcinoid midgut NOS|Mal carcinoid midgut NOS
C2349329|T191|PT|209.26|ICD9CM|Malignant carcinoid tumor of midgut, not otherwise specified|Malignant carcinoid tumor of midgut, not otherwise specified
C2349330|T191|AB|209.27|ICD9CM|Mal carcnoid hindgut NOS|Mal carcnoid hindgut NOS
C2349330|T191|PT|209.27|ICD9CM|Malignant carcinoid tumor of hindgut, not otherwise specified|Malignant carcinoid tumor of hindgut, not otherwise specified
C2349331|T191|AB|209.29|ICD9CM|Malig carcinoid oth site|Malig carcinoid oth site
C2349331|T191|PT|209.29|ICD9CM|Malignant carcinoid tumor of other sites|Malignant carcinoid tumor of other sites
C2349335|T191|HT|209.3|ICD9CM|Malignant poorly differentiated neuroendocrine tumors|Malignant poorly differentiated neuroendocrine tumors
C2349333|T191|AB|209.30|ICD9CM|Malig neuroendo ca NOS|Malig neuroendo ca NOS
C2349333|T191|PT|209.30|ICD9CM|Malignant poorly differentiated neuroendocrine carcinoma, any site|Malignant poorly differentiated neuroendocrine carcinoma, any site
C2712672|T191|AB|209.31|ICD9CM|Merkel cell ca-face|Merkel cell ca-face
C2712672|T191|PT|209.31|ICD9CM|Merkel cell carcinoma of the face|Merkel cell carcinoma of the face
C2712692|T191|AB|209.32|ICD9CM|Merkel cell ca-sclp/neck|Merkel cell ca-sclp/neck
C2712692|T191|PT|209.32|ICD9CM|Merkel cell carcinoma of the scalp and neck|Merkel cell carcinoma of the scalp and neck
C4076715|T191|AB|209.33|ICD9CM|Merkel cell ca-up limb|Merkel cell ca-up limb
C4076715|T191|PT|209.33|ICD9CM|Merkel cell carcinoma of the upper limb|Merkel cell carcinoma of the upper limb
C4076723|T191|AB|209.34|ICD9CM|Merkel cell ca-low limb|Merkel cell ca-low limb
C4076723|T191|PT|209.34|ICD9CM|Merkel cell carcinoma of the lower limb|Merkel cell carcinoma of the lower limb
C2712728|T191|AB|209.35|ICD9CM|Merkel cell ca-trunk|Merkel cell ca-trunk
C2712728|T191|PT|209.35|ICD9CM|Merkel cell carcinoma of the trunk|Merkel cell carcinoma of the trunk
C2712734|T191|AB|209.36|ICD9CM|Merkel cell ca-oth sites|Merkel cell ca-oth sites
C2712734|T191|PT|209.36|ICD9CM|Merkel cell carcinoma of other sites|Merkel cell carcinoma of other sites
C2349340|T191|HT|209.4|ICD9CM|Benign carcinoid tumors of the small intestine|Benign carcinoid tumors of the small intestine
C2349336|T191|AB|209.40|ICD9CM|Ben crcnoid sm intst NOS|Ben crcnoid sm intst NOS
C2349336|T191|PT|209.40|ICD9CM|Benign carcinoid tumor of the small intestine, unspecified portion|Benign carcinoid tumor of the small intestine, unspecified portion
C2349337|T191|AB|209.41|ICD9CM|Ben carcinoid duodenum|Ben carcinoid duodenum
C2349337|T191|PT|209.41|ICD9CM|Benign carcinoid tumor of the duodenum|Benign carcinoid tumor of the duodenum
C2349338|T191|AB|209.42|ICD9CM|Benign carcinoid jejunum|Benign carcinoid jejunum
C2349338|T191|PT|209.42|ICD9CM|Benign carcinoid tumor of the jejunum|Benign carcinoid tumor of the jejunum
C2349339|T191|AB|209.43|ICD9CM|Benign carcinoid ileum|Benign carcinoid ileum
C2349339|T191|PT|209.43|ICD9CM|Benign carcinoid tumor of the ileum|Benign carcinoid tumor of the ileum
C2349349|T191|HT|209.5|ICD9CM|Benign carcinoid tumors of the appendix, large intestine, and rectum|Benign carcinoid tumors of the appendix, large intestine, and rectum
C2349341|T191|AB|209.50|ICD9CM|Ben crcnoid lg intst NOS|Ben crcnoid lg intst NOS
C2349341|T191|PT|209.50|ICD9CM|Benign carcinoid tumor of the large intestine, unspecified portion|Benign carcinoid tumor of the large intestine, unspecified portion
C2349342|T191|AB|209.51|ICD9CM|Ben carcinoid appendix|Ben carcinoid appendix
C2349342|T191|PT|209.51|ICD9CM|Benign carcinoid tumor of the appendix|Benign carcinoid tumor of the appendix
C2349343|T191|AB|209.52|ICD9CM|Benign carcinoid cecum|Benign carcinoid cecum
C2349343|T191|PT|209.52|ICD9CM|Benign carcinoid tumor of the cecum|Benign carcinoid tumor of the cecum
C2349344|T191|AB|209.53|ICD9CM|Ben carcinoid asc colon|Ben carcinoid asc colon
C2349344|T191|PT|209.53|ICD9CM|Benign carcinoid tumor of the ascending colon|Benign carcinoid tumor of the ascending colon
C2349345|T191|AB|209.54|ICD9CM|Ben crcinoid trans colon|Ben crcinoid trans colon
C2349345|T191|PT|209.54|ICD9CM|Benign carcinoid tumor of the transverse colon|Benign carcinoid tumor of the transverse colon
C2349346|T191|AB|209.55|ICD9CM|Ben carcinoid desc colon|Ben carcinoid desc colon
C2349346|T191|PT|209.55|ICD9CM|Benign carcinoid tumor of the descending colon|Benign carcinoid tumor of the descending colon
C2349347|T191|AB|209.56|ICD9CM|Ben carcinoid sig colon|Ben carcinoid sig colon
C2349347|T191|PT|209.56|ICD9CM|Benign carcinoid tumor of the sigmoid colon|Benign carcinoid tumor of the sigmoid colon
C2349348|T191|AB|209.57|ICD9CM|Benign carcinoid rectum|Benign carcinoid rectum
C2349348|T191|PT|209.57|ICD9CM|Benign carcinoid tumor of the rectum|Benign carcinoid tumor of the rectum
C2349359|T191|HT|209.6|ICD9CM|Benign carcinoid tumors of other and unspecified sites|Benign carcinoid tumors of other and unspecified sites
C2349350|T191|AB|209.60|ICD9CM|Ben crcnd prim site unkn|Ben crcnd prim site unkn
C2349350|T191|PT|209.60|ICD9CM|Benign carcinoid tumor of unknown primary site|Benign carcinoid tumor of unknown primary site
C2349351|T191|AB|209.61|ICD9CM|Ben carcinoid bronc/lung|Ben carcinoid bronc/lung
C2349351|T191|PT|209.61|ICD9CM|Benign carcinoid tumor of the bronchus and lung|Benign carcinoid tumor of the bronchus and lung
C2349352|T191|AB|209.62|ICD9CM|Benign carcinoid thymus|Benign carcinoid thymus
C2349352|T191|PT|209.62|ICD9CM|Benign carcinoid tumor of the thymus|Benign carcinoid tumor of the thymus
C2349353|T191|AB|209.63|ICD9CM|Benign carcinoid stomach|Benign carcinoid stomach
C2349353|T191|PT|209.63|ICD9CM|Benign carcinoid tumor of the stomach|Benign carcinoid tumor of the stomach
C2349354|T191|AB|209.64|ICD9CM|Benign carcinoid kidney|Benign carcinoid kidney
C2349354|T191|PT|209.64|ICD9CM|Benign carcinoid tumor of the kidney|Benign carcinoid tumor of the kidney
C2349355|T191|AB|209.65|ICD9CM|Ben crcinoid foregut NOS|Ben crcinoid foregut NOS
C2349355|T191|PT|209.65|ICD9CM|Benign carcinoid tumor of foregut, not otherwise specified|Benign carcinoid tumor of foregut, not otherwise specified
C2349356|T191|AB|209.66|ICD9CM|Ben crcinoid midgut NOS|Ben crcinoid midgut NOS
C2349356|T191|PT|209.66|ICD9CM|Benign carcinoid tumor of midgut, not otherwise specified|Benign carcinoid tumor of midgut, not otherwise specified
C2349357|T191|AB|209.67|ICD9CM|Ben crcnoid hindgut NOS|Ben crcnoid hindgut NOS
C2349357|T191|PT|209.67|ICD9CM|Benign carcinoid tumor of hindgut, not otherwise specified|Benign carcinoid tumor of hindgut, not otherwise specified
C2349358|T191|AB|209.69|ICD9CM|Bengn carcinoid oth site|Bengn carcinoid oth site
C2349358|T191|PT|209.69|ICD9CM|Benign carcinoid tumor of other sites|Benign carcinoid tumor of other sites
C2712917|T191|HT|209.7|ICD9CM|Secondary neuroendocrine tumors|Secondary neuroendocrine tumors
C2712749|T191|AB|209.70|ICD9CM|Sec neuroendo tumor NOS|Sec neuroendo tumor NOS
C2712749|T191|PT|209.70|ICD9CM|Secondary neuroendocrine tumor, unspecified site|Secondary neuroendocrine tumor, unspecified site
C2712873|T191|AB|209.71|ICD9CM|Sec neuroend tu dist lym|Sec neuroend tu dist lym
C2712873|T191|PT|209.71|ICD9CM|Secondary neuroendocrine tumor of distant lymph nodes|Secondary neuroendocrine tumor of distant lymph nodes
C2712885|T191|AB|209.72|ICD9CM|Sec neuroend tumor-liver|Sec neuroend tumor-liver
C2712885|T191|PT|209.72|ICD9CM|Secondary neuroendocrine tumor of liver|Secondary neuroendocrine tumor of liver
C2712897|T191|AB|209.73|ICD9CM|Sec neuroendo tumor-bone|Sec neuroendo tumor-bone
C2712897|T191|PT|209.73|ICD9CM|Secondary neuroendocrine tumor of bone|Secondary neuroendocrine tumor of bone
C2712904|T191|AB|209.74|ICD9CM|Sec neuroendo tu-periton|Sec neuroendo tu-periton
C2712904|T191|PT|209.74|ICD9CM|Secondary neuroendocrine tumor of peritoneum|Secondary neuroendocrine tumor of peritoneum
C2712933|T191|AB|209.75|ICD9CM|Secondary Merkel cell ca|Secondary Merkel cell ca
C2712933|T191|PT|209.75|ICD9CM|Secondary Merkel cell carcinoma|Secondary Merkel cell carcinoma
C2712796|T191|AB|209.79|ICD9CM|Sec neuroend tu oth site|Sec neuroend tu oth site
C2712796|T191|PT|209.79|ICD9CM|Secondary neuroendocrine tumor of other sites|Secondary neuroendocrine tumor of other sites
C0153931|T191|HT|210|ICD9CM|Benign neoplasm of lip, oral cavity, and pharynx|Benign neoplasm of lip, oral cavity, and pharynx
C0086692|T191|HT|210-229.99|ICD9CM|BENIGN NEOPLASMS|BENIGN NEOPLASMS
C0153932|T191|AB|210.0|ICD9CM|Benign neoplasm lip|Benign neoplasm lip
C0153932|T191|PT|210.0|ICD9CM|Benign neoplasm of lip|Benign neoplasm of lip
C0153933|T191|PT|210.1|ICD9CM|Benign neoplasm of tongue|Benign neoplasm of tongue
C0153933|T191|AB|210.1|ICD9CM|Benign neoplasm tongue|Benign neoplasm tongue
C0496858|T191|AB|210.2|ICD9CM|Ben neo major salivary|Ben neo major salivary
C0496858|T191|PT|210.2|ICD9CM|Benign neoplasm of major salivary glands|Benign neoplasm of major salivary glands
C0153934|T191|AB|210.3|ICD9CM|Benign neo mouth floor|Benign neo mouth floor
C0153934|T191|PT|210.3|ICD9CM|Benign neoplasm of floor of mouth|Benign neoplasm of floor of mouth
C0153935|T191|AB|210.4|ICD9CM|Benign neo mouth NEC/NOS|Benign neo mouth NEC/NOS
C0153935|T191|PT|210.4|ICD9CM|Benign neoplasm of other and unspecified parts of mouth|Benign neoplasm of other and unspecified parts of mouth
C0153936|T191|PT|210.5|ICD9CM|Benign neoplasm of tonsil|Benign neoplasm of tonsil
C0153936|T191|AB|210.5|ICD9CM|Benign neoplasm tonsil|Benign neoplasm tonsil
C0153937|T191|AB|210.6|ICD9CM|Benign neo oropharyn NEC|Benign neo oropharyn NEC
C0153937|T191|PT|210.6|ICD9CM|Benign neoplasm of other parts of oropharynx|Benign neoplasm of other parts of oropharynx
C0153938|T191|AB|210.7|ICD9CM|Benign neo nasopharynx|Benign neo nasopharynx
C0153938|T191|PT|210.7|ICD9CM|Benign neoplasm of nasopharynx|Benign neoplasm of nasopharynx
C0153939|T191|AB|210.8|ICD9CM|Benign neo hypopharynx|Benign neo hypopharynx
C0153939|T191|PT|210.8|ICD9CM|Benign neoplasm of hypopharynx|Benign neoplasm of hypopharynx
C0153940|T191|AB|210.9|ICD9CM|Benign neo pharynx NOS|Benign neo pharynx NOS
C0153940|T191|PT|210.9|ICD9CM|Benign neoplasm of pharynx, unspecified|Benign neoplasm of pharynx, unspecified
C0497538|T191|HT|211|ICD9CM|Benign neoplasm of other parts of digestive system|Benign neoplasm of other parts of digestive system
C0153942|T191|AB|211.0|ICD9CM|Benign neo esophagus|Benign neo esophagus
C0153942|T191|PT|211.0|ICD9CM|Benign neoplasm of esophagus|Benign neoplasm of esophagus
C0153943|T191|PT|211.1|ICD9CM|Benign neoplasm of stomach|Benign neoplasm of stomach
C0153943|T191|AB|211.1|ICD9CM|Benign neoplasm stomach|Benign neoplasm stomach
C0153944|T191|PT|211.2|ICD9CM|Benign neoplasm of duodenum, jejunum, and ileum|Benign neoplasm of duodenum, jejunum, and ileum
C0153944|T191|AB|211.2|ICD9CM|Benign neoplasm sm bowel|Benign neoplasm sm bowel
C0004991|T191|AB|211.3|ICD9CM|Benign neoplasm lg bowel|Benign neoplasm lg bowel
C0004991|T191|PT|211.3|ICD9CM|Benign neoplasm of colon|Benign neoplasm of colon
C0153945|T191|AB|211.4|ICD9CM|Benign neopl rectum/anus|Benign neopl rectum/anus
C0153945|T191|PT|211.4|ICD9CM|Benign neoplasm of rectum and anal canal|Benign neoplasm of rectum and anal canal
C0347277|T191|AB|211.5|ICD9CM|Ben neo liver/bile ducts|Ben neo liver/bile ducts
C0347277|T191|PT|211.5|ICD9CM|Benign neoplasm of liver and biliary passages|Benign neoplasm of liver and biliary passages
C0347924|T191|PT|211.6|ICD9CM|Benign neoplasm of pancreas, except islets of Langerhans|Benign neoplasm of pancreas, except islets of Langerhans
C0347924|T191|AB|211.6|ICD9CM|Benign neoplasm pancreas|Benign neoplasm pancreas
C0496872|T191|AB|211.7|ICD9CM|Ben neo islets langerhan|Ben neo islets langerhan
C0496872|T191|PT|211.7|ICD9CM|Benign neoplasm of islets of Langerhans|Benign neoplasm of islets of Langerhans
C0347406|T191|AB|211.8|ICD9CM|Ben neo peritoneum|Ben neo peritoneum
C0347406|T191|PT|211.8|ICD9CM|Benign neoplasm of retroperitoneum and peritoneum|Benign neoplasm of retroperitoneum and peritoneum
C0497538|T191|AB|211.9|ICD9CM|Ben neo GI tract NEC/NOS|Ben neo GI tract NEC/NOS
C0497538|T191|PT|211.9|ICD9CM|Benign neoplasm of other and unspecified site in the digestive system|Benign neoplasm of other and unspecified site in the digestive system
C0347243|T191|HT|212|ICD9CM|Benign neoplasm of respiratory and intrathoracic organs|Benign neoplasm of respiratory and intrathoracic organs
C0153951|T191|AB|212.0|ICD9CM|Ben neo nasal cav/sinus|Ben neo nasal cav/sinus
C0153951|T191|PT|212.0|ICD9CM|Benign neoplasm of nasal cavities, middle ear, and accessory sinuses|Benign neoplasm of nasal cavities, middle ear, and accessory sinuses
C0153952|T191|AB|212.1|ICD9CM|Benign neo larynx|Benign neo larynx
C0153952|T191|PT|212.1|ICD9CM|Benign neoplasm of larynx|Benign neoplasm of larynx
C0153953|T191|AB|212.2|ICD9CM|Benign neo trachea|Benign neo trachea
C0153953|T191|PT|212.2|ICD9CM|Benign neoplasm of trachea|Benign neoplasm of trachea
C0153954|T191|AB|212.3|ICD9CM|Benign neo bronchus/lung|Benign neo bronchus/lung
C0153954|T191|PT|212.3|ICD9CM|Benign neoplasm of bronchus and lung|Benign neoplasm of bronchus and lung
C0153955|T191|PT|212.4|ICD9CM|Benign neoplasm of pleura|Benign neoplasm of pleura
C0153955|T191|AB|212.4|ICD9CM|Benign neoplasm pleura|Benign neoplasm pleura
C0153956|T191|AB|212.5|ICD9CM|Benign neo mediastinum|Benign neo mediastinum
C0153956|T191|PT|212.5|ICD9CM|Benign neoplasm of mediastinum|Benign neoplasm of mediastinum
C0345975|T191|PT|212.6|ICD9CM|Benign neoplasm of thymus|Benign neoplasm of thymus
C0345975|T191|AB|212.6|ICD9CM|Benign neoplasm thymus|Benign neoplasm thymus
C0153957|T191|AB|212.7|ICD9CM|Benign neoplasm heart|Benign neoplasm heart
C0153957|T191|PT|212.7|ICD9CM|Benign neoplasm of heart|Benign neoplasm of heart
C0153958|T191|AB|212.8|ICD9CM|Benign neo resp sys NEC|Benign neo resp sys NEC
C0153958|T191|PT|212.8|ICD9CM|Benign neoplasm of other specified sites of respiratory and intrathoracic organs|Benign neoplasm of other specified sites of respiratory and intrathoracic organs
C0347243|T191|AB|212.9|ICD9CM|Benign neo resp sys NOS|Benign neo resp sys NOS
C0347243|T191|PT|212.9|ICD9CM|Benign neoplasm of respiratory and intrathoracic organs, site unspecified|Benign neoplasm of respiratory and intrathoracic organs, site unspecified
C0153959|T191|HT|213|ICD9CM|Benign neoplasm of bone and articular cartilage|Benign neoplasm of bone and articular cartilage
C0153960|T191|AB|213.0|ICD9CM|Ben neo skull/face bone|Ben neo skull/face bone
C0153960|T191|PT|213.0|ICD9CM|Benign neoplasm of bones of skull and face|Benign neoplasm of bones of skull and face
C0004994|T191|AB|213.1|ICD9CM|Ben neo lower jaw bone|Ben neo lower jaw bone
C0004994|T191|PT|213.1|ICD9CM|Benign neoplasm of lower jaw bone|Benign neoplasm of lower jaw bone
C0702197|T191|AB|213.2|ICD9CM|Benign neo vertebrae|Benign neo vertebrae
C0702197|T191|PT|213.2|ICD9CM|Benign neoplasm of vertebral column, excluding sacrum and coccyx|Benign neoplasm of vertebral column, excluding sacrum and coccyx
C0153962|T191|AB|213.3|ICD9CM|Ben neo ribs/stern/clav|Ben neo ribs/stern/clav
C0153962|T191|PT|213.3|ICD9CM|Benign neoplasm of ribs, sternum, and clavicle|Benign neoplasm of ribs, sternum, and clavicle
C0153963|T191|AB|213.4|ICD9CM|Ben neo long bones arm|Ben neo long bones arm
C0153963|T191|PT|213.4|ICD9CM|Benign neoplasm of scapula and long bones of upper limb|Benign neoplasm of scapula and long bones of upper limb
C0153964|T191|AB|213.5|ICD9CM|Ben neo bones wrist/hand|Ben neo bones wrist/hand
C0153964|T191|PT|213.5|ICD9CM|Benign neoplasm of short bones of upper limb|Benign neoplasm of short bones of upper limb
C0153965|T191|AB|213.6|ICD9CM|Benign neo pelvic girdle|Benign neo pelvic girdle
C0153965|T191|PT|213.6|ICD9CM|Benign neoplasm of pelvic bones, sacrum, and coccyx|Benign neoplasm of pelvic bones, sacrum, and coccyx
C0153966|T191|AB|213.7|ICD9CM|Ben neo long bones leg|Ben neo long bones leg
C0153966|T191|PT|213.7|ICD9CM|Benign neoplasm of long bones of lower limb|Benign neoplasm of long bones of lower limb
C0153967|T191|AB|213.8|ICD9CM|Ben neo bones ankle/foot|Ben neo bones ankle/foot
C0153967|T191|PT|213.8|ICD9CM|Benign neoplasm of short bones of lower limb|Benign neoplasm of short bones of lower limb
C0153959|T191|AB|213.9|ICD9CM|Benign neo bone NOS|Benign neo bone NOS
C0153959|T191|PT|213.9|ICD9CM|Benign neoplasm of bone and articular cartilage, site unspecified|Benign neoplasm of bone and articular cartilage, site unspecified
C0023798|T191|HT|214|ICD9CM|Lipoma|Lipoma
C0153968|T191|PT|214.0|ICD9CM|Lipoma of skin and subcutaneous tissue of face|Lipoma of skin and subcutaneous tissue of face
C0153968|T191|AB|214.0|ICD9CM|Lipoma skin face|Lipoma skin face
C0153969|T191|PT|214.1|ICD9CM|Lipoma of other skin and subcutaneous tissue|Lipoma of other skin and subcutaneous tissue
C0153969|T191|AB|214.1|ICD9CM|Lipoma skin NEC|Lipoma skin NEC
C0153970|T191|AB|214.2|ICD9CM|Lipoma intrathoracic|Lipoma intrathoracic
C0153970|T191|PT|214.2|ICD9CM|Lipoma of intrathoracic organs|Lipoma of intrathoracic organs
C0153971|T191|AB|214.3|ICD9CM|Lipoma intra-abdominal|Lipoma intra-abdominal
C0153971|T191|PT|214.3|ICD9CM|Lipoma of intra-abdominal organs|Lipoma of intra-abdominal organs
C0153972|T191|PT|214.4|ICD9CM|Lipoma of spermatic cord|Lipoma of spermatic cord
C0153972|T191|AB|214.4|ICD9CM|Lipoma spermatic cord|Lipoma spermatic cord
C0023800|T191|AB|214.8|ICD9CM|Lipoma NEC|Lipoma NEC
C0023800|T191|PT|214.8|ICD9CM|Lipoma of other specified sites|Lipoma of other specified sites
C0023798|T191|AB|214.9|ICD9CM|Lipoma NOS|Lipoma NOS
C0023798|T191|PT|214.9|ICD9CM|Lipoma, unspecified site|Lipoma, unspecified site
C0496876|T191|HT|215|ICD9CM|Other benign neoplasm of connective and other soft tissue|Other benign neoplasm of connective and other soft tissue
C0153974|T191|AB|215.0|ICD9CM|Ben neo soft tissue head|Ben neo soft tissue head
C0153974|T191|PT|215.0|ICD9CM|Other benign neoplasm of connective and other soft tissue of head, face, and neck|Other benign neoplasm of connective and other soft tissue of head, face, and neck
C0153975|T191|AB|215.2|ICD9CM|Ben neo soft tissue arm|Ben neo soft tissue arm
C0153975|T191|PT|215.2|ICD9CM|Other benign neoplasm of connective and other soft tissue of upper limb, including shoulder|Other benign neoplasm of connective and other soft tissue of upper limb, including shoulder
C0153976|T191|AB|215.3|ICD9CM|Ben neo soft tissue leg|Ben neo soft tissue leg
C0153976|T191|PT|215.3|ICD9CM|Other benign neoplasm of connective and other soft tissue of lower limb, including hip|Other benign neoplasm of connective and other soft tissue of lower limb, including hip
C0153977|T191|AB|215.4|ICD9CM|Ben neo soft tis thorax|Ben neo soft tis thorax
C0153977|T191|PT|215.4|ICD9CM|Other benign neoplasm of connective and other soft tissue of thorax|Other benign neoplasm of connective and other soft tissue of thorax
C0153978|T191|AB|215.5|ICD9CM|Ben neo soft tis abdomen|Ben neo soft tis abdomen
C0153978|T191|PT|215.5|ICD9CM|Other benign neoplasm of connective and other soft tissue of abdomen|Other benign neoplasm of connective and other soft tissue of abdomen
C0153979|T191|AB|215.6|ICD9CM|Ben neo soft tis pelvis|Ben neo soft tis pelvis
C0153979|T191|PT|215.6|ICD9CM|Other benign neoplasm of connective and other soft tissue of pelvis|Other benign neoplasm of connective and other soft tissue of pelvis
C0375098|T191|AB|215.7|ICD9CM|Benign neo trunk NOS|Benign neo trunk NOS
C0375098|T191|PT|215.7|ICD9CM|Other benign neoplasm of connective and other soft tissue of trunk, unspecified|Other benign neoplasm of connective and other soft tissue of trunk, unspecified
C0153981|T191|AB|215.8|ICD9CM|Ben neo soft tissue NEC|Ben neo soft tissue NEC
C0153981|T191|PT|215.8|ICD9CM|Other benign neoplasm of connective and other soft tissue of other specified sites|Other benign neoplasm of connective and other soft tissue of other specified sites
C0496876|T191|AB|215.9|ICD9CM|Ben neo soft tissue NOS|Ben neo soft tissue NOS
C0496876|T191|PT|215.9|ICD9CM|Other benign neoplasm of connective and other soft tissue, site unspecified|Other benign neoplasm of connective and other soft tissue, site unspecified
C0004998|T191|HT|216|ICD9CM|Benign neoplasm of skin|Benign neoplasm of skin
C0153982|T191|AB|216.0|ICD9CM|Benign neo skin lip|Benign neo skin lip
C0153982|T191|PT|216.0|ICD9CM|Benign neoplasm of skin of lip|Benign neoplasm of skin of lip
C0153983|T191|AB|216.1|ICD9CM|Benign neo skin eyelid|Benign neo skin eyelid
C0153983|T191|PT|216.1|ICD9CM|Benign neoplasm of eyelid, including canthus|Benign neoplasm of eyelid, including canthus
C0153984|T191|AB|216.2|ICD9CM|Benign neo skin ear|Benign neo skin ear
C0153984|T191|PT|216.2|ICD9CM|Benign neoplasm of ear and external auditory canal|Benign neoplasm of ear and external auditory canal
C0153985|T191|AB|216.3|ICD9CM|Benign neo skin face NEC|Benign neo skin face NEC
C0153985|T191|PT|216.3|ICD9CM|Benign neoplasm of skin of other and unspecified parts of face|Benign neoplasm of skin of other and unspecified parts of face
C0153986|T191|AB|216.4|ICD9CM|Ben neo scalp/skin neck|Ben neo scalp/skin neck
C0153986|T191|PT|216.4|ICD9CM|Benign neoplasm of scalp and skin of neck|Benign neoplasm of scalp and skin of neck
C0153987|T191|AB|216.5|ICD9CM|Benign neo skin trunk|Benign neo skin trunk
C0153987|T191|PT|216.5|ICD9CM|Benign neoplasm of skin of trunk, except scrotum|Benign neoplasm of skin of trunk, except scrotum
C0153988|T191|AB|216.6|ICD9CM|Benign neo skin arm|Benign neo skin arm
C0153988|T191|PT|216.6|ICD9CM|Benign neoplasm of skin of upper limb, including shoulder|Benign neoplasm of skin of upper limb, including shoulder
C0153989|T191|AB|216.7|ICD9CM|Benign neo skin leg|Benign neo skin leg
C0153989|T191|PT|216.7|ICD9CM|Benign neoplasm of skin of lower limb, including hip|Benign neoplasm of skin of lower limb, including hip
C0153990|T191|PT|216.8|ICD9CM|Benign neoplasm of other specified sites of skin|Benign neoplasm of other specified sites of skin
C0153990|T191|AB|216.8|ICD9CM|Benign neoplasm skin NEC|Benign neoplasm skin NEC
C0004998|T191|PT|216.9|ICD9CM|Benign neoplasm of skin, site unspecified|Benign neoplasm of skin, site unspecified
C0004998|T191|AB|216.9|ICD9CM|Benign neoplasm skin NOS|Benign neoplasm skin NOS
C0346156|T191|AB|217|ICD9CM|Benign neoplasm breast|Benign neoplasm breast
C0346156|T191|PT|217|ICD9CM|Benign neoplasm of breast|Benign neoplasm of breast
C0042133|T191|HT|218|ICD9CM|Uterine leiomyoma|Uterine leiomyoma
C0153993|T191|AB|218.0|ICD9CM|Submucous leiomyoma|Submucous leiomyoma
C0153993|T191|PT|218.0|ICD9CM|Submucous leiomyoma of uterus|Submucous leiomyoma of uterus
C0153994|T191|AB|218.1|ICD9CM|Intramural leiomyoma|Intramural leiomyoma
C0153994|T191|PT|218.1|ICD9CM|Intramural leiomyoma of uterus|Intramural leiomyoma of uterus
C0153995|T191|AB|218.2|ICD9CM|Subserous leiomyoma|Subserous leiomyoma
C0153995|T191|PT|218.2|ICD9CM|Subserous leiomyoma of uterus|Subserous leiomyoma of uterus
C0042133|T191|PT|218.9|ICD9CM|Leiomyoma of uterus, unspecified|Leiomyoma of uterus, unspecified
C0042133|T191|AB|218.9|ICD9CM|Uterine leiomyoma NOS|Uterine leiomyoma NOS
C0153996|T191|HT|219|ICD9CM|Other benign neoplasm of uterus|Other benign neoplasm of uterus
C0153997|T191|AB|219.0|ICD9CM|Benign neo cervix uteri|Benign neo cervix uteri
C0153997|T191|PT|219.0|ICD9CM|Benign neoplasm of cervix uteri|Benign neoplasm of cervix uteri
C0153998|T191|AB|219.1|ICD9CM|Benign neo corpus uteri|Benign neo corpus uteri
C0153998|T191|PT|219.1|ICD9CM|Benign neoplasm of corpus uteri|Benign neoplasm of corpus uteri
C0347491|T191|AB|219.8|ICD9CM|Benign neo uterus NEC|Benign neo uterus NEC
C0347491|T191|PT|219.8|ICD9CM|Benign neoplasm of other specified parts of uterus|Benign neoplasm of other specified parts of uterus
C0153999|T191|AB|219.9|ICD9CM|Benign neo uterus NOS|Benign neo uterus NOS
C0153999|T191|PT|219.9|ICD9CM|Benign neoplasm of uterus, part unspecified|Benign neoplasm of uterus, part unspecified
C0004997|T191|PT|220|ICD9CM|Benign neoplasm of ovary|Benign neoplasm of ovary
C0004997|T191|AB|220|ICD9CM|Benign neoplasm ovary|Benign neoplasm ovary
C0154000|T191|HT|221|ICD9CM|Benign neoplasm of other female genital organs|Benign neoplasm of other female genital organs
C0496889|T191|AB|221.0|ICD9CM|Ben neo fallopian tube|Ben neo fallopian tube
C0496889|T191|PT|221.0|ICD9CM|Benign neoplasm of fallopian tube and uterine ligaments|Benign neoplasm of fallopian tube and uterine ligaments
C0154002|T191|PT|221.1|ICD9CM|Benign neoplasm of vagina|Benign neoplasm of vagina
C0154002|T191|AB|221.1|ICD9CM|Benign neoplasm vagina|Benign neoplasm vagina
C0154003|T191|PT|221.2|ICD9CM|Benign neoplasm of vulva|Benign neoplasm of vulva
C0154003|T191|AB|221.2|ICD9CM|Benign neoplasm vulva|Benign neoplasm vulva
C0154004|T191|AB|221.8|ICD9CM|Ben neo fem genital NEC|Ben neo fem genital NEC
C0154004|T191|PT|221.8|ICD9CM|Benign neoplasm of other specified sites of female genital organs|Benign neoplasm of other specified sites of female genital organs
C0154005|T191|AB|221.9|ICD9CM|Ben neo fem genital NOS|Ben neo fem genital NOS
C0154005|T191|PT|221.9|ICD9CM|Benign neoplasm of female genital organ, site unspecified|Benign neoplasm of female genital organ, site unspecified
C0496891|T191|HT|222|ICD9CM|Benign neoplasm of male genital organs|Benign neoplasm of male genital organs
C0154007|T191|PT|222.0|ICD9CM|Benign neoplasm of testis|Benign neoplasm of testis
C0154007|T191|AB|222.0|ICD9CM|Benign neoplasm testis|Benign neoplasm testis
C0149627|T191|PT|222.1|ICD9CM|Benign neoplasm of penis|Benign neoplasm of penis
C0149627|T191|AB|222.1|ICD9CM|Benign neoplasm penis|Benign neoplasm penis
C0154009|T191|PT|222.2|ICD9CM|Benign neoplasm of prostate|Benign neoplasm of prostate
C0154009|T191|AB|222.2|ICD9CM|Benign neoplasm prostate|Benign neoplasm prostate
C0154010|T191|AB|222.3|ICD9CM|Benign neo epididymis|Benign neo epididymis
C0154010|T191|PT|222.3|ICD9CM|Benign neoplasm of epididymis|Benign neoplasm of epididymis
C0154011|T191|PT|222.4|ICD9CM|Benign neoplasm of scrotum|Benign neoplasm of scrotum
C0154011|T191|AB|222.4|ICD9CM|Benign neoplasm scrotum|Benign neoplasm scrotum
C0154012|T191|AB|222.8|ICD9CM|Ben neo male genital NEC|Ben neo male genital NEC
C0154012|T191|PT|222.8|ICD9CM|Benign neoplasm of other specified sites of male genital organs|Benign neoplasm of other specified sites of male genital organs
C0496891|T191|AB|222.9|ICD9CM|Ben neo male genital NOS|Ben neo male genital NOS
C0496891|T191|PT|222.9|ICD9CM|Benign neoplasm of male genital organ, site unspecified|Benign neoplasm of male genital organ, site unspecified
C0154013|T191|HT|223|ICD9CM|Benign neoplasm of kidney and other urinary organs|Benign neoplasm of kidney and other urinary organs
C0154014|T191|AB|223.0|ICD9CM|Benign neoplasm kidney|Benign neoplasm kidney
C0154014|T191|PT|223.0|ICD9CM|Benign neoplasm of kidney, except pelvis|Benign neoplasm of kidney, except pelvis
C0154015|T191|AB|223.1|ICD9CM|Benign neo renal pelvis|Benign neo renal pelvis
C0154015|T191|PT|223.1|ICD9CM|Benign neoplasm of renal pelvis|Benign neoplasm of renal pelvis
C0154016|T191|PT|223.2|ICD9CM|Benign neoplasm of ureter|Benign neoplasm of ureter
C0154016|T191|AB|223.2|ICD9CM|Benign neoplasm ureter|Benign neoplasm ureter
C0154017|T191|AB|223.3|ICD9CM|Benign neoplasm bladder|Benign neoplasm bladder
C0154017|T191|PT|223.3|ICD9CM|Benign neoplasm of bladder|Benign neoplasm of bladder
C0154018|T191|HT|223.8|ICD9CM|Benign neoplasm of other specified sites of urinary organs|Benign neoplasm of other specified sites of urinary organs
C0154019|T191|PT|223.81|ICD9CM|Benign neoplasm of urethra|Benign neoplasm of urethra
C0154019|T191|AB|223.81|ICD9CM|Benign neoplasm urethra|Benign neoplasm urethra
C0154018|T191|AB|223.89|ICD9CM|Benign neo urinary NEC|Benign neo urinary NEC
C0154018|T191|PT|223.89|ICD9CM|Benign neoplasm of other specified sites of urinary organs|Benign neoplasm of other specified sites of urinary organs
C0496893|T191|AB|223.9|ICD9CM|Benign neo urinary NOS|Benign neo urinary NOS
C0496893|T191|PT|223.9|ICD9CM|Benign neoplasm of urinary organ, site unspecified|Benign neoplasm of urinary organ, site unspecified
C0496897|T191|HT|224|ICD9CM|Benign neoplasm of eye|Benign neoplasm of eye
C0154022|T191|AB|224.0|ICD9CM|Benign neoplasm eyeball|Benign neoplasm eyeball
C0154022|T191|PT|224.0|ICD9CM|Benign neoplasm of eyeball, except conjunctiva, cornea, retina, and choroid|Benign neoplasm of eyeball, except conjunctiva, cornea, retina, and choroid
C0154023|T191|PT|224.1|ICD9CM|Benign neoplasm of orbit|Benign neoplasm of orbit
C0154023|T191|AB|224.1|ICD9CM|Benign neoplasm orbit|Benign neoplasm orbit
C0154024|T191|AB|224.2|ICD9CM|Ben neo lacrimal gland|Ben neo lacrimal gland
C0154024|T191|PT|224.2|ICD9CM|Benign neoplasm of lacrimal gland|Benign neoplasm of lacrimal gland
C0154025|T191|AB|224.3|ICD9CM|Benign neo conjunctiva|Benign neo conjunctiva
C0154025|T191|PT|224.3|ICD9CM|Benign neoplasm of conjunctiva|Benign neoplasm of conjunctiva
C0154026|T191|AB|224.4|ICD9CM|Benign neoplasm cornea|Benign neoplasm cornea
C0154026|T191|PT|224.4|ICD9CM|Benign neoplasm of cornea|Benign neoplasm of cornea
C0154027|T191|PT|224.5|ICD9CM|Benign neoplasm of retina|Benign neoplasm of retina
C0154027|T191|AB|224.5|ICD9CM|Benign neoplasm retina|Benign neoplasm retina
C0154028|T191|AB|224.6|ICD9CM|Benign neoplasm choroid|Benign neoplasm choroid
C0154028|T191|PT|224.6|ICD9CM|Benign neoplasm of choroid|Benign neoplasm of choroid
C0154029|T191|AB|224.7|ICD9CM|Ben neo lacrimal duct|Ben neo lacrimal duct
C0154029|T191|PT|224.7|ICD9CM|Benign neoplasm of lacrimal duct|Benign neoplasm of lacrimal duct
C0154030|T191|AB|224.8|ICD9CM|Benign neoplasm eye NEC|Benign neoplasm eye NEC
C0154030|T191|PT|224.8|ICD9CM|Benign neoplasm of other specified parts of eye|Benign neoplasm of other specified parts of eye
C0496897|T191|AB|224.9|ICD9CM|Benign neoplasm eye NOS|Benign neoplasm eye NOS
C0496897|T191|PT|224.9|ICD9CM|Benign neoplasm of eye, part unspecified|Benign neoplasm of eye, part unspecified
C0497550|T191|HT|225|ICD9CM|Benign neoplasm of brain and other parts of nervous system|Benign neoplasm of brain and other parts of nervous system
C0496899|T191|AB|225.0|ICD9CM|Benign neoplasm brain|Benign neoplasm brain
C0496899|T191|PT|225.0|ICD9CM|Benign neoplasm of brain|Benign neoplasm of brain
C0004992|T191|AB|225.1|ICD9CM|Benign neo cranial nerve|Benign neo cranial nerve
C0004992|T191|PT|225.1|ICD9CM|Benign neoplasm of cranial nerves|Benign neoplasm of cranial nerves
C0154033|T191|AB|225.2|ICD9CM|Ben neo cerebr meninges|Ben neo cerebr meninges
C0154033|T191|PT|225.2|ICD9CM|Benign neoplasm of cerebral meninges|Benign neoplasm of cerebral meninges
C0154034|T191|AB|225.3|ICD9CM|Benign neo spinal cord|Benign neo spinal cord
C0154034|T191|PT|225.3|ICD9CM|Benign neoplasm of spinal cord|Benign neoplasm of spinal cord
C0154035|T191|AB|225.4|ICD9CM|Ben neo spinal meninges|Ben neo spinal meninges
C0154035|T191|PT|225.4|ICD9CM|Benign neoplasm of spinal meninges|Benign neoplasm of spinal meninges
C0154036|T191|AB|225.8|ICD9CM|Benign neo nerv sys NEC|Benign neo nerv sys NEC
C0154036|T191|PT|225.8|ICD9CM|Benign neoplasm of other specified sites of nervous system|Benign neoplasm of other specified sites of nervous system
C0497550|T191|AB|225.9|ICD9CM|Benign neo nerv sys NOS|Benign neo nerv sys NOS
C0497550|T191|PT|225.9|ICD9CM|Benign neoplasm of nervous system, part unspecified|Benign neoplasm of nervous system, part unspecified
C0154038|T191|PT|226|ICD9CM|Benign neoplasm of thyroid glands|Benign neoplasm of thyroid glands
C0154038|T191|AB|226|ICD9CM|Benign neoplasm thyroid|Benign neoplasm thyroid
C0154039|T191|HT|227|ICD9CM|Benign neoplasm of other endocrine glands and related structures|Benign neoplasm of other endocrine glands and related structures
C0154040|T191|AB|227.0|ICD9CM|Benign neoplasm adrenal|Benign neoplasm adrenal
C0154040|T191|PT|227.0|ICD9CM|Benign neoplasm of adrenal gland|Benign neoplasm of adrenal gland
C0154041|T191|AB|227.1|ICD9CM|Benign neo parathyroid|Benign neo parathyroid
C0154041|T191|PT|227.1|ICD9CM|Benign neoplasm of parathyroid gland|Benign neoplasm of parathyroid gland
C0347525|T191|AB|227.3|ICD9CM|Benign neo pituitary|Benign neo pituitary
C0347525|T191|PT|227.3|ICD9CM|Benign neoplasm of pituitary gland and craniopharyngeal duct|Benign neoplasm of pituitary gland and craniopharyngeal duct
C0154043|T191|AB|227.4|ICD9CM|Ben neopl pineal gland|Ben neopl pineal gland
C0154043|T191|PT|227.4|ICD9CM|Benign neoplasm of pineal gland|Benign neoplasm of pineal gland
C0154044|T191|AB|227.5|ICD9CM|Benign neo carotid body|Benign neo carotid body
C0154044|T191|PT|227.5|ICD9CM|Benign neoplasm of carotid body|Benign neoplasm of carotid body
C0154045|T191|AB|227.6|ICD9CM|Ben neo paraganglia NEC|Ben neo paraganglia NEC
C0154045|T191|PT|227.6|ICD9CM|Benign neoplasm of aortic body and other paraganglia|Benign neoplasm of aortic body and other paraganglia
C0154039|T191|AB|227.8|ICD9CM|Benign neo endocrine NEC|Benign neo endocrine NEC
C0154039|T191|PT|227.8|ICD9CM|Benign neoplasm of other endocrine glands and related structures|Benign neoplasm of other endocrine glands and related structures
C0347524|T191|AB|227.9|ICD9CM|Benign neo endocrine NOS|Benign neo endocrine NOS
C0347524|T191|PT|227.9|ICD9CM|Benign neoplasm of endocrine gland, site unspecified|Benign neoplasm of endocrine gland, site unspecified
C0851225|T191|HT|228|ICD9CM|Hemangioma and lymphangioma, any site|Hemangioma and lymphangioma, any site
C0018916|T191|HT|228.0|ICD9CM|Hemangioma, any site|Hemangioma, any site
C0018916|T191|AB|228.00|ICD9CM|Hemangioma NOS|Hemangioma NOS
C0018916|T191|PT|228.00|ICD9CM|Hemangioma of unspecified site|Hemangioma of unspecified site
C0154049|T191|PT|228.01|ICD9CM|Hemangioma of skin and subcutaneous tissue|Hemangioma of skin and subcutaneous tissue
C0154049|T191|AB|228.01|ICD9CM|Hemangioma skin|Hemangioma skin
C0154050|T191|AB|228.02|ICD9CM|Hemangioma intracranial|Hemangioma intracranial
C0154050|T191|PT|228.02|ICD9CM|Hemangioma of intracranial structures|Hemangioma of intracranial structures
C0154051|T191|PT|228.03|ICD9CM|Hemangioma of retina|Hemangioma of retina
C0154051|T191|AB|228.03|ICD9CM|Hemangioma retina|Hemangioma retina
C0154052|T191|AB|228.04|ICD9CM|Hemangioma intra-abdom|Hemangioma intra-abdom
C0154052|T191|PT|228.04|ICD9CM|Hemangioma of intra-abdominal structures|Hemangioma of intra-abdominal structures
C0018918|T191|AB|228.09|ICD9CM|Hemangioma NEC|Hemangioma NEC
C0018918|T191|PT|228.09|ICD9CM|Hemangioma of other sites|Hemangioma of other sites
C0024221|T191|AB|228.1|ICD9CM|Lymphangioma, any site|Lymphangioma, any site
C0024221|T191|PT|228.1|ICD9CM|Lymphangioma, any site|Lymphangioma, any site
C0154053|T191|HT|229|ICD9CM|Benign neoplasm of other and unspecified sites|Benign neoplasm of other and unspecified sites
C0154054|T191|AB|229.0|ICD9CM|Benign neo lymph nodes|Benign neo lymph nodes
C0154054|T191|PT|229.0|ICD9CM|Benign neoplasm of lymph nodes|Benign neoplasm of lymph nodes
C0154055|T191|AB|229.8|ICD9CM|Benign neoplasm NEC|Benign neoplasm NEC
C0154055|T191|PT|229.8|ICD9CM|Benign neoplasm of other specified sites|Benign neoplasm of other specified sites
C0086692|T191|AB|229.9|ICD9CM|Benign neoplasm NOS|Benign neoplasm NOS
C0086692|T191|PT|229.9|ICD9CM|Benign neoplasm of unspecified site|Benign neoplasm of unspecified site
C0154057|T191|HT|230|ICD9CM|Carcinoma in situ of digestive organs|Carcinoma in situ of digestive organs
C0007099|T191|HT|230-234.99|ICD9CM|CARCINOMA IN SITU|CARCINOMA IN SITU
C0154058|T191|AB|230.0|ICD9CM|Ca in situ oral cav/phar|Ca in situ oral cav/phar
C0154058|T191|PT|230.0|ICD9CM|Carcinoma in situ of lip, oral cavity, and pharynx|Carcinoma in situ of lip, oral cavity, and pharynx
C0154059|T191|AB|230.1|ICD9CM|Ca in situ esophagus|Ca in situ esophagus
C0154059|T191|PT|230.1|ICD9CM|Carcinoma in situ of esophagus|Carcinoma in situ of esophagus
C0154060|T191|AB|230.2|ICD9CM|Ca in situ stomach|Ca in situ stomach
C0154060|T191|PT|230.2|ICD9CM|Carcinoma in situ of stomach|Carcinoma in situ of stomach
C0154061|T191|AB|230.3|ICD9CM|Ca in situ colon|Ca in situ colon
C0154061|T191|PT|230.3|ICD9CM|Carcinoma in situ of colon|Carcinoma in situ of colon
C0154062|T191|AB|230.4|ICD9CM|Ca in situ rectum|Ca in situ rectum
C0154062|T191|PT|230.4|ICD9CM|Carcinoma in situ of rectum|Carcinoma in situ of rectum
C2242854|T191|AB|230.5|ICD9CM|Ca in situ anal canal|Ca in situ anal canal
C2242854|T191|PT|230.5|ICD9CM|Carcinoma in situ of anal canal|Carcinoma in situ of anal canal
C0154064|T191|AB|230.6|ICD9CM|Ca in situ anus NOS|Ca in situ anus NOS
C0154064|T191|PT|230.6|ICD9CM|Carcinoma in situ of anus, unspecified|Carcinoma in situ of anus, unspecified
C0154065|T191|AB|230.7|ICD9CM|Ca in situ bowel NEC/NOS|Ca in situ bowel NEC/NOS
C0154065|T191|PT|230.7|ICD9CM|Carcinoma in situ of other and unspecified parts of intestine|Carcinoma in situ of other and unspecified parts of intestine
C0496854|T191|AB|230.8|ICD9CM|Ca in situ liver/biliary|Ca in situ liver/biliary
C0496854|T191|PT|230.8|ICD9CM|Carcinoma in situ of liver and biliary system|Carcinoma in situ of liver and biliary system
C0154067|T191|AB|230.9|ICD9CM|Ca in situ GI NEC/NOS|Ca in situ GI NEC/NOS
C0154067|T191|PT|230.9|ICD9CM|Carcinoma in situ of other and unspecified digestive organs|Carcinoma in situ of other and unspecified digestive organs
C0348402|T191|HT|231|ICD9CM|Carcinoma in situ of respiratory system|Carcinoma in situ of respiratory system
C0154069|T191|AB|231.0|ICD9CM|Ca in situ larynx|Ca in situ larynx
C0154069|T191|PT|231.0|ICD9CM|Carcinoma in situ of larynx|Carcinoma in situ of larynx
C0154070|T191|AB|231.1|ICD9CM|Ca in situ trachea|Ca in situ trachea
C0154070|T191|PT|231.1|ICD9CM|Carcinoma in situ of trachea|Carcinoma in situ of trachea
C0154071|T191|AB|231.2|ICD9CM|Ca in situ bronchus/lung|Ca in situ bronchus/lung
C0154071|T191|PT|231.2|ICD9CM|Carcinoma in situ of bronchus and lung|Carcinoma in situ of bronchus and lung
C0154072|T191|AB|231.8|ICD9CM|Ca in situ resp sys NEC|Ca in situ resp sys NEC
C0154072|T191|PT|231.8|ICD9CM|Carcinoma in situ of other specified parts of respiratory system|Carcinoma in situ of other specified parts of respiratory system
C0348402|T191|AB|231.9|ICD9CM|Ca in situ resp sys NOS|Ca in situ resp sys NOS
C0348402|T191|PT|231.9|ICD9CM|Carcinoma in situ of respiratory system, part unspecified|Carcinoma in situ of respiratory system, part unspecified
C0154073|T191|HT|232|ICD9CM|Carcinoma in situ of skin|Carcinoma in situ of skin
C0154074|T191|AB|232.0|ICD9CM|Ca in situ skin lip|Ca in situ skin lip
C0154074|T191|PT|232.0|ICD9CM|Carcinoma in situ of skin of lip|Carcinoma in situ of skin of lip
C0347138|T191|AB|232.1|ICD9CM|Ca in situ eyelid|Ca in situ eyelid
C0347138|T191|PT|232.1|ICD9CM|Carcinoma in situ of eyelid, including canthus|Carcinoma in situ of eyelid, including canthus
C0347139|T191|AB|232.2|ICD9CM|Ca in situ skin ear|Ca in situ skin ear
C0347139|T191|PT|232.2|ICD9CM|Carcinoma in situ of skin of ear and external auditory canal|Carcinoma in situ of skin of ear and external auditory canal
C0154077|T191|AB|232.3|ICD9CM|Ca in situ skin face NEC|Ca in situ skin face NEC
C0154077|T191|PT|232.3|ICD9CM|Carcinoma in situ of skin of other and unspecified parts of face|Carcinoma in situ of skin of other and unspecified parts of face
C0154078|T191|AB|232.4|ICD9CM|Ca in situ scalp|Ca in situ scalp
C0154078|T191|PT|232.4|ICD9CM|Carcinoma in situ of scalp and skin of neck|Carcinoma in situ of scalp and skin of neck
C0154079|T191|AB|232.5|ICD9CM|Ca in situ skin trunk|Ca in situ skin trunk
C0154079|T191|PT|232.5|ICD9CM|Carcinoma in situ of skin of trunk, except scrotum|Carcinoma in situ of skin of trunk, except scrotum
C0154080|T191|AB|232.6|ICD9CM|Ca in situ skin arm|Ca in situ skin arm
C0154080|T191|PT|232.6|ICD9CM|Carcinoma in situ of skin of upper limb, including shoulder|Carcinoma in situ of skin of upper limb, including shoulder
C0154081|T191|AB|232.7|ICD9CM|Ca in situ skin leg|Ca in situ skin leg
C0154081|T191|PT|232.7|ICD9CM|Carcinoma in situ of skin of lower limb, including hip|Carcinoma in situ of skin of lower limb, including hip
C0154082|T191|AB|232.8|ICD9CM|Ca in situ skin NEC|Ca in situ skin NEC
C0154082|T191|PT|232.8|ICD9CM|Carcinoma in situ of other specified sites of skin|Carcinoma in situ of other specified sites of skin
C0154073|T191|AB|232.9|ICD9CM|Ca in situ skin NOS|Ca in situ skin NOS
C0154073|T191|PT|232.9|ICD9CM|Carcinoma in situ of skin, site unspecified|Carcinoma in situ of skin, site unspecified
C0154083|T191|HT|233|ICD9CM|Carcinoma in situ of breast and genitourinary system|Carcinoma in situ of breast and genitourinary system
C0154084|T191|AB|233.0|ICD9CM|Ca in situ breast|Ca in situ breast
C0154084|T191|PT|233.0|ICD9CM|Carcinoma in situ of breast|Carcinoma in situ of breast
C0851140|T191|AB|233.1|ICD9CM|Ca in situ cervix uteri|Ca in situ cervix uteri
C0851140|T191|PT|233.1|ICD9CM|Carcinoma in situ of cervix uteri|Carcinoma in situ of cervix uteri
C0154086|T191|AB|233.2|ICD9CM|Ca in situ uterus NEC|Ca in situ uterus NEC
C0154086|T191|PT|233.2|ICD9CM|Carcinoma in situ of other and unspecified parts of uterus|Carcinoma in situ of other and unspecified parts of uterus
C0154087|T191|HT|233.3|ICD9CM|Carcinoma in situ of other and unspecified female genital organs|Carcinoma in situ of other and unspecified female genital organs
C1955737|T191|AB|233.30|ICD9CM|Ca in situ fem gen NOS|Ca in situ fem gen NOS
C1955737|T191|PT|233.30|ICD9CM|Carcinoma in situ, unspecified female genital organ|Carcinoma in situ, unspecified female genital organ
C0686277|T191|AB|233.31|ICD9CM|Carcinoma in situ vagina|Carcinoma in situ vagina
C0686277|T191|PT|233.31|ICD9CM|Carcinoma in situ, vagina|Carcinoma in situ, vagina
C0278729|T191|AB|233.32|ICD9CM|Carcinoma in situ vulva|Carcinoma in situ vulva
C0278729|T191|PT|233.32|ICD9CM|Carcinoma in situ, vulva|Carcinoma in situ, vulva
C1955739|T191|AB|233.39|ICD9CM|Ca in situ fem gen NEC|Ca in situ fem gen NEC
C1955739|T191|PT|233.39|ICD9CM|Carcinoma in situ, other female genital organ|Carcinoma in situ, other female genital organ
C0154088|T191|AB|233.4|ICD9CM|Ca in situ prostate|Ca in situ prostate
C0154088|T191|PT|233.4|ICD9CM|Carcinoma in situ of prostate|Carcinoma in situ of prostate
C0154089|T191|AB|233.5|ICD9CM|Ca in situ penis|Ca in situ penis
C0154089|T191|PT|233.5|ICD9CM|Carcinoma in situ of penis|Carcinoma in situ of penis
C0154090|T191|AB|233.6|ICD9CM|Ca in situ male gen NEC|Ca in situ male gen NEC
C0154090|T191|PT|233.6|ICD9CM|Carcinoma in situ of other and unspecified male genital organs|Carcinoma in situ of other and unspecified male genital organs
C0154091|T191|AB|233.7|ICD9CM|Ca in situ bladder|Ca in situ bladder
C0154091|T191|PT|233.7|ICD9CM|Carcinoma in situ of bladder|Carcinoma in situ of bladder
C0154092|T191|AB|233.9|ICD9CM|Ca in situ urinary NEC|Ca in situ urinary NEC
C0154092|T191|PT|233.9|ICD9CM|Carcinoma in situ of other and unspecified urinary organs|Carcinoma in situ of other and unspecified urinary organs
C0154093|T191|HT|234|ICD9CM|Carcinoma in situ of other and unspecified sites|Carcinoma in situ of other and unspecified sites
C0154094|T191|AB|234.0|ICD9CM|Ca in situ eye|Ca in situ eye
C0154094|T191|PT|234.0|ICD9CM|Carcinoma in situ of eye|Carcinoma in situ of eye
C0007100|T191|AB|234.8|ICD9CM|Ca in situ NEC|Ca in situ NEC
C0007100|T191|PT|234.8|ICD9CM|Carcinoma in situ of other specified sites|Carcinoma in situ of other specified sites
C0007099|T191|AB|234.9|ICD9CM|Ca in situ NOS|Ca in situ NOS
C0007099|T191|PT|234.9|ICD9CM|Carcinoma in situ, site unspecified|Carcinoma in situ, site unspecified
C0154095|T191|HT|235|ICD9CM|Neoplasm of uncertain behavior of digestive and respiratory systems|Neoplasm of uncertain behavior of digestive and respiratory systems
C0154129|T191|HT|235-238.99|ICD9CM|NEOPLASMS OF UNCERTAIN BEHAVIOR|NEOPLASMS OF UNCERTAIN BEHAVIOR
C0154096|T191|PT|235.0|ICD9CM|Neoplasm of uncertain behavior of major salivary glands|Neoplasm of uncertain behavior of major salivary glands
C0154096|T191|AB|235.0|ICD9CM|Unc behav neo salivary|Unc behav neo salivary
C0154097|T191|PT|235.1|ICD9CM|Neoplasm of uncertain behavior of lip, oral cavity, and pharynx|Neoplasm of uncertain behavior of lip, oral cavity, and pharynx
C0154097|T191|AB|235.1|ICD9CM|Unc behav neo oral/phar|Unc behav neo oral/phar
C0154098|T191|PT|235.2|ICD9CM|Neoplasm of uncertain behavior of stomach, intestines, and rectum|Neoplasm of uncertain behavior of stomach, intestines, and rectum
C0154098|T191|AB|235.2|ICD9CM|Unc behav neo intestine|Unc behav neo intestine
C0496909|T191|PT|235.3|ICD9CM|Neoplasm of uncertain behavior of liver and biliary passages|Neoplasm of uncertain behavior of liver and biliary passages
C0496909|T191|AB|235.3|ICD9CM|Unc behav neo liver|Unc behav neo liver
C0154100|T191|PT|235.4|ICD9CM|Neoplasm of uncertain behavior of retroperitoneum and peritoneum|Neoplasm of uncertain behavior of retroperitoneum and peritoneum
C0154100|T191|AB|235.4|ICD9CM|Unc behav neo peritoneum|Unc behav neo peritoneum
C0154101|T191|PT|235.5|ICD9CM|Neoplasm of uncertain behavior of other and unspecified digestive organs|Neoplasm of uncertain behavior of other and unspecified digestive organs
C0154101|T191|AB|235.5|ICD9CM|Unc behav neo GI NEC|Unc behav neo GI NEC
C0496912|T191|PT|235.6|ICD9CM|Neoplasm of uncertain behavior of larynx|Neoplasm of uncertain behavior of larynx
C0496912|T191|AB|235.6|ICD9CM|Unc behav neo larynx|Unc behav neo larynx
C0154103|T191|PT|235.7|ICD9CM|Neoplasm of uncertain behavior of trachea, bronchus, and lung|Neoplasm of uncertain behavior of trachea, bronchus, and lung
C0154103|T191|AB|235.7|ICD9CM|Unc behav neo lung|Unc behav neo lung
C0154104|T191|PT|235.8|ICD9CM|Neoplasm of uncertain behavior of pleura, thymus, and mediastinum|Neoplasm of uncertain behavior of pleura, thymus, and mediastinum
C0154104|T191|AB|235.8|ICD9CM|Unc behav neo pleura|Unc behav neo pleura
C0154105|T191|PT|235.9|ICD9CM|Neoplasm of uncertain behavior of other and unspecified respiratory organs|Neoplasm of uncertain behavior of other and unspecified respiratory organs
C0154105|T191|AB|235.9|ICD9CM|Unc behav neo resp NEC|Unc behav neo resp NEC
C0154106|T191|HT|236|ICD9CM|Neoplasm of uncertain behavior of genitourinary organs|Neoplasm of uncertain behavior of genitourinary organs
C0496919|T191|PT|236.0|ICD9CM|Neoplasm of uncertain behavior of uterus|Neoplasm of uncertain behavior of uterus
C0496919|T191|AB|236.0|ICD9CM|Uncert behav neo uterus|Uncert behav neo uterus
C0496921|T191|PT|236.1|ICD9CM|Neoplasm of uncertain behavior of placenta|Neoplasm of uncertain behavior of placenta
C0496921|T191|AB|236.1|ICD9CM|Unc behav neo placenta|Unc behav neo placenta
C0496920|T191|PT|236.2|ICD9CM|Neoplasm of uncertain behavior of ovary|Neoplasm of uncertain behavior of ovary
C0496920|T191|AB|236.2|ICD9CM|Unc behav neo ovary|Unc behav neo ovary
C2869595|T191|PT|236.3|ICD9CM|Neoplasm of uncertain behavior of other and unspecified female genital organs|Neoplasm of uncertain behavior of other and unspecified female genital organs
C2869595|T191|AB|236.3|ICD9CM|Unc behav neo female NEC|Unc behav neo female NEC
C0496924|T191|PT|236.4|ICD9CM|Neoplasm of uncertain behavior of testis|Neoplasm of uncertain behavior of testis
C0496924|T191|AB|236.4|ICD9CM|Unc behav neo testis|Unc behav neo testis
C0496923|T191|PT|236.5|ICD9CM|Neoplasm of uncertain behavior of prostate|Neoplasm of uncertain behavior of prostate
C0496923|T191|AB|236.5|ICD9CM|Unc behav neo prostate|Unc behav neo prostate
C2869603|T191|PT|236.6|ICD9CM|Neoplasm of uncertain behavior of other and unspecified male genital organs|Neoplasm of uncertain behavior of other and unspecified male genital organs
C2869603|T191|AB|236.6|ICD9CM|Unc behav neo male NEC|Unc behav neo male NEC
C0496930|T191|PT|236.7|ICD9CM|Neoplasm of uncertain behavior of bladder|Neoplasm of uncertain behavior of bladder
C0496930|T191|AB|236.7|ICD9CM|Unc behav neo bladder|Unc behav neo bladder
C0154113|T191|HT|236.9|ICD9CM|Neoplasm of uncertain behavior of other and unspecified urinary organs|Neoplasm of uncertain behavior of other and unspecified urinary organs
C0496932|T191|PT|236.90|ICD9CM|Neoplasm of uncertain behavior of urinary organ, unspecified|Neoplasm of uncertain behavior of urinary organ, unspecified
C0496932|T191|AB|236.90|ICD9CM|Unc behav neo urinar NOS|Unc behav neo urinar NOS
C0154115|T191|PT|236.91|ICD9CM|Neoplasm of uncertain behavior of kidney and ureter|Neoplasm of uncertain behavior of kidney and ureter
C0154115|T191|AB|236.91|ICD9CM|Unc behav neo kidney|Unc behav neo kidney
C2873698|T191|PT|236.99|ICD9CM|Neoplasm of uncertain behavior of other and unspecified urinary organs|Neoplasm of uncertain behavior of other and unspecified urinary organs
C2873698|T191|AB|236.99|ICD9CM|Unc behav neo urinar NEC|Unc behav neo urinar NEC
C0154116|T191|HT|237|ICD9CM|Neoplasm of uncertain behavior of endocrine glands and nervous system|Neoplasm of uncertain behavior of endocrine glands and nervous system
C0027636|T191|PT|237.0|ICD9CM|Neoplasm of uncertain behavior of pituitary gland and craniopharyngeal duct|Neoplasm of uncertain behavior of pituitary gland and craniopharyngeal duct
C0027636|T191|AB|237.0|ICD9CM|Unc behav neo pituitary|Unc behav neo pituitary
C0496946|T191|PT|237.1|ICD9CM|Neoplasm of uncertain behavior of pineal gland|Neoplasm of uncertain behavior of pineal gland
C0496946|T191|AB|237.1|ICD9CM|Unc behav neo pineal|Unc behav neo pineal
C0154117|T191|PT|237.2|ICD9CM|Neoplasm of uncertain behavior of adrenal gland|Neoplasm of uncertain behavior of adrenal gland
C0154117|T191|AB|237.2|ICD9CM|Unc behav neo adrenal|Unc behav neo adrenal
C0027634|T191|PT|237.3|ICD9CM|Neoplasm of uncertain behavior of paraganglia|Neoplasm of uncertain behavior of paraganglia
C0027634|T191|AB|237.3|ICD9CM|Unc behav neo paragang|Unc behav neo paragang
C0154118|T191|PT|237.4|ICD9CM|Neoplasm of uncertain behavior of other and unspecified endocrine glands|Neoplasm of uncertain behavior of other and unspecified endocrine glands
C0154118|T191|AB|237.4|ICD9CM|Uncer neo endocrine NEC|Uncer neo endocrine NEC
C0154119|T191|PT|237.5|ICD9CM|Neoplasm of uncertain behavior of brain and spinal cord|Neoplasm of uncertain behavior of brain and spinal cord
C0154119|T191|AB|237.5|ICD9CM|Unc beh neo brain/spinal|Unc beh neo brain/spinal
C0154120|T191|PT|237.6|ICD9CM|Neoplasm of uncertain behavior of meninges|Neoplasm of uncertain behavior of meninges
C0154120|T191|AB|237.6|ICD9CM|Unc behav neo meninges|Unc behav neo meninges
C0162678|T191|HT|237.7|ICD9CM|Neurofibromatosis|Neurofibromatosis
C0162678|T191|AB|237.70|ICD9CM|Neurofibromatosis NOS|Neurofibromatosis NOS
C0162678|T191|PT|237.70|ICD9CM|Neurofibromatosis, unspecified|Neurofibromatosis, unspecified
C0027831|T191|AB|237.71|ICD9CM|Neurofibromatosis type I|Neurofibromatosis type I
C0027831|T191|PT|237.71|ICD9CM|Neurofibromatosis, type 1 [von recklinghausen's disease]|Neurofibromatosis, type 1 [von recklinghausen's disease]
C0027832|T191|AB|237.72|ICD9CM|Neurofibromatosis typ II|Neurofibromatosis typ II
C0027832|T191|PT|237.72|ICD9CM|Neurofibromatosis, type 2 [acoustic neurofibromatosis]|Neurofibromatosis, type 2 [acoustic neurofibromatosis]
C1335929|T191|PT|237.73|ICD9CM|Schwannomatosis|Schwannomatosis
C1335929|T191|AB|237.73|ICD9CM|Schwannomatosis|Schwannomatosis
C2921012|T047|AB|237.79|ICD9CM|Neurofibromatosis NEC|Neurofibromatosis NEC
C2921012|T047|PT|237.79|ICD9CM|Other neurofibromatosis|Other neurofibromatosis
C0154123|T191|PT|237.9|ICD9CM|Neoplasm of uncertain behavior of other and unspecified parts of nervous system|Neoplasm of uncertain behavior of other and unspecified parts of nervous system
C0154123|T191|AB|237.9|ICD9CM|Unc beh neo nerv sys NEC|Unc beh neo nerv sys NEC
C0154124|T191|HT|238|ICD9CM|Neoplasm of uncertain behavior of other and unspecified sites and tissues|Neoplasm of uncertain behavior of other and unspecified sites and tissues
C0027630|T191|PT|238.0|ICD9CM|Neoplasm of uncertain behavior of bone and articular cartilage|Neoplasm of uncertain behavior of bone and articular cartilage
C0027630|T191|AB|238.0|ICD9CM|Unc behav neo bone|Unc behav neo bone
C0154125|T191|PT|238.1|ICD9CM|Neoplasm of uncertain behavior of connective and other soft tissue|Neoplasm of uncertain behavior of connective and other soft tissue
C0154125|T191|AB|238.1|ICD9CM|Unc behav neo soft tissu|Unc behav neo soft tissu
C0496955|T191|PT|238.2|ICD9CM|Neoplasm of uncertain behavior of skin|Neoplasm of uncertain behavior of skin
C0496955|T191|AB|238.2|ICD9CM|Unc behav neo skin|Unc behav neo skin
C0496956|T191|PT|238.3|ICD9CM|Neoplasm of uncertain behavior of breast|Neoplasm of uncertain behavior of breast
C0496956|T191|AB|238.3|ICD9CM|Unc behav neo breast|Unc behav neo breast
C0032463|T191|AB|238.4|ICD9CM|Polycythemia vera|Polycythemia vera
C0032463|T191|PT|238.4|ICD9CM|Polycythemia vera|Polycythemia vera
C0154127|T191|AB|238.5|ICD9CM|Mastocytoma NOS|Mastocytoma NOS
C0154127|T191|PT|238.5|ICD9CM|Neoplasm of uncertain behavior of histiocytic and mast cells|Neoplasm of uncertain behavior of histiocytic and mast cells
C0027638|T191|PT|238.6|ICD9CM|Neoplasm of uncertain behavior of plasma cells|Neoplasm of uncertain behavior of plasma cells
C0027638|T191|AB|238.6|ICD9CM|Plasmacytoma NOS|Plasmacytoma NOS
C0027632|T191|HT|238.7|ICD9CM|Neoplasm of uncertain behavior of other lymphatic and hematopoietic tissues|Neoplasm of uncertain behavior of other lymphatic and hematopoietic tissues
C0040028|T047|PT|238.71|ICD9CM|Essential thrombocythemia|Essential thrombocythemia
C0040028|T047|AB|238.71|ICD9CM|Essntial thrombocythemia|Essntial thrombocythemia
C1719305|T047|PT|238.72|ICD9CM|Low grade myelodysplastic syndrome lesions|Low grade myelodysplastic syndrome lesions
C1719305|T047|AB|238.72|ICD9CM|Low grde myelody syn les|Low grde myelody syn les
C1719308|T047|AB|238.73|ICD9CM|Hi grde myelodys syn les|Hi grde myelodys syn les
C1719308|T047|PT|238.73|ICD9CM|High grade myelodysplastic syndrome lesions|High grade myelodysplastic syndrome lesions
C1292779|T191|PT|238.74|ICD9CM|Myelodysplastic syndrome with 5q deletion|Myelodysplastic syndrome with 5q deletion
C1292779|T191|AB|238.74|ICD9CM|Myelodyspls syn w 5q del|Myelodyspls syn w 5q del
C3463824|T191|AB|238.75|ICD9CM|Myelodysplastic synd NOS|Myelodysplastic synd NOS
C3463824|T191|PT|238.75|ICD9CM|Myelodysplastic syndrome, unspecified|Myelodysplastic syndrome, unspecified
C0001815|T191|AB|238.76|ICD9CM|Myelofi w myelo metaplas|Myelofi w myelo metaplas
C0001815|T191|PT|238.76|ICD9CM|Myelofibrosis with myeloid metaplasia|Myelofibrosis with myeloid metaplasia
C0432487|T191|AB|238.77|ICD9CM|Post tp lymphprolif dis|Post tp lymphprolif dis
C0432487|T191|PT|238.77|ICD9CM|Post-transplant lymphoproliferative disorder (PTLD)|Post-transplant lymphoproliferative disorder (PTLD)
C1706492|T191|AB|238.79|ICD9CM|Lymph/hematpoitc tis NEC|Lymph/hematpoitc tis NEC
C1706492|T191|PT|238.79|ICD9CM|Other lymphatic and hematopoietic tissues|Other lymphatic and hematopoietic tissues
C2873733|T191|PT|238.8|ICD9CM|Neoplasm of uncertain behavior of other specified sites|Neoplasm of uncertain behavior of other specified sites
C2873733|T191|AB|238.8|ICD9CM|Uncert behavior neo NEC|Uncert behavior neo NEC
C0375110|T191|PT|238.9|ICD9CM|Neoplasm of uncertain behavior, site unspecified|Neoplasm of uncertain behavior, site unspecified
C0375110|T191|AB|238.9|ICD9CM|Uncert behavior neo NOS|Uncert behavior neo NOS
C3665668|T191|HT|239|ICD9CM|Neoplasms of unspecified nature|Neoplasms of unspecified nature
C3665668|T191|HT|239-239.99|ICD9CM|NEOPLASMS OF UNSPECIFIED NATURE|NEOPLASMS OF UNSPECIFIED NATURE
C0012243|T191|AB|239.0|ICD9CM|Digestive neoplasm NOS|Digestive neoplasm NOS
C0012243|T191|PT|239.0|ICD9CM|Neoplasm of unspecified nature of digestive system|Neoplasm of unspecified nature of digestive system
C0154131|T191|PT|239.1|ICD9CM|Neoplasm of unspecified nature of respiratory system|Neoplasm of unspecified nature of respiratory system
C0154131|T191|AB|239.1|ICD9CM|Respiratory neoplasm NOS|Respiratory neoplasm NOS
C0154132|T191|AB|239.2|ICD9CM|Bone/skin neoplasm NOS|Bone/skin neoplasm NOS
C0154132|T191|PT|239.2|ICD9CM|Neoplasm of unspecified nature of bone, soft tissue, and skin|Neoplasm of unspecified nature of bone, soft tissue, and skin
C0027641|T191|AB|239.3|ICD9CM|Breast neoplasm NOS|Breast neoplasm NOS
C0027641|T191|PT|239.3|ICD9CM|Neoplasm of unspecified nature of breast|Neoplasm of unspecified nature of breast
C0027639|T191|AB|239.4|ICD9CM|Bladder neoplasm NOS|Bladder neoplasm NOS
C0027639|T191|PT|239.4|ICD9CM|Neoplasm of unspecified nature of bladder|Neoplasm of unspecified nature of bladder
C0154133|T191|PT|239.5|ICD9CM|Neoplasm of unspecified nature of other genitourinary organs|Neoplasm of unspecified nature of other genitourinary organs
C0154133|T191|AB|239.5|ICD9CM|Other gu neoplasm NOS|Other gu neoplasm NOS
C0006118|T191|AB|239.6|ICD9CM|Brain neoplasm NOS|Brain neoplasm NOS
C0006118|T191|PT|239.6|ICD9CM|Neoplasm of unspecified nature of brain|Neoplasm of unspecified nature of brain
C0154134|T191|AB|239.7|ICD9CM|Endocrine/nerv neo NOS|Endocrine/nerv neo NOS
C0154134|T191|PT|239.7|ICD9CM|Neoplasm of unspecified nature of endocrine glands and other parts of nervous system|Neoplasm of unspecified nature of endocrine glands and other parts of nervous system
C0154135|T191|HT|239.8|ICD9CM|Neoplasm of unspecified nature of other specified sites|Neoplasm of unspecified nature of other specified sites
C2712911|T191|AB|239.81|ICD9CM|Neo retina/choroid NOS|Neo retina/choroid NOS
C2712911|T191|PT|239.81|ICD9CM|Neoplasms of unspecified nature, retina and choroid|Neoplasms of unspecified nature, retina and choroid
C0154135|T191|AB|239.89|ICD9CM|Neoplasm other sites NOS|Neoplasm other sites NOS
C0154135|T191|PT|239.89|ICD9CM|Neoplasms of unspecified nature, other specified sites|Neoplasms of unspecified nature, other specified sites
C0375111|T191|AB|239.9|ICD9CM|Neoplasm NOS|Neoplasm NOS
C0375111|T191|PT|239.9|ICD9CM|Neoplasm of unspecified nature, site unspecified|Neoplasm of unspecified nature, site unspecified
C0037158|T047|HT|240|ICD9CM|Simple and unspecified goiter|Simple and unspecified goiter
C0040128|T047|HT|240-246.99|ICD9CM|DISORDERS OF THYROID GLAND|DISORDERS OF THYROID GLAND
C0342105|T047|HT|240-279.99|ICD9CM|ENDOCRINE, NUTRITIONAL AND METABOLIC DISEASES, AND IMMUNITY DISORDERS|ENDOCRINE, NUTRITIONAL AND METABOLIC DISEASES, AND IMMUNITY DISORDERS
C0018022|T047|PT|240.0|ICD9CM|Goiter, specified as simple|Goiter, specified as simple
C0018022|T047|AB|240.0|ICD9CM|Simple goiter|Simple goiter
C0018021|T047|AB|240.9|ICD9CM|Goiter NOS|Goiter NOS
C0018021|T047|PT|240.9|ICD9CM|Goiter, unspecified|Goiter, unspecified
C1318500|T047|HT|241|ICD9CM|Nontoxic nodular goiter|Nontoxic nodular goiter
C0342115|T047|AB|241.0|ICD9CM|Nontox uninodular goiter|Nontox uninodular goiter
C0342115|T047|PT|241.0|ICD9CM|Nontoxic uninodular goiter|Nontoxic uninodular goiter
C0271761|T047|AB|241.1|ICD9CM|Nontox multinodul goiter|Nontox multinodul goiter
C0271761|T047|PT|241.1|ICD9CM|Nontoxic multinodular goiter|Nontoxic multinodular goiter
C1318500|T047|AB|241.9|ICD9CM|Nontox nodul goiter NOS|Nontox nodul goiter NOS
C1318500|T047|PT|241.9|ICD9CM|Unspecified nontoxic nodular goiter|Unspecified nontoxic nodular goiter
C0040156|T047|HT|242|ICD9CM|Thyrotoxicosis with or without goiter|Thyrotoxicosis with or without goiter
C0342122|T047|HT|242.0|ICD9CM|Toxic diffuse goiter|Toxic diffuse goiter
C0154138|T047|AB|242.00|ICD9CM|Tox dif goiter no crisis|Tox dif goiter no crisis
C0154138|T047|PT|242.00|ICD9CM|Toxic diffuse goiter without mention of thyrotoxic crisis or storm|Toxic diffuse goiter without mention of thyrotoxic crisis or storm
C0154139|T047|AB|242.01|ICD9CM|Tox dif goiter w crisis|Tox dif goiter w crisis
C0154139|T047|PT|242.01|ICD9CM|Toxic diffuse goiter with mention of thyrotoxic crisis or storm|Toxic diffuse goiter with mention of thyrotoxic crisis or storm
C0154141|T047|HT|242.1|ICD9CM|Toxic uninodular goiter|Toxic uninodular goiter
C0489955|T047|AB|242.10|ICD9CM|Tox uninod goit no cris|Tox uninod goit no cris
C0489955|T047|PT|242.10|ICD9CM|Toxic uninodular goiter without mention of thyrotoxic crisis or storm|Toxic uninodular goiter without mention of thyrotoxic crisis or storm
C0154142|T047|AB|242.11|ICD9CM|Tox uninod goit w crisis|Tox uninod goit w crisis
C0154142|T047|PT|242.11|ICD9CM|Toxic uninodular goiter with mention of thyrotoxic crisis or storm|Toxic uninodular goiter with mention of thyrotoxic crisis or storm
C0154143|T047|HT|242.2|ICD9CM|Toxic multinodular goiter|Toxic multinodular goiter
C0154144|T047|AB|242.20|ICD9CM|Tox multnod goit no cris|Tox multnod goit no cris
C0154144|T047|PT|242.20|ICD9CM|Toxic multinodular goiter without mention of thyrotoxic crisis or storm|Toxic multinodular goiter without mention of thyrotoxic crisis or storm
C0154145|T047|AB|242.21|ICD9CM|Tox multnod goit w cris|Tox multnod goit w cris
C0154145|T047|PT|242.21|ICD9CM|Toxic multinodular goiter with mention of thyrotoxic crisis or storm|Toxic multinodular goiter with mention of thyrotoxic crisis or storm
C0342127|T047|HT|242.3|ICD9CM|Toxic nodular goiter, unspecified type|Toxic nodular goiter, unspecified type
C0154146|T047|AB|242.30|ICD9CM|Tox nod goiter no crisis|Tox nod goiter no crisis
C0154146|T047|PT|242.30|ICD9CM|Toxic nodular goiter, unspecified type, without mention of thyrotoxic crisis or storm|Toxic nodular goiter, unspecified type, without mention of thyrotoxic crisis or storm
C0154147|T047|AB|242.31|ICD9CM|Tox nod goiter w crisis|Tox nod goiter w crisis
C0154147|T047|PT|242.31|ICD9CM|Toxic nodular goiter, unspecified type, with mention of thyrotoxic crisis or storm|Toxic nodular goiter, unspecified type, with mention of thyrotoxic crisis or storm
C0154148|T047|HT|242.4|ICD9CM|Thyrotoxicosis from ectopic thyroid nodule|Thyrotoxicosis from ectopic thyroid nodule
C0342132|T047|AB|242.40|ICD9CM|Thyrotox-ect nod no cris|Thyrotox-ect nod no cris
C0342132|T047|PT|242.40|ICD9CM|Thyrotoxicosis from ectopic thyroid nodule without mention of thyrotoxic crisis or storm|Thyrotoxicosis from ectopic thyroid nodule without mention of thyrotoxic crisis or storm
C0342133|T047|AB|242.41|ICD9CM|Thyrotox-ect nod w cris|Thyrotox-ect nod w cris
C0342133|T047|PT|242.41|ICD9CM|Thyrotoxicosis from ectopic thyroid nodule with mention of thyrotoxic crisis or storm|Thyrotoxicosis from ectopic thyroid nodule with mention of thyrotoxic crisis or storm
C0154151|T047|HT|242.8|ICD9CM|Thyrotoxicosis of other specified origin|Thyrotoxicosis of other specified origin
C0154152|T047|PT|242.80|ICD9CM|Thyrotoxicosis of other specified origin without mention of thyrotoxic crisis or storm|Thyrotoxicosis of other specified origin without mention of thyrotoxic crisis or storm
C0154152|T047|AB|242.80|ICD9CM|Thyrtox orig NEC no cris|Thyrtox orig NEC no cris
C0154153|T047|AB|242.81|ICD9CM|Thyrotox orig NEC w cris|Thyrotox orig NEC w cris
C0154153|T047|PT|242.81|ICD9CM|Thyrotoxicosis of other specified origin with mention of thyrotoxic crisis or storm|Thyrotoxicosis of other specified origin with mention of thyrotoxic crisis or storm
C0271763|T047|HT|242.9|ICD9CM|Thyrotoxicosis without mention of goiter or other cause|Thyrotoxicosis without mention of goiter or other cause
C0154154|T047|AB|242.90|ICD9CM|Thyrotox NOS no crisis|Thyrotox NOS no crisis
C0154155|T047|AB|242.91|ICD9CM|Thyrotox NOS w crisis|Thyrotox NOS w crisis
C0154155|T047|PT|242.91|ICD9CM|Thyrotoxicosis without mention of goiter or other cause, with mention of thyrotoxic crisis or storm|Thyrotoxicosis without mention of goiter or other cause, with mention of thyrotoxic crisis or storm
C0010308|T047|PT|243|ICD9CM|Congenital hypothyroidism|Congenital hypothyroidism
C0010308|T047|AB|243|ICD9CM|Congenital hypothyroidsm|Congenital hypothyroidsm
C0700502|T047|HT|244|ICD9CM|Acquired hypothyroidism|Acquired hypothyroidism
C0154157|T047|AB|244.0|ICD9CM|Postsurgical hypothyroid|Postsurgical hypothyroid
C0154157|T047|PT|244.0|ICD9CM|Postsurgical hypothyroidism|Postsurgical hypothyroidism
C0154158|T047|PT|244.1|ICD9CM|Other postablative hypothyroidism|Other postablative hypothyroidism
C0154158|T047|AB|244.1|ICD9CM|Postablat hypothyr NEC|Postablat hypothyr NEC
C0154159|T047|AB|244.2|ICD9CM|Iodine hypothyroidism|Iodine hypothyroidism
C0154159|T047|PT|244.2|ICD9CM|Iodine hypothyroidism|Iodine hypothyroidism
C0154160|T047|AB|244.3|ICD9CM|Iatrogen hypothyroid NEC|Iatrogen hypothyroid NEC
C0154160|T047|PT|244.3|ICD9CM|Other iatrogenic hypothyroidism|Other iatrogenic hypothyroidism
C0154161|T047|AB|244.8|ICD9CM|Acquired hypothyroid NEC|Acquired hypothyroid NEC
C0154161|T047|PT|244.8|ICD9CM|Other specified acquired hypothyroidism|Other specified acquired hypothyroidism
C0020676|T047|AB|244.9|ICD9CM|Hypothyroidism NOS|Hypothyroidism NOS
C0020676|T047|PT|244.9|ICD9CM|Unspecified acquired hypothyroidism|Unspecified acquired hypothyroidism
C0040147|T047|HT|245|ICD9CM|Thyroiditis|Thyroiditis
C0001360|T047|AB|245.0|ICD9CM|Acute thyroiditis|Acute thyroiditis
C0001360|T047|PT|245.0|ICD9CM|Acute thyroiditis|Acute thyroiditis
C0040149|T047|AB|245.1|ICD9CM|Subacute thyroiditis|Subacute thyroiditis
C0040149|T047|PT|245.1|ICD9CM|Subacute thyroiditis|Subacute thyroiditis
C0677607|T047|AB|245.2|ICD9CM|Chr lymphocyt thyroidit|Chr lymphocyt thyroidit
C0677607|T047|PT|245.2|ICD9CM|Chronic lymphocytic thyroiditis|Chronic lymphocytic thyroiditis
C3887878|T047|AB|245.3|ICD9CM|Chr fibrous thyroiditis|Chr fibrous thyroiditis
C3887878|T047|PT|245.3|ICD9CM|Chronic fibrous thyroiditis|Chronic fibrous thyroiditis
C0154163|T047|AB|245.4|ICD9CM|Iatrogenic thyroiditis|Iatrogenic thyroiditis
C0154163|T047|PT|245.4|ICD9CM|Iatrogenic thyroiditis|Iatrogenic thyroiditis
C0029495|T047|AB|245.8|ICD9CM|Chr thyroiditis NEC/NOS|Chr thyroiditis NEC/NOS
C0029495|T047|PT|245.8|ICD9CM|Other and unspecified chronic thyroiditis|Other and unspecified chronic thyroiditis
C0040147|T047|AB|245.9|ICD9CM|Thyroiditis NOS|Thyroiditis NOS
C0040147|T047|PT|245.9|ICD9CM|Thyroiditis, unspecified|Thyroiditis, unspecified
C0154164|T047|HT|246|ICD9CM|Other disorders of thyroid|Other disorders of thyroid
C0701822|T047|AB|246.0|ICD9CM|Dis thyrocalciton secret|Dis thyrocalciton secret
C0701822|T047|PT|246.0|ICD9CM|Disorders of thyrocalcitonin secretion|Disorders of thyrocalcitonin secretion
C0152077|T047|AB|246.1|ICD9CM|Dyshormonogenic goiter|Dyshormonogenic goiter
C0152077|T047|PT|246.1|ICD9CM|Dyshormonogenic goiter|Dyshormonogenic goiter
C0162299|T047|AB|246.2|ICD9CM|Cyst of thyroid|Cyst of thyroid
C0162299|T047|PT|246.2|ICD9CM|Cyst of thyroid|Cyst of thyroid
C0154166|T046|AB|246.3|ICD9CM|Hemorr/infarc thyroid|Hemorr/infarc thyroid
C0154166|T046|PT|246.3|ICD9CM|Hemorrhage and infarction of thyroid|Hemorrhage and infarction of thyroid
C0154167|T047|AB|246.8|ICD9CM|Disorders of thyroid NEC|Disorders of thyroid NEC
C0154167|T047|PT|246.8|ICD9CM|Other specified disorders of thyroid|Other specified disorders of thyroid
C0040128|T047|AB|246.9|ICD9CM|Disorder of thyroid NOS|Disorder of thyroid NOS
C0040128|T047|PT|246.9|ICD9CM|Unspecified disorder of thyroid|Unspecified disorder of thyroid
C0271640|T047|HT|249|ICD9CM|Secondary diabetes mellitus|Secondary diabetes mellitus
C0178257|T047|HT|249-259.99|ICD9CM|DISEASES OF OTHER ENDOCRINE GLANDS|DISEASES OF OTHER ENDOCRINE GLANDS
C2349363|T047|HT|249.0|ICD9CM|Secondary diabetes mellitus, without mention of complication|Secondary diabetes mellitus, without mention of complication
C2349361|T047|AB|249.00|ICD9CM|Sec DM wo cmp nt st uncn|Sec DM wo cmp nt st uncn
C2349362|T047|AB|249.01|ICD9CM|Sec DM wo comp uncontrld|Sec DM wo comp uncontrld
C2349362|T047|PT|249.01|ICD9CM|Secondary diabetes mellitus without mention of complication, uncontrolled|Secondary diabetes mellitus without mention of complication, uncontrolled
C2349367|T047|HT|249.1|ICD9CM|Secondary diabetes mellitus with ketoacidosis|Secondary diabetes mellitus with ketoacidosis
C2349365|T047|AB|249.10|ICD9CM|Sec DM keto nt st uncntr|Sec DM keto nt st uncntr
C2349365|T047|PT|249.10|ICD9CM|Secondary diabetes mellitus with ketoacidosis, not stated as uncontrolled, or unspecified|Secondary diabetes mellitus with ketoacidosis, not stated as uncontrolled, or unspecified
C2349366|T047|AB|249.11|ICD9CM|Sec DM ketoacd uncntrld|Sec DM ketoacd uncntrld
C2349366|T047|PT|249.11|ICD9CM|Secondary diabetes mellitus with ketoacidosis, uncontrolled|Secondary diabetes mellitus with ketoacidosis, uncontrolled
C2349372|T047|HT|249.2|ICD9CM|Secondary diabetes mellitus with hyperosmolarity|Secondary diabetes mellitus with hyperosmolarity
C2349370|T047|AB|249.20|ICD9CM|Sec DM hpros nt st uncnr|Sec DM hpros nt st uncnr
C2349370|T047|PT|249.20|ICD9CM|Secondary diabetes mellitus with hyperosmolarity, not stated as uncontrolled, or unspecified|Secondary diabetes mellitus with hyperosmolarity, not stated as uncontrolled, or unspecified
C2349371|T047|AB|249.21|ICD9CM|Sec DM hprosmlr uncntrld|Sec DM hprosmlr uncntrld
C2349371|T047|PT|249.21|ICD9CM|Secondary diabetes mellitus with hyperosmolarity, uncontrolled|Secondary diabetes mellitus with hyperosmolarity, uncontrolled
C2349376|T047|HT|249.3|ICD9CM|Secondary diabetes mellitus with other coma|Secondary diabetes mellitus with other coma
C2349374|T047|AB|249.30|ICD9CM|Sec DM ot cma nt st uncn|Sec DM ot cma nt st uncn
C2349374|T047|PT|249.30|ICD9CM|Secondary diabetes mellitus with other coma, not stated as uncontrolled, or unspecified|Secondary diabetes mellitus with other coma, not stated as uncontrolled, or unspecified
C2349375|T047|AB|249.31|ICD9CM|Sec DM oth coma uncntrld|Sec DM oth coma uncntrld
C2349375|T047|PT|249.31|ICD9CM|Secondary diabetes mellitus with other coma, uncontrolled|Secondary diabetes mellitus with other coma, uncontrolled
C2349382|T047|HT|249.4|ICD9CM|Secondary diabetes mellitus with renal manifestations|Secondary diabetes mellitus with renal manifestations
C2349380|T047|AB|249.40|ICD9CM|Sec DM renl nt st uncntr|Sec DM renl nt st uncntr
C2349380|T047|PT|249.40|ICD9CM|Secondary diabetes mellitus with renal manifestations, not stated as uncontrolled, or unspecified|Secondary diabetes mellitus with renal manifestations, not stated as uncontrolled, or unspecified
C2349381|T047|AB|249.41|ICD9CM|Sec DM renal uncontrld|Sec DM renal uncontrld
C2349381|T047|PT|249.41|ICD9CM|Secondary diabetes mellitus with renal manifestations, uncontrolled|Secondary diabetes mellitus with renal manifestations, uncontrolled
C2349385|T047|HT|249.5|ICD9CM|Secondary diabetes mellitus with ophthalmic manifestations|Secondary diabetes mellitus with ophthalmic manifestations
C2349383|T047|AB|249.50|ICD9CM|Sec DM ophth nt st uncn|Sec DM ophth nt st uncn
C2349384|T047|AB|249.51|ICD9CM|Sec DM ophth uncontrld|Sec DM ophth uncontrld
C2349384|T047|PT|249.51|ICD9CM|Secondary diabetes mellitus with ophthalmic manifestations, uncontrolled|Secondary diabetes mellitus with ophthalmic manifestations, uncontrolled
C2349388|T047|HT|249.6|ICD9CM|Secondary diabetes mellitus with neurological manifestations|Secondary diabetes mellitus with neurological manifestations
C2349386|T047|AB|249.60|ICD9CM|Sec DM neuro nt st uncn|Sec DM neuro nt st uncn
C2349387|T047|AB|249.61|ICD9CM|Sec DM neuro uncontrld|Sec DM neuro uncontrld
C2349387|T047|PT|249.61|ICD9CM|Secondary diabetes mellitus with neurological manifestations, uncontrolled|Secondary diabetes mellitus with neurological manifestations, uncontrolled
C2349391|T047|HT|249.7|ICD9CM|Secondary diabetes mellitus with peripheral circulatory disorders|Secondary diabetes mellitus with peripheral circulatory disorders
C2349389|T047|AB|249.70|ICD9CM|Sec DM circ nt st uncntr|Sec DM circ nt st uncntr
C2349390|T047|AB|249.71|ICD9CM|Sec DM circ uncontrld|Sec DM circ uncontrld
C2349390|T047|PT|249.71|ICD9CM|Secondary diabetes mellitus with peripheral circulatory disorders, uncontrolled|Secondary diabetes mellitus with peripheral circulatory disorders, uncontrolled
C2349394|T047|HT|249.8|ICD9CM|Secondary diabetes mellitus with other specified manifestations|Secondary diabetes mellitus with other specified manifestations
C2349392|T047|AB|249.80|ICD9CM|Sec DM oth nt st uncontr|Sec DM oth nt st uncontr
C2349393|T047|AB|249.81|ICD9CM|Sec DM other uncontrld|Sec DM other uncontrld
C2349393|T047|PT|249.81|ICD9CM|Secondary diabetes mellitus with other specified manifestations, uncontrolled|Secondary diabetes mellitus with other specified manifestations, uncontrolled
C2349399|T047|HT|249.9|ICD9CM|Secondary diabetes mellitus with unspecified complication|Secondary diabetes mellitus with unspecified complication
C2349397|T047|AB|249.90|ICD9CM|Sec DM unsp nt st uncon|Sec DM unsp nt st uncon
C2349398|T047|AB|249.91|ICD9CM|Sec DM unsp uncontrold|Sec DM unsp uncontrold
C2349398|T047|PT|249.91|ICD9CM|Secondary diabetes mellitus with unspecified complication, uncontrolled|Secondary diabetes mellitus with unspecified complication, uncontrolled
C0011849|T047|HT|250|ICD9CM|Diabetes mellitus|Diabetes mellitus
C0271635|T047|HT|250.0|ICD9CM|Diabetes mellitus without mention of complication|Diabetes mellitus without mention of complication
C0375113|T047|AB|250.00|ICD9CM|DMII wo cmp nt st uncntr|DMII wo cmp nt st uncntr
C0375114|T047|AB|250.01|ICD9CM|DMI wo cmp nt st uncntrl|DMI wo cmp nt st uncntrl
C0375115|T047|PT|250.02|ICD9CM|Diabetes mellitus without mention of complication, type II or unspecified type, uncontrolled|Diabetes mellitus without mention of complication, type II or unspecified type, uncontrolled
C0375115|T047|AB|250.02|ICD9CM|DMII wo cmp uncntrld|DMII wo cmp uncntrld
C0375116|T047|PT|250.03|ICD9CM|Diabetes mellitus without mention of complication, type I [juvenile type], uncontrolled|Diabetes mellitus without mention of complication, type I [juvenile type], uncontrolled
C0375116|T047|AB|250.03|ICD9CM|DMI wo cmp uncntrld|DMI wo cmp uncntrld
C0011880|T047|HT|250.1|ICD9CM|Diabetes with ketoacidosis|Diabetes with ketoacidosis
C0375117|T047|PT|250.10|ICD9CM|Diabetes with ketoacidosis, type II or unspecified type, not stated as uncontrolled|Diabetes with ketoacidosis, type II or unspecified type, not stated as uncontrolled
C0375117|T047|AB|250.10|ICD9CM|DMII keto nt st uncntrld|DMII keto nt st uncntrld
C0375118|T047|PT|250.11|ICD9CM|Diabetes with ketoacidosis, type I [juvenile type], not stated as uncontrolled|Diabetes with ketoacidosis, type I [juvenile type], not stated as uncontrolled
C0375118|T047|AB|250.11|ICD9CM|DMI keto nt st uncntrld|DMI keto nt st uncntrld
C0375119|T047|PT|250.12|ICD9CM|Diabetes with ketoacidosis, type II or unspecified type, uncontrolled|Diabetes with ketoacidosis, type II or unspecified type, uncontrolled
C0375119|T047|AB|250.12|ICD9CM|DMII ketoacd uncontrold|DMII ketoacd uncontrold
C0375120|T047|PT|250.13|ICD9CM|Diabetes with ketoacidosis, type I [juvenile type], uncontrolled|Diabetes with ketoacidosis, type I [juvenile type], uncontrolled
C0375120|T047|AB|250.13|ICD9CM|DMI ketoacd uncontrold|DMI ketoacd uncontrold
C0375121|T047|HT|250.2|ICD9CM|Diabetes mellitus with hyperosmolarity|Diabetes mellitus with hyperosmolarity
C0375122|T047|PT|250.20|ICD9CM|Diabetes with hyperosmolarity, type II or unspecified type, not stated as uncontrolled|Diabetes with hyperosmolarity, type II or unspecified type, not stated as uncontrolled
C0375122|T047|AB|250.20|ICD9CM|DMII hprsm nt st uncntrl|DMII hprsm nt st uncntrl
C0375123|T047|PT|250.21|ICD9CM|Diabetes with hyperosmolarity, type I [juvenile type], not stated as uncontrolled|Diabetes with hyperosmolarity, type I [juvenile type], not stated as uncontrolled
C0375123|T047|AB|250.21|ICD9CM|DMI hprsm nt st uncntrld|DMI hprsm nt st uncntrld
C0375124|T047|PT|250.22|ICD9CM|Diabetes with hyperosmolarity, type II or unspecified type, uncontrolled|Diabetes with hyperosmolarity, type II or unspecified type, uncontrolled
C0375124|T047|AB|250.22|ICD9CM|DMII hprosmlr uncontrold|DMII hprosmlr uncontrold
C0375125|T047|PT|250.23|ICD9CM|Diabetes with hyperosmolarity, type I [juvenile type], uncontrolled|Diabetes with hyperosmolarity, type I [juvenile type], uncontrolled
C0375125|T047|AB|250.23|ICD9CM|DMI hprosmlr uncontrold|DMI hprosmlr uncontrold
C0011870|T047|HT|250.3|ICD9CM|Diabetes with other coma|Diabetes with other coma
C0375126|T047|PT|250.30|ICD9CM|Diabetes with other coma, type II or unspecified type, not stated as uncontrolled|Diabetes with other coma, type II or unspecified type, not stated as uncontrolled
C0375126|T047|AB|250.30|ICD9CM|DMII o cm nt st uncntrld|DMII o cm nt st uncntrld
C0375127|T047|PT|250.31|ICD9CM|Diabetes with other coma, type I [juvenile type], not stated as uncontrolled|Diabetes with other coma, type I [juvenile type], not stated as uncontrolled
C0375127|T047|AB|250.31|ICD9CM|DMI o cm nt st uncntrld|DMI o cm nt st uncntrld
C0375128|T047|PT|250.32|ICD9CM|Diabetes with other coma, type II or unspecified type, uncontrolled|Diabetes with other coma, type II or unspecified type, uncontrolled
C0375128|T047|AB|250.32|ICD9CM|DMII oth coma uncontrold|DMII oth coma uncontrold
C0375129|T047|PT|250.33|ICD9CM|Diabetes with other coma, type I [juvenile type], uncontrolled|Diabetes with other coma, type I [juvenile type], uncontrolled
C0375129|T047|AB|250.33|ICD9CM|DMI oth coma uncontrold|DMI oth coma uncontrold
C0011881|T047|HT|250.4|ICD9CM|Diabetes with renal manifestations|Diabetes with renal manifestations
C0375130|T047|PT|250.40|ICD9CM|Diabetes with renal manifestations, type II or unspecified type, not stated as uncontrolled|Diabetes with renal manifestations, type II or unspecified type, not stated as uncontrolled
C0375130|T047|AB|250.40|ICD9CM|DMII renl nt st uncntrld|DMII renl nt st uncntrld
C0375131|T047|PT|250.41|ICD9CM|Diabetes with renal manifestations, type I [juvenile type], not stated as uncontrolled|Diabetes with renal manifestations, type I [juvenile type], not stated as uncontrolled
C0375131|T047|AB|250.41|ICD9CM|DMI renl nt st uncntrld|DMI renl nt st uncntrld
C0375132|T047|PT|250.42|ICD9CM|Diabetes with renal manifestations, type II or unspecified type, uncontrolled|Diabetes with renal manifestations, type II or unspecified type, uncontrolled
C0375132|T047|AB|250.42|ICD9CM|DMII renal uncntrld|DMII renal uncntrld
C0375133|T047|PT|250.43|ICD9CM|Diabetes with renal manifestations, type I [juvenile type], uncontrolled|Diabetes with renal manifestations, type I [juvenile type], uncontrolled
C0375133|T047|AB|250.43|ICD9CM|DMI renal uncntrld|DMI renal uncntrld
C0342245|T047|HT|250.5|ICD9CM|Diabetes with ophthalmic manifestations|Diabetes with ophthalmic manifestations
C0375134|T047|PT|250.50|ICD9CM|Diabetes with ophthalmic manifestations, type II or unspecified type, not stated as uncontrolled|Diabetes with ophthalmic manifestations, type II or unspecified type, not stated as uncontrolled
C0375134|T047|AB|250.50|ICD9CM|DMII ophth nt st uncntrl|DMII ophth nt st uncntrl
C0375135|T047|PT|250.51|ICD9CM|Diabetes with ophthalmic manifestations, type I [juvenile type], not stated as uncontrolled|Diabetes with ophthalmic manifestations, type I [juvenile type], not stated as uncontrolled
C0375135|T047|AB|250.51|ICD9CM|DMI ophth nt st uncntrld|DMI ophth nt st uncntrld
C0376128|T047|PT|250.52|ICD9CM|Diabetes with ophthalmic manifestations, type II or unspecified type, uncontrolled|Diabetes with ophthalmic manifestations, type II or unspecified type, uncontrolled
C0376128|T047|AB|250.52|ICD9CM|DMII ophth uncntrld|DMII ophth uncntrld
C0375136|T047|PT|250.53|ICD9CM|Diabetes with ophthalmic manifestations, type I [juvenile type], uncontrolled|Diabetes with ophthalmic manifestations, type I [juvenile type], uncontrolled
C0375136|T047|AB|250.53|ICD9CM|DMI ophth uncntrld|DMI ophth uncntrld
C0011882|T047|HT|250.6|ICD9CM|Diabetes with neurological manifestations|Diabetes with neurological manifestations
C0375137|T047|PT|250.60|ICD9CM|Diabetes with neurological manifestations, type II or unspecified type, not stated as uncontrolled|Diabetes with neurological manifestations, type II or unspecified type, not stated as uncontrolled
C0375137|T047|AB|250.60|ICD9CM|DMII neuro nt st uncntrl|DMII neuro nt st uncntrl
C0375138|T047|PT|250.61|ICD9CM|Diabetes with neurological manifestations, type I [juvenile type], not stated as uncontrolled|Diabetes with neurological manifestations, type I [juvenile type], not stated as uncontrolled
C0375138|T047|AB|250.61|ICD9CM|DMI neuro nt st uncntrld|DMI neuro nt st uncntrld
C0375139|T047|PT|250.62|ICD9CM|Diabetes with neurological manifestations, type II or unspecified type, uncontrolled|Diabetes with neurological manifestations, type II or unspecified type, uncontrolled
C0375139|T047|AB|250.62|ICD9CM|DMII neuro uncntrld|DMII neuro uncntrld
C0375140|T047|PT|250.63|ICD9CM|Diabetes with neurological manifestations, type I [juvenile type], uncontrolled|Diabetes with neurological manifestations, type I [juvenile type], uncontrolled
C0375140|T047|AB|250.63|ICD9CM|DMI neuro uncntrld|DMI neuro uncntrld
C0011871|T047|HT|250.7|ICD9CM|Diabetes with peripheral circulatory disorders|Diabetes with peripheral circulatory disorders
C0375141|T047|AB|250.70|ICD9CM|DMII circ nt st uncntrld|DMII circ nt st uncntrld
C0375142|T047|PT|250.71|ICD9CM|Diabetes with peripheral circulatory disorders, type I [juvenile type], not stated as uncontrolled|Diabetes with peripheral circulatory disorders, type I [juvenile type], not stated as uncontrolled
C0375142|T047|AB|250.71|ICD9CM|DMI circ nt st uncntrld|DMI circ nt st uncntrld
C0375143|T047|PT|250.72|ICD9CM|Diabetes with peripheral circulatory disorders, type II or unspecified type, uncontrolled|Diabetes with peripheral circulatory disorders, type II or unspecified type, uncontrolled
C0375143|T047|AB|250.72|ICD9CM|DMII circ uncntrld|DMII circ uncntrld
C0375144|T047|PT|250.73|ICD9CM|Diabetes with peripheral circulatory disorders, type I [juvenile type], uncontrolled|Diabetes with peripheral circulatory disorders, type I [juvenile type], uncontrolled
C0375144|T047|AB|250.73|ICD9CM|DMI circ uncntrld|DMI circ uncntrld
C0154183|T047|HT|250.8|ICD9CM|Diabetes with other specified manifestations|Diabetes with other specified manifestations
C0375145|T047|AB|250.80|ICD9CM|DMII oth nt st uncntrld|DMII oth nt st uncntrld
C0375146|T047|PT|250.81|ICD9CM|Diabetes with other specified manifestations, type I [juvenile type], not stated as uncontrolled|Diabetes with other specified manifestations, type I [juvenile type], not stated as uncontrolled
C0375146|T047|AB|250.81|ICD9CM|DMI oth nt st uncntrld|DMI oth nt st uncntrld
C0375147|T047|PT|250.82|ICD9CM|Diabetes with other specified manifestations, type II or unspecified type, uncontrolled|Diabetes with other specified manifestations, type II or unspecified type, uncontrolled
C0375147|T047|AB|250.82|ICD9CM|DMII oth uncntrld|DMII oth uncntrld
C0375148|T047|PT|250.83|ICD9CM|Diabetes with other specified manifestations, type I [juvenile type], uncontrolled|Diabetes with other specified manifestations, type I [juvenile type], uncontrolled
C0375148|T047|AB|250.83|ICD9CM|DMI oth uncntrld|DMI oth uncntrld
C0342257|T047|HT|250.9|ICD9CM|Diabetes with unspecified complication|Diabetes with unspecified complication
C0375149|T047|PT|250.90|ICD9CM|Diabetes with unspecified complication, type II or unspecified type, not stated as uncontrolled|Diabetes with unspecified complication, type II or unspecified type, not stated as uncontrolled
C0375149|T047|AB|250.90|ICD9CM|DMII unspf nt st uncntrl|DMII unspf nt st uncntrl
C0375150|T047|PT|250.91|ICD9CM|Diabetes with unspecified complication, type I [juvenile type], not stated as uncontrolled|Diabetes with unspecified complication, type I [juvenile type], not stated as uncontrolled
C0375150|T047|AB|250.91|ICD9CM|DMI unspf nt st uncntrld|DMI unspf nt st uncntrld
C0375151|T047|PT|250.92|ICD9CM|Diabetes with unspecified complication, type II or unspecified type, uncontrolled|Diabetes with unspecified complication, type II or unspecified type, uncontrolled
C0375151|T047|AB|250.92|ICD9CM|DMII unspf uncntrld|DMII unspf uncntrld
C0375152|T047|PT|250.93|ICD9CM|Diabetes with unspecified complication, type I [juvenile type], uncontrolled|Diabetes with unspecified complication, type I [juvenile type], uncontrolled
C0375152|T047|AB|250.93|ICD9CM|DMI unspf uncntrld|DMI unspf uncntrld
C0154189|T047|HT|251|ICD9CM|Other disorders of pancreatic internal secretion|Other disorders of pancreatic internal secretion
C0020617|T047|AB|251.0|ICD9CM|Hypoglycemic coma|Hypoglycemic coma
C0020617|T047|PT|251.0|ICD9CM|Hypoglycemic coma|Hypoglycemic coma
C0375153|T047|AB|251.1|ICD9CM|Oth spcf hypoglycemia|Oth spcf hypoglycemia
C0375153|T047|PT|251.1|ICD9CM|Other specified hypoglycemia|Other specified hypoglycemia
C0020615|T047|AB|251.2|ICD9CM|Hypoglycemia NOS|Hypoglycemia NOS
C0020615|T047|PT|251.2|ICD9CM|Hypoglycemia, unspecified|Hypoglycemia, unspecified
C0154190|T047|AB|251.3|ICD9CM|Postsurg hypoinsulinemia|Postsurg hypoinsulinemia
C0154190|T047|PT|251.3|ICD9CM|Postsurgical hypoinsulinemia|Postsurgical hypoinsulinemia
C0154191|T047|AB|251.4|ICD9CM|Abn secretion glucagon|Abn secretion glucagon
C0154191|T047|PT|251.4|ICD9CM|Abnormality of secretion of glucagon|Abnormality of secretion of glucagon
C0000774|T047|AB|251.5|ICD9CM|Abnorm secretion gastrin|Abnorm secretion gastrin
C0000774|T047|PT|251.5|ICD9CM|Abnormality of secretion of gastrin|Abnormality of secretion of gastrin
C0154192|T047|PT|251.8|ICD9CM|Other specified disorders of pancreatic internal secretion|Other specified disorders of pancreatic internal secretion
C0154192|T047|AB|251.8|ICD9CM|Pancreatic disorder NEC|Pancreatic disorder NEC
C1263961|T047|AB|251.9|ICD9CM|Pancreatic disorder NOS|Pancreatic disorder NOS
C1263961|T047|PT|251.9|ICD9CM|Unspecified disorder of pancreatic internal secretion|Unspecified disorder of pancreatic internal secretion
C0030517|T047|HT|252|ICD9CM|Disorders of parathyroid gland|Disorders of parathyroid gland
C0020502|T047|HT|252.0|ICD9CM|Hyperparathyroidism|Hyperparathyroidism
C0020502|T047|AB|252.00|ICD9CM|Hyperparathyroidism NOS|Hyperparathyroidism NOS
C0020502|T047|PT|252.00|ICD9CM|Hyperparathyroidism, unspecified|Hyperparathyroidism, unspecified
C0221002|T047|AB|252.01|ICD9CM|Primary hyperparathyroid|Primary hyperparathyroid
C0221002|T047|PT|252.01|ICD9CM|Primary hyperparathyroidism|Primary hyperparathyroidism
C1456268|T047|AB|252.02|ICD9CM|Sec hyprprthyrd nonrenal|Sec hyprprthyrd nonrenal
C1456268|T047|PT|252.02|ICD9CM|Secondary hyperparathyroidism, non-renal|Secondary hyperparathyroidism, non-renal
C0348455|T047|AB|252.08|ICD9CM|Hyperparathyroidism NEC|Hyperparathyroidism NEC
C0348455|T047|PT|252.08|ICD9CM|Other hyperparathyroidism|Other hyperparathyroidism
C0020626|T047|AB|252.1|ICD9CM|Hypoparathyroidism|Hypoparathyroidism
C0020626|T047|PT|252.1|ICD9CM|Hypoparathyroidism|Hypoparathyroidism
C0154195|T047|PT|252.8|ICD9CM|Other specified disorders of parathyroid gland|Other specified disorders of parathyroid gland
C0154195|T047|AB|252.8|ICD9CM|Parathyroid disorder NEC|Parathyroid disorder NEC
C0030517|T047|AB|252.9|ICD9CM|Parathyroid disorder NOS|Parathyroid disorder NOS
C0030517|T047|PT|252.9|ICD9CM|Unspecified disorder of parathyroid gland|Unspecified disorder of parathyroid gland
C0859058|T047|HT|253|ICD9CM|Disorders of the pituitary gland and its hypothalamic control|Disorders of the pituitary gland and its hypothalamic control
C0405578|T047|AB|253.0|ICD9CM|Acromegaly and gigantism|Acromegaly and gigantism
C0405578|T047|PT|253.0|ICD9CM|Acromegaly and gigantism|Acromegaly and gigantism
C0029493|T047|AB|253.1|ICD9CM|Ant pituit hyperfunc NEC|Ant pituit hyperfunc NEC
C0029493|T047|PT|253.1|ICD9CM|Other and unspecified anterior pituitary hyperfunction|Other and unspecified anterior pituitary hyperfunction
C0242343|T047|AB|253.2|ICD9CM|Panhypopituitarism|Panhypopituitarism
C0242343|T047|PT|253.2|ICD9CM|Panhypopituitarism|Panhypopituitarism
C0013338|T047|AB|253.3|ICD9CM|Pituitary dwarfism|Pituitary dwarfism
C0013338|T047|PT|253.3|ICD9CM|Pituitary dwarfism|Pituitary dwarfism
C0701162|T047|AB|253.4|ICD9CM|Anter pituitary dis NEC|Anter pituitary dis NEC
C0701162|T047|PT|253.4|ICD9CM|Other anterior pituitary disorders|Other anterior pituitary disorders
C0011848|T047|AB|253.5|ICD9CM|Diabetes insipidus|Diabetes insipidus
C0011848|T047|PT|253.5|ICD9CM|Diabetes insipidus|Diabetes insipidus
C0029593|T047|AB|253.6|ICD9CM|Neurohypophysis dis NEC|Neurohypophysis dis NEC
C0029593|T047|PT|253.6|ICD9CM|Other disorders of neurohypophysis|Other disorders of neurohypophysis
C0154198|T047|AB|253.7|ICD9CM|Iatrogenic pituitary dis|Iatrogenic pituitary dis
C0154198|T047|PT|253.7|ICD9CM|Iatrogenic pituitary disorders|Iatrogenic pituitary disorders
C0029597|T047|PT|253.8|ICD9CM|Other disorders of the pituitary and other syndromes of diencephalohypophyseal origin|Other disorders of the pituitary and other syndromes of diencephalohypophyseal origin
C0029597|T047|AB|253.8|ICD9CM|Pituitary disorder NEC|Pituitary disorder NEC
C0859058|T047|AB|253.9|ICD9CM|Pituitary disorder NOS|Pituitary disorder NOS
C0859058|T047|PT|253.9|ICD9CM|Unspecified disorder of the pituitary gland and its hypothalamic control|Unspecified disorder of the pituitary gland and its hypothalamic control
C0154199|T047|HT|254|ICD9CM|Diseases of thymus gland|Diseases of thymus gland
C3887666|T047|AB|254.0|ICD9CM|Persist hyperplas thymus|Persist hyperplas thymus
C3887666|T047|PT|254.0|ICD9CM|Persistent hyperplasia of thymus|Persistent hyperplasia of thymus
C0154200|T047|AB|254.1|ICD9CM|Abscess of thymus|Abscess of thymus
C0154200|T047|PT|254.1|ICD9CM|Abscess of thymus|Abscess of thymus
C0342565|T047|AB|254.8|ICD9CM|Diseases of thymus NEC|Diseases of thymus NEC
C0342565|T047|PT|254.8|ICD9CM|Other specified diseases of thymus gland|Other specified diseases of thymus gland
C0154199|T047|AB|254.9|ICD9CM|Disease of thymus NOS|Disease of thymus NOS
C0154199|T047|PT|254.9|ICD9CM|Unspecified disease of thymus gland|Unspecified disease of thymus gland
C0001621|T047|HT|255|ICD9CM|Disorders of adrenal glands|Disorders of adrenal glands
C0010481|T047|AB|255.0|ICD9CM|Cushing's syndrome|Cushing's syndrome
C0010481|T047|PT|255.0|ICD9CM|Cushing's syndrome|Cushing's syndrome
C0020428|T047|HT|255.1|ICD9CM|Hyperaldosteronism|Hyperaldosteronism
C0020428|T047|AB|255.10|ICD9CM|Hyperaldosteronism NOS|Hyperaldosteronism NOS
C0020428|T047|PT|255.10|ICD9CM|Hyperaldosteronism, unspecified|Hyperaldosteronism, unspecified
C1260386|T047|PT|255.11|ICD9CM|Glucocorticoid-remediable aldosteronism|Glucocorticoid-remediable aldosteronism
C1260386|T047|AB|255.11|ICD9CM|Glucrtcod-rem aldsternsm|Glucrtcod-rem aldsternsm
C1384514|T047|AB|255.12|ICD9CM|Conn's syndrome|Conn's syndrome
C1384514|T047|PT|255.12|ICD9CM|Conn's syndrome|Conn's syndrome
C0004775|T047|AB|255.13|ICD9CM|Bartter's syndrome|Bartter's syndrome
C0004775|T047|PT|255.13|ICD9CM|Bartter's syndrome|Bartter's syndrome
C1260387|T047|PT|255.14|ICD9CM|Other secondary aldosteronism|Other secondary aldosteronism
C1260387|T047|AB|255.14|ICD9CM|Secondry aldosternsm NEC|Secondry aldosternsm NEC
C0701163|T047|AB|255.2|ICD9CM|Adrenogenital disorders|Adrenogenital disorders
C0701163|T047|PT|255.2|ICD9CM|Adrenogenital disorders|Adrenogenital disorders
C0348461|T047|AB|255.3|ICD9CM|Corticoadren overact NEC|Corticoadren overact NEC
C0348461|T047|PT|255.3|ICD9CM|Other corticoadrenal overactivity|Other corticoadrenal overactivity
C0405580|T047|HT|255.4|ICD9CM|Corticoadrenal insufficiency|Corticoadrenal insufficiency
C1955741|T047|PT|255.41|ICD9CM|Glucocorticoid deficiency|Glucocorticoid deficiency
C1955741|T047|AB|255.41|ICD9CM|Glucocorticoid deficient|Glucocorticoid deficient
C1955743|T047|AB|255.42|ICD9CM|Mineralcorticoid defcnt|Mineralcorticoid defcnt
C1955743|T047|PT|255.42|ICD9CM|Mineralocorticoid deficiency|Mineralocorticoid deficiency
C0154205|T047|AB|255.5|ICD9CM|Adrenal hypofunction NEC|Adrenal hypofunction NEC
C0154205|T047|PT|255.5|ICD9CM|Other adrenal hypofunction|Other adrenal hypofunction
C0154206|T047|AB|255.6|ICD9CM|Medulloadrenal hyperfunc|Medulloadrenal hyperfunc
C0154206|T047|PT|255.6|ICD9CM|Medulloadrenal hyperfunction|Medulloadrenal hyperfunction
C0154207|T047|AB|255.8|ICD9CM|Adrenal disorder NEC|Adrenal disorder NEC
C0154207|T047|PT|255.8|ICD9CM|Other specified disorders of adrenal glands|Other specified disorders of adrenal glands
C0001621|T047|AB|255.9|ICD9CM|Adrenal disorder NOS|Adrenal disorder NOS
C0001621|T047|PT|255.9|ICD9CM|Unspecified disorder of adrenal glands|Unspecified disorder of adrenal glands
C0154208|T047|HT|256|ICD9CM|Ovarian dysfunction|Ovarian dysfunction
C0154209|T047|AB|256.0|ICD9CM|Hyperestrogenism|Hyperestrogenism
C0154209|T047|PT|256.0|ICD9CM|Hyperestrogenism|Hyperestrogenism
C0154210|T047|PT|256.1|ICD9CM|Other ovarian hyperfunction|Other ovarian hyperfunction
C0154210|T047|AB|256.1|ICD9CM|Ovarian hyperfunc NEC|Ovarian hyperfunc NEC
C0154211|T033|AB|256.2|ICD9CM|Postablativ ovarian fail|Postablativ ovarian fail
C0154211|T033|PT|256.2|ICD9CM|Postablative ovarian failure|Postablative ovarian failure
C0029697|T047|HT|256.3|ICD9CM|Other ovarian failure|Other ovarian failure
C0025322|T047|AB|256.31|ICD9CM|Premature menopause|Premature menopause
C0025322|T047|PT|256.31|ICD9CM|Premature menopause|Premature menopause
C0029697|T047|PT|256.39|ICD9CM|Other ovarian failure|Other ovarian failure
C0029697|T047|AB|256.39|ICD9CM|Ovarian failure NEC|Ovarian failure NEC
C0032460|T047|AB|256.4|ICD9CM|Polycystic ovaries|Polycystic ovaries
C0032460|T047|PT|256.4|ICD9CM|Polycystic ovaries|Polycystic ovaries
C0154212|T047|PT|256.8|ICD9CM|Other ovarian dysfunction|Other ovarian dysfunction
C0154212|T047|AB|256.8|ICD9CM|Ovarian dysfunction NEC|Ovarian dysfunction NEC
C0154208|T047|AB|256.9|ICD9CM|Ovarian dysfunction NOS|Ovarian dysfunction NOS
C0154208|T047|PT|256.9|ICD9CM|Unspecified ovarian dysfunction|Unspecified ovarian dysfunction
C0405581|T047|HT|257|ICD9CM|Testicular dysfunction|Testicular dysfunction
C0154215|T047|AB|257.0|ICD9CM|Testicular hyperfunction|Testicular hyperfunction
C0154215|T047|PT|257.0|ICD9CM|Testicular hyperfunction|Testicular hyperfunction
C0154216|T047|AB|257.1|ICD9CM|Postablat testic hypofun|Postablat testic hypofun
C0154216|T047|PT|257.1|ICD9CM|Postablative testicular hypofunction|Postablative testicular hypofunction
C0029858|T047|PT|257.2|ICD9CM|Other testicular hypofunction|Other testicular hypofunction
C0029858|T047|AB|257.2|ICD9CM|Testicular hypofunc NEC|Testicular hypofunc NEC
C0029857|T046|PT|257.8|ICD9CM|Other testicular dysfunction|Other testicular dysfunction
C0029857|T046|AB|257.8|ICD9CM|Testicular dysfunct NEC|Testicular dysfunct NEC
C0405581|T047|AB|257.9|ICD9CM|Testicular dysfunct NOS|Testicular dysfunct NOS
C0405581|T047|PT|257.9|ICD9CM|Unspecified testicular dysfunction|Unspecified testicular dysfunction
C0154218|T047|HT|258|ICD9CM|Polyglandular dysfunction and related disorders|Polyglandular dysfunction and related disorders
C0311355|T191|HT|258.0|ICD9CM|Polyglandular activity in multiple endocrine adenomatosis|Polyglandular activity in multiple endocrine adenomatosis
C0025267|T191|AB|258.01|ICD9CM|Mult endo neoplas type I|Mult endo neoplas type I
C0025267|T191|PT|258.01|ICD9CM|Multiple endocrine neoplasia [MEN] type I|Multiple endocrine neoplasia [MEN] type I
C0025268|T191|AB|258.02|ICD9CM|Mult endo neop type IIA|Mult endo neop type IIA
C0025268|T191|PT|258.02|ICD9CM|Multiple endocrine neoplasia [MEN] type IIA|Multiple endocrine neoplasia [MEN] type IIA
C0025269|T191|AB|258.03|ICD9CM|Mult endo neop type IIB|Mult endo neop type IIB
C0025269|T191|PT|258.03|ICD9CM|Multiple endocrine neoplasia [MEN] type IIB|Multiple endocrine neoplasia [MEN] type IIB
C0154220|T047|AB|258.1|ICD9CM|Comb endocr dysfunct NEC|Comb endocr dysfunct NEC
C0154220|T047|PT|258.1|ICD9CM|Other combinations of endocrine dysfunction|Other combinations of endocrine dysfunction
C0154221|T047|PT|258.8|ICD9CM|Other specified polyglandular dysfunction|Other specified polyglandular dysfunction
C0154221|T047|AB|258.8|ICD9CM|Polyglandul dysfunc NEC|Polyglandul dysfunc NEC
C0154222|T047|AB|258.9|ICD9CM|Polyglandul dysfunc NOS|Polyglandul dysfunc NOS
C0154222|T047|PT|258.9|ICD9CM|Polyglandular dysfunction, unspecified|Polyglandular dysfunction, unspecified
C0154223|T047|HT|259|ICD9CM|Other endocrine disorders|Other endocrine disorders
C0869499|T047|PT|259.0|ICD9CM|Delay in sexual development and puberty, not elsewhere classified|Delay in sexual development and puberty, not elsewhere classified
C0869499|T047|AB|259.0|ICD9CM|Delay sexual develop NEC|Delay sexual develop NEC
C0869515|T047|PT|259.1|ICD9CM|Precocious sexual development and puberty, not elsewhere classified|Precocious sexual development and puberty, not elsewhere classified
C0869515|T047|AB|259.1|ICD9CM|Sexual precocity NEC|Sexual precocity NEC
C0024586|T047|AB|259.2|ICD9CM|Carcinoid syndrome|Carcinoid syndrome
C0024586|T047|PT|259.2|ICD9CM|Carcinoid syndrome|Carcinoid syndrome
C0869496|T047|AB|259.3|ICD9CM|Ectopic hormone secr NEC|Ectopic hormone secr NEC
C0869496|T047|PT|259.3|ICD9CM|Ectopic hormone secretion, not elsewhere classified|Ectopic hormone secretion, not elsewhere classified
C0677577|T019|AB|259.4|ICD9CM|Dwarfism NEC|Dwarfism NEC
C0677577|T019|PT|259.4|ICD9CM|Dwarfism, not elsewhere classified|Dwarfism, not elsewhere classified
C0039585|T047|HT|259.5|ICD9CM|Androgen insensitivity syndrome|Androgen insensitivity syndrome
C2349400|T047|PT|259.50|ICD9CM|Androgen insensitivity, unspecified|Androgen insensitivity, unspecified
C2349400|T047|AB|259.50|ICD9CM|Androgen insensitvty NOS|Androgen insensitvty NOS
C0039585|T047|PT|259.51|ICD9CM|Androgen insensitivity syndrome|Androgen insensitivity syndrome
C0039585|T047|AB|259.51|ICD9CM|Androgen insensitvty syn|Androgen insensitvty syn
C0268301|T047|AB|259.52|ICD9CM|Part androgen insnsitvty|Part androgen insnsitvty
C0268301|T047|PT|259.52|ICD9CM|Partial androgen insensitivity|Partial androgen insensitivity
C0029793|T047|AB|259.8|ICD9CM|Endocrine disorders NEC|Endocrine disorders NEC
C0029793|T047|PT|259.8|ICD9CM|Other specified endocrine disorders|Other specified endocrine disorders
C0014130|T047|AB|259.9|ICD9CM|Endocrine disorder NOS|Endocrine disorder NOS
C0014130|T047|PT|259.9|ICD9CM|Unspecified endocrine disorder|Unspecified endocrine disorder
C0022806|T047|AB|260|ICD9CM|Kwashiorkor|Kwashiorkor
C0022806|T047|PT|260|ICD9CM|Kwashiorkor|Kwashiorkor
C4761312|T047|HT|260-269.99|ICD9CM|NUTRITIONAL DEFICIENCIES|NUTRITIONAL DEFICIENCIES
C0086588|T047|AB|261|ICD9CM|Nutritional marasmus|Nutritional marasmus
C0086588|T047|PT|261|ICD9CM|Nutritional marasmus|Nutritional marasmus
C0267981|T047|AB|262|ICD9CM|Oth severe malnutrition|Oth severe malnutrition
C0267981|T047|PT|262|ICD9CM|Other severe protein-calorie malnutrition|Other severe protein-calorie malnutrition
C0687762|T047|HT|263|ICD9CM|Other and unspecified protein-calorie malnutrition|Other and unspecified protein-calorie malnutrition
C0154227|T047|AB|263.0|ICD9CM|Malnutrition mod degree|Malnutrition mod degree
C0154227|T047|PT|263.0|ICD9CM|Malnutrition of moderate degree|Malnutrition of moderate degree
C0154228|T047|AB|263.1|ICD9CM|Malnutrition mild degree|Malnutrition mild degree
C0154228|T047|PT|263.1|ICD9CM|Malnutrition of mild degree|Malnutrition of mild degree
C0154229|T047|AB|263.2|ICD9CM|Arrest devel d/t malnutr|Arrest devel d/t malnutr
C0154229|T047|PT|263.2|ICD9CM|Arrested development following protein-calorie malnutrition|Arrested development following protein-calorie malnutrition
C0154230|T047|PT|263.8|ICD9CM|Other protein-calorie malnutrition|Other protein-calorie malnutrition
C0154230|T047|AB|263.8|ICD9CM|Protein-cal malnutr NEC|Protein-cal malnutr NEC
C0033677|T046|AB|263.9|ICD9CM|Protein-cal malnutr NOS|Protein-cal malnutr NOS
C0033677|T046|PT|263.9|ICD9CM|Unspecified protein-calorie malnutrition|Unspecified protein-calorie malnutrition
C0042842|T047|HT|264|ICD9CM|Vitamin A deficiency|Vitamin A deficiency
C0154231|T047|AB|264.0|ICD9CM|Vit A conjunctiv xerosis|Vit A conjunctiv xerosis
C0154231|T047|PT|264.0|ICD9CM|Vitamin A deficiency with conjunctival xerosis|Vitamin A deficiency with conjunctival xerosis
C0154232|T047|AB|264.1|ICD9CM|Vit A bitot's spot|Vit A bitot's spot
C0154232|T047|PT|264.1|ICD9CM|Vitamin A deficiency with conjunctival xerosis and Bitot's spot|Vitamin A deficiency with conjunctival xerosis and Bitot's spot
C0154233|T047|AB|264.2|ICD9CM|Vit A corneal xerosis|Vit A corneal xerosis
C0154233|T047|PT|264.2|ICD9CM|Vitamin A deficiency with corneal xerosis|Vitamin A deficiency with corneal xerosis
C0154234|T047|AB|264.3|ICD9CM|Vit A cornea ulcer/xeros|Vit A cornea ulcer/xeros
C0154234|T047|PT|264.3|ICD9CM|Vitamin A deficiency with corneal ulceration and xerosis|Vitamin A deficiency with corneal ulceration and xerosis
C0154235|T047|AB|264.4|ICD9CM|Vit A keratomalacia|Vit A keratomalacia
C0154235|T047|PT|264.4|ICD9CM|Vitamin A deficiency with keratomalacia|Vitamin A deficiency with keratomalacia
C0154236|T047|AB|264.5|ICD9CM|Vit A night blindness|Vit A night blindness
C0154236|T047|PT|264.5|ICD9CM|Vitamin A deficiency with night blindness|Vitamin A deficiency with night blindness
C0154237|T047|AB|264.6|ICD9CM|Vit A def w corneal scar|Vit A def w corneal scar
C0154237|T047|PT|264.6|ICD9CM|Vitamin A deficiency with xerophthalmic scars of cornea|Vitamin A deficiency with xerophthalmic scars of cornea
C0154238|T047|PT|264.7|ICD9CM|Other ocular manifestations of vitamin A deficiency|Other ocular manifestations of vitamin A deficiency
C0154238|T047|AB|264.7|ICD9CM|Vit A ocular defic NEC|Vit A ocular defic NEC
C0029665|T047|PT|264.8|ICD9CM|Other manifestations of vitamin A deficiency|Other manifestations of vitamin A deficiency
C0029665|T047|AB|264.8|ICD9CM|Vitamin A deficiency NEC|Vitamin A deficiency NEC
C0042842|T047|PT|264.9|ICD9CM|Unspecified vitamin A deficiency|Unspecified vitamin A deficiency
C0042842|T047|AB|264.9|ICD9CM|Vitamin A deficiency NOS|Vitamin A deficiency NOS
C0154239|T047|HT|265|ICD9CM|Thiamine and niacin deficiency states|Thiamine and niacin deficiency states
C0005122|T047|AB|265.0|ICD9CM|Beriberi|Beriberi
C0005122|T047|PT|265.0|ICD9CM|Beriberi|Beriberi
C0029510|T047|PT|265.1|ICD9CM|Other and unspecified manifestations of thiamine deficiency|Other and unspecified manifestations of thiamine deficiency
C0029510|T047|AB|265.1|ICD9CM|Thiamine defic NEC/NOS|Thiamine defic NEC/NOS
C0030783|T047|AB|265.2|ICD9CM|Pellagra|Pellagra
C0030783|T047|PT|265.2|ICD9CM|Pellagra|Pellagra
C0042850|T047|HT|266|ICD9CM|Deficiency of B-complex components|Deficiency of B-complex components
C0035528|T047|AB|266.0|ICD9CM|Ariboflavinosis|Ariboflavinosis
C0035528|T047|PT|266.0|ICD9CM|Ariboflavinosis|Ariboflavinosis
C0936215|T047|PT|266.1|ICD9CM|Vitamin B6 deficiency|Vitamin B6 deficiency
C0936215|T047|AB|266.1|ICD9CM|Vitamin b6 deficiency|Vitamin b6 deficiency
C0029523|T047|AB|266.2|ICD9CM|B-complex defic NEC|B-complex defic NEC
C0029523|T047|PT|266.2|ICD9CM|Other B-complex deficiencies|Other B-complex deficiencies
C0042850|T047|PT|266.9|ICD9CM|Unspecified vitamin B deficiency|Unspecified vitamin B deficiency
C0042850|T047|AB|266.9|ICD9CM|Vitamin b deficiency NOS|Vitamin b deficiency NOS
C0003969|T047|AB|267|ICD9CM|Ascorbic acid deficiency|Ascorbic acid deficiency
C0003969|T047|PT|267|ICD9CM|Ascorbic acid deficiency|Ascorbic acid deficiency
C0042870|T047|HT|268|ICD9CM|Vitamin D deficiency|Vitamin D deficiency
C0221468|T047|AB|268.0|ICD9CM|Rickets, active|Rickets, active
C0221468|T047|PT|268.0|ICD9CM|Rickets, active|Rickets, active
C0154240|T046|AB|268.1|ICD9CM|Rickets, late effect|Rickets, late effect
C0154240|T046|PT|268.1|ICD9CM|Rickets, late effect|Rickets, late effect
C0029442|T047|AB|268.2|ICD9CM|Osteomalacia NOS|Osteomalacia NOS
C0029442|T047|PT|268.2|ICD9CM|Osteomalacia, unspecified|Osteomalacia, unspecified
C0042870|T047|PT|268.9|ICD9CM|Unspecified vitamin D deficiency|Unspecified vitamin D deficiency
C0042870|T047|AB|268.9|ICD9CM|Vitamin D deficiency NOS|Vitamin D deficiency NOS
C0154241|T047|HT|269|ICD9CM|Other nutritional deficiencies|Other nutritional deficiencies
C0042880|T047|PT|269.0|ICD9CM|Deficiency of vitamin K|Deficiency of vitamin K
C0042880|T047|AB|269.0|ICD9CM|Deficiency of vitamin k|Deficiency of vitamin k
C0011157|T047|PT|269.1|ICD9CM|Deficiency of other vitamins|Deficiency of other vitamins
C0011157|T047|AB|269.1|ICD9CM|Vitamin Deficiency NEC|Vitamin Deficiency NEC
C1510471|T047|PT|269.2|ICD9CM|Unspecified vitamin deficiency|Unspecified vitamin deficiency
C1510471|T047|AB|269.2|ICD9CM|Vitamin Deficiency NOS|Vitamin Deficiency NOS
C0869423|T047|AB|269.3|ICD9CM|Mineral deficiency NEC|Mineral deficiency NEC
C0869423|T047|PT|269.3|ICD9CM|Mineral deficiency, not elsewhere classified|Mineral deficiency, not elsewhere classified
C0154241|T047|AB|269.8|ICD9CM|Nutrition deficiency NEC|Nutrition deficiency NEC
C0154241|T047|PT|269.8|ICD9CM|Other nutritional deficiency|Other nutritional deficiency
C4761312|T047|AB|269.9|ICD9CM|Nutrition deficiency NOS|Nutrition deficiency NOS
C4761312|T047|PT|269.9|ICD9CM|Unspecified nutritional deficiency|Unspecified nutritional deficiency
C0002514|T047|HT|270|ICD9CM|Disorders of amino-acid transport and metabolism|Disorders of amino-acid transport and metabolism
C0178259|T046|HT|270-279.99|ICD9CM|OTHER METABOLIC AND IMMUNITY DISORDERS|OTHER METABOLIC AND IMMUNITY DISORDERS
C0268641|T047|AB|270.0|ICD9CM|Amino-acid transport dis|Amino-acid transport dis
C0268641|T047|PT|270.0|ICD9CM|Disturbances of amino-acid transport|Disturbances of amino-acid transport
C0031485|T047|AB|270.1|ICD9CM|Phenylketonuria - pku|Phenylketonuria - pku
C0031485|T047|PT|270.1|ICD9CM|Phenylketonuria [PKU]|Phenylketonuria [PKU]
C0348483|T047|AB|270.2|ICD9CM|Arom amin-acid metab NEC|Arom amin-acid metab NEC
C0348483|T047|PT|270.2|ICD9CM|Other disturbances of aromatic amino-acid metabolism|Other disturbances of aromatic amino-acid metabolism
C0342712|T047|AB|270.3|ICD9CM|Bran-chain amin-acid dis|Bran-chain amin-acid dis
C0342712|T047|PT|270.3|ICD9CM|Disturbances of branched-chain amino-acid metabolism|Disturbances of branched-chain amino-acid metabolism
C0268613|T047|PT|270.4|ICD9CM|Disturbances of sulphur-bearing amino-acid metabolism|Disturbances of sulphur-bearing amino-acid metabolism
C0268613|T047|AB|270.4|ICD9CM|Sulph amino-acid met dis|Sulph amino-acid met dis
C0268512|T047|AB|270.5|ICD9CM|Dis histidine metabolism|Dis histidine metabolism
C0268512|T047|PT|270.5|ICD9CM|Disturbances of histidine metabolism|Disturbances of histidine metabolism
C0154246|T047|AB|270.6|ICD9CM|Dis urea cycle metabol|Dis urea cycle metabol
C0154246|T047|PT|270.6|ICD9CM|Disorders of urea cycle metabolism|Disorders of urea cycle metabolism
C0154247|T047|PT|270.7|ICD9CM|Other disturbances of straight-chain amino-acid metabolism|Other disturbances of straight-chain amino-acid metabolism
C0154247|T047|AB|270.7|ICD9CM|Straig amin-acid met NEC|Straig amin-acid met NEC
C0029774|T047|AB|270.8|ICD9CM|Dis amino-acid metab NEC|Dis amino-acid metab NEC
C0029774|T047|PT|270.8|ICD9CM|Other specified disorders of amino-acid metabolism|Other specified disorders of amino-acid metabolism
C0002514|T047|AB|270.9|ICD9CM|Dis amino-acid metab NOS|Dis amino-acid metab NOS
C0002514|T047|PT|270.9|ICD9CM|Unspecified disorder of amino-acid metabolism|Unspecified disorder of amino-acid metabolism
C0154249|T047|HT|271|ICD9CM|Disorders of carbohydrate transport and metabolism|Disorders of carbohydrate transport and metabolism
C0017919|T047|AB|271.0|ICD9CM|Glycogenosis|Glycogenosis
C0017919|T047|PT|271.0|ICD9CM|Glycogenosis|Glycogenosis
C0016952|T047|AB|271.1|ICD9CM|Galactosemia|Galactosemia
C0016952|T047|PT|271.1|ICD9CM|Galactosemia|Galactosemia
C0016751|T047|AB|271.2|ICD9CM|Hered fructose intoleran|Hered fructose intoleran
C0016751|T047|PT|271.2|ICD9CM|Hereditary fructose intolerance|Hereditary fructose intolerance
C0021830|T047|AB|271.3|ICD9CM|Disaccharidase def/malab|Disaccharidase def/malab
C0021830|T047|PT|271.3|ICD9CM|Intestinal disaccharidase deficiencies and disaccharide malabsorption|Intestinal disaccharidase deficiencies and disaccharide malabsorption
C0017980|T047|AB|271.4|ICD9CM|Renal glycosuria|Renal glycosuria
C0017980|T047|PT|271.4|ICD9CM|Renal glycosuria|Renal glycosuria
C0029777|T047|AB|271.8|ICD9CM|Dis carbohydr metab NEC|Dis carbohydr metab NEC
C0029777|T047|PT|271.8|ICD9CM|Other specified disorders of carbohydrate transport and metabolism|Other specified disorders of carbohydrate transport and metabolism
C0154249|T047|AB|271.9|ICD9CM|Dis carbohydr metab NOS|Dis carbohydr metab NOS
C0154249|T047|PT|271.9|ICD9CM|Unspecified disorder of carbohydrate transport and metabolism|Unspecified disorder of carbohydrate transport and metabolism
C0154251|T047|HT|272|ICD9CM|Disorders of lipoid metabolism|Disorders of lipoid metabolism
C0678189|T047|AB|272.0|ICD9CM|Pure hypercholesterolem|Pure hypercholesterolem
C0678189|T047|PT|272.0|ICD9CM|Pure hypercholesterolemia|Pure hypercholesterolemia
C0020480|T047|AB|272.1|ICD9CM|Pure hyperglyceridemia|Pure hyperglyceridemia
C0020480|T047|PT|272.1|ICD9CM|Pure hyperglyceridemia|Pure hyperglyceridemia
C2047520|T047|AB|272.2|ICD9CM|Mixed hyperlipidemia|Mixed hyperlipidemia
C2047520|T047|PT|272.2|ICD9CM|Mixed hyperlipidemia|Mixed hyperlipidemia
C0023817|T047|AB|272.3|ICD9CM|Hyperchylomicronemia|Hyperchylomicronemia
C0023817|T047|PT|272.3|ICD9CM|Hyperchylomicronemia|Hyperchylomicronemia
C0348494|T047|AB|272.4|ICD9CM|Hyperlipidemia NEC/NOS|Hyperlipidemia NEC/NOS
C0348494|T047|PT|272.4|ICD9CM|Other and unspecified hyperlipidemia|Other and unspecified hyperlipidemia
C0020623|T033|AB|272.5|ICD9CM|Lipoprotein deficiencies|Lipoprotein deficiencies
C0020623|T033|PT|272.5|ICD9CM|Lipoprotein deficiencies|Lipoprotein deficiencies
C0023787|T047|AB|272.6|ICD9CM|Lipodystrophy|Lipodystrophy
C0023787|T047|PT|272.6|ICD9CM|Lipodystrophy|Lipodystrophy
C0023794|T047|AB|272.7|ICD9CM|Lipidoses|Lipidoses
C0023794|T047|PT|272.7|ICD9CM|Lipidoses|Lipidoses
C0029591|T047|AB|272.8|ICD9CM|Lipoid metabol dis NEC|Lipoid metabol dis NEC
C0029591|T047|PT|272.8|ICD9CM|Other disorders of lipoid metabolism|Other disorders of lipoid metabolism
C0154251|T047|AB|272.9|ICD9CM|Lipoid metabol dis NOS|Lipoid metabol dis NOS
C0154251|T047|PT|272.9|ICD9CM|Unspecified disorder of lipoid metabolism|Unspecified disorder of lipoid metabolism
C3875058|T047|HT|273|ICD9CM|Disorders of plasma protein metabolism|Disorders of plasma protein metabolism
C0154254|T047|AB|273.0|ICD9CM|Polyclon hypergammaglobu|Polyclon hypergammaglobu
C0154254|T047|PT|273.0|ICD9CM|Polyclonal hypergammaglobulinemia|Polyclonal hypergammaglobulinemia
C0026471|T191|AB|273.1|ICD9CM|Monoclon paraproteinemia|Monoclon paraproteinemia
C0026471|T191|PT|273.1|ICD9CM|Monoclonal paraproteinemia|Monoclonal paraproteinemia
C0029698|T191|PT|273.2|ICD9CM|Other paraproteinemias|Other paraproteinemias
C0029698|T191|AB|273.2|ICD9CM|Paraproteinemia NEC|Paraproteinemia NEC
C0024419|T191|AB|273.3|ICD9CM|Macroglobulinemia|Macroglobulinemia
C0024419|T191|PT|273.3|ICD9CM|Macroglobulinemia|Macroglobulinemia
C0221757|T047|AB|273.4|ICD9CM|Alpha-1-antitrypsin def|Alpha-1-antitrypsin def
C0221757|T047|PT|273.4|ICD9CM|Alpha-1-antitrypsin deficiency|Alpha-1-antitrypsin deficiency
C0029594|T047|AB|273.8|ICD9CM|Dis plas protein met NEC|Dis plas protein met NEC
C0029594|T047|PT|273.8|ICD9CM|Other disorders of plasma protein metabolism|Other disorders of plasma protein metabolism
C3875058|T047|AB|273.9|ICD9CM|Dis plas protein met NOS|Dis plas protein met NOS
C3875058|T047|PT|273.9|ICD9CM|Unspecified disorder of plasma protein metabolism|Unspecified disorder of plasma protein metabolism
C0018099|T047|HT|274|ICD9CM|Gout|Gout
C0003868|T047|HT|274.0|ICD9CM|Gouty arthropathy|Gouty arthropathy
C0003868|T047|AB|274.00|ICD9CM|Gouty arthropathy NOS|Gouty arthropathy NOS
C0003868|T047|PT|274.00|ICD9CM|Gouty arthropathy, unspecified|Gouty arthropathy, unspecified
C0149896|T047|AB|274.01|ICD9CM|Acute gouty arthropathy|Acute gouty arthropathy
C0149896|T047|PT|274.01|ICD9CM|Acute gouty arthropathy|Acute gouty arthropathy
C2712886|T047|AB|274.02|ICD9CM|Chr gouty atrph wo tophi|Chr gouty atrph wo tophi
C2712886|T047|PT|274.02|ICD9CM|Chronic gouty arthropathy without mention of tophus (tophi)|Chronic gouty arthropathy without mention of tophus (tophi)
C2712899|T047|AB|274.03|ICD9CM|Chr gouty atroph w tophi|Chr gouty atroph w tophi
C2712899|T047|PT|274.03|ICD9CM|Chronic gouty arthropathy with tophus (tophi)|Chronic gouty arthropathy with tophus (tophi)
C0391820|T047|HT|274.1|ICD9CM|Gouty nephropathy|Gouty nephropathy
C0391820|T047|AB|274.10|ICD9CM|Gouty nephropathy NOS|Gouty nephropathy NOS
C0391820|T047|PT|274.10|ICD9CM|Gouty nephropathy, unspecified|Gouty nephropathy, unspecified
C0403719|T047|AB|274.11|ICD9CM|Uric acid nephrolithias|Uric acid nephrolithias
C0403719|T047|PT|274.11|ICD9CM|Uric acid nephrolithiasis|Uric acid nephrolithiasis
C0154256|T047|AB|274.19|ICD9CM|Gouty nephropathy NEC|Gouty nephropathy NEC
C0154256|T047|PT|274.19|ICD9CM|Other gouty nephropathy|Other gouty nephropathy
C0154257|T047|HT|274.8|ICD9CM|Gout with other specified manifestations|Gout with other specified manifestations
C0154258|T033|AB|274.81|ICD9CM|Gouty tophi of ear|Gouty tophi of ear
C0154258|T033|PT|274.81|ICD9CM|Gouty tophi of ear|Gouty tophi of ear
C0154259|T047|PT|274.82|ICD9CM|Gouty tophi of other sites, except ear|Gouty tophi of other sites, except ear
C0154259|T047|AB|274.82|ICD9CM|Gouty tophi site NEC|Gouty tophi site NEC
C0154257|T047|AB|274.89|ICD9CM|Gout w manifestation NEC|Gout w manifestation NEC
C0154257|T047|PT|274.89|ICD9CM|Gout with other specified manifestations|Gout with other specified manifestations
C0018099|T047|AB|274.9|ICD9CM|Gout NOS|Gout NOS
C0018099|T047|PT|274.9|ICD9CM|Gout, unspecified|Gout, unspecified
C0154260|T046|HT|275|ICD9CM|Disorders of mineral metabolism|Disorders of mineral metabolism
C0012715|T047|HT|275.0|ICD9CM|Disorders of iron metabolism|Disorders of iron metabolism
C0392514|T047|AB|275.01|ICD9CM|Heredit hemochromatosis|Heredit hemochromatosis
C0392514|T047|PT|275.01|ICD9CM|Hereditary hemochromatosis|Hereditary hemochromatosis
C2921014|T047|AB|275.02|ICD9CM|Hemochromatos-rbc trans|Hemochromatos-rbc trans
C2921014|T047|PT|275.02|ICD9CM|Hemochromatosis due to repeated red blood cell transfusions|Hemochromatosis due to repeated red blood cell transfusions
C2921018|T047|AB|275.03|ICD9CM|Hemochromatosis NEC|Hemochromatosis NEC
C2921018|T047|PT|275.03|ICD9CM|Other hemochromatosis|Other hemochromatosis
C2874299|T047|AB|275.09|ICD9CM|Disord iron metablsm NEC|Disord iron metablsm NEC
C2874299|T047|PT|275.09|ICD9CM|Other disorders of iron metabolism|Other disorders of iron metabolism
C0012714|T047|AB|275.1|ICD9CM|Dis copper metabolism|Dis copper metabolism
C0012714|T047|PT|275.1|ICD9CM|Disorders of copper metabolism|Disorders of copper metabolism
C0012716|T047|AB|275.2|ICD9CM|Dis magnesium metabolism|Dis magnesium metabolism
C0012716|T047|PT|275.2|ICD9CM|Disorders of magnesium metabolism|Disorders of magnesium metabolism
C0031707|T047|AB|275.3|ICD9CM|Dis phosphorus metabol|Dis phosphorus metabol
C0031707|T047|PT|275.3|ICD9CM|Disorders of phosphorus metabolism|Disorders of phosphorus metabolism
C0006705|T047|HT|275.4|ICD9CM|Disorders of calcium metabolism|Disorders of calcium metabolism
C0006705|T047|AB|275.40|ICD9CM|Dis calcium metablsm NOS|Dis calcium metablsm NOS
C0006705|T047|PT|275.40|ICD9CM|Unspecified disorder of calcium metabolism|Unspecified disorder of calcium metabolism
C0020598|T047|AB|275.41|ICD9CM|Hypocalcemia|Hypocalcemia
C0020598|T047|PT|275.41|ICD9CM|Hypocalcemia|Hypocalcemia
C0020437|T047|AB|275.42|ICD9CM|Hypercalcemia|Hypercalcemia
C0020437|T047|PT|275.42|ICD9CM|Hypercalcemia|Hypercalcemia
C0489982|T047|AB|275.49|ICD9CM|Dis calcium metablsm NEC|Dis calcium metablsm NEC
C0489982|T047|PT|275.49|ICD9CM|Other disorders of calcium metabolism|Other disorders of calcium metabolism
C0342635|T047|PT|275.5|ICD9CM|Hungry bone syndrome|Hungry bone syndrome
C0342635|T047|AB|275.5|ICD9CM|Hungry bone syndrome|Hungry bone syndrome
C0154261|T046|AB|275.8|ICD9CM|Dis mineral metabol NEC|Dis mineral metabol NEC
C0154261|T046|PT|275.8|ICD9CM|Other specified disorders of mineral metabolism|Other specified disorders of mineral metabolism
C0154260|T046|AB|275.9|ICD9CM|Dis mineral metabol NOS|Dis mineral metabol NOS
C0154260|T046|PT|275.9|ICD9CM|Unspecified disorder of mineral metabolism|Unspecified disorder of mineral metabolism
C0267994|T046|HT|276|ICD9CM|Disorders of fluid, electrolyte, and acid-base balance|Disorders of fluid, electrolyte, and acid-base balance
C0342580|T047|AB|276.0|ICD9CM|Hyperosmolality|Hyperosmolality
C0342580|T047|PT|276.0|ICD9CM|Hyperosmolality and/or hypernatremia|Hyperosmolality and/or hypernatremia
C0020645|T033|AB|276.1|ICD9CM|Hyposmolality|Hyposmolality
C0020645|T033|PT|276.1|ICD9CM|Hyposmolality and/or hyponatremia|Hyposmolality and/or hyponatremia
C0001122|T046|AB|276.2|ICD9CM|Acidosis|Acidosis
C0001122|T046|PT|276.2|ICD9CM|Acidosis|Acidosis
C0002063|T047|AB|276.3|ICD9CM|Alkalosis|Alkalosis
C0002063|T047|PT|276.3|ICD9CM|Alkalosis|Alkalosis
C0154264|T047|AB|276.4|ICD9CM|Mixed acid-base bal dis|Mixed acid-base bal dis
C0154264|T047|PT|276.4|ICD9CM|Mixed acid-base balance disorder|Mixed acid-base balance disorder
C0546884|T033|HT|276.5|ICD9CM|Volume depletion|Volume depletion
C0546884|T033|AB|276.50|ICD9CM|Volume depletion NOS|Volume depletion NOS
C0546884|T033|PT|276.50|ICD9CM|Volume depletion, unspecified|Volume depletion, unspecified
C0011175|T047|AB|276.51|ICD9CM|Dehydration|Dehydration
C0011175|T047|PT|276.51|ICD9CM|Dehydration|Dehydration
C0546884|T033|AB|276.52|ICD9CM|Hypovolemia|Hypovolemia
C0546884|T033|PT|276.52|ICD9CM|Hypovolemia|Hypovolemia
C0546817|T046|HT|276.6|ICD9CM|Fluid overload|Fluid overload
C2921022|T046|AB|276.61|ICD9CM|Transfsn w circ overload|Transfsn w circ overload
C2921022|T046|PT|276.61|ICD9CM|Transfusion associated circulatory overload|Transfusion associated circulatory overload
C2921023|T047|AB|276.69|ICD9CM|Fluid overload NEC|Fluid overload NEC
C2921023|T047|PT|276.69|ICD9CM|Other fluid overload|Other fluid overload
C0020461|T033|AB|276.7|ICD9CM|Hyperpotassemia|Hyperpotassemia
C0020461|T033|PT|276.7|ICD9CM|Hyperpotassemia|Hyperpotassemia
C0020621|T033|AB|276.8|ICD9CM|Hypopotassemia|Hypopotassemia
C0020621|T033|PT|276.8|ICD9CM|Hypopotassemia|Hypopotassemia
C0868890|T046|AB|276.9|ICD9CM|Electrolyt/fluid dis NEC|Electrolyt/fluid dis NEC
C0868890|T046|PT|276.9|ICD9CM|Electrolyte and fluid disorders not elsewhere classified|Electrolyte and fluid disorders not elsewhere classified
C0268329|T047|HT|277|ICD9CM|Other and unspecified disorders of metabolism|Other and unspecified disorders of metabolism
C0010674|T047|HT|277.0|ICD9CM|Cystic fibrosis|Cystic fibrosis
C0010676|T047|AB|277.00|ICD9CM|Cystic fibros w/o ileus|Cystic fibros w/o ileus
C0010676|T047|PT|277.00|ICD9CM|Cystic fibrosis without mention of meconium ileus|Cystic fibrosis without mention of meconium ileus
C0546982|T047|AB|277.01|ICD9CM|Cystic fibrosis w ileus|Cystic fibrosis w ileus
C0546982|T047|PT|277.01|ICD9CM|Cystic fibrosis with meconium ileus|Cystic fibrosis with meconium ileus
C0348815|T047|AB|277.02|ICD9CM|Cystic fibros w pul man|Cystic fibros w pul man
C0348815|T047|PT|277.02|ICD9CM|Cystic fibrosis with pulmonary manifestations|Cystic fibrosis with pulmonary manifestations
C1135187|T047|AB|277.03|ICD9CM|Cystic fibrosis w GI man|Cystic fibrosis w GI man
C1135187|T047|PT|277.03|ICD9CM|Cystic fibrosis with gastrointestinal manifestations|Cystic fibrosis with gastrointestinal manifestations
C0494350|T047|AB|277.09|ICD9CM|Cystic fibrosis NEC|Cystic fibrosis NEC
C0494350|T047|PT|277.09|ICD9CM|Cystic fibrosis with other manifestations|Cystic fibrosis with other manifestations
C0032708|T047|AB|277.1|ICD9CM|Dis porphyrin metabolism|Dis porphyrin metabolism
C0032708|T047|PT|277.1|ICD9CM|Disorders of porphyrin metabolism|Disorders of porphyrin metabolism
C0029595|T047|PT|277.2|ICD9CM|Other disorders of purine and pyrimidine metabolism|Other disorders of purine and pyrimidine metabolism
C0029595|T047|AB|277.2|ICD9CM|Purine/pyrimid dis NEC|Purine/pyrimid dis NEC
C0002726|T047|HT|277.3|ICD9CM|Amyloidosis|Amyloidosis
C0002726|T047|AB|277.30|ICD9CM|Amyloidosis NOS|Amyloidosis NOS
C0002726|T047|PT|277.30|ICD9CM|Amyloidosis, unspecified|Amyloidosis, unspecified
C0031069|T047|AB|277.31|ICD9CM|Fam Mediterranean fever|Fam Mediterranean fever
C0031069|T047|PT|277.31|ICD9CM|Familial Mediterranean fever|Familial Mediterranean fever
C0348499|T047|AB|277.39|ICD9CM|Amyloidosis NEC|Amyloidosis NEC
C0348499|T047|PT|277.39|ICD9CM|Other amyloidosis|Other amyloidosis
C0012711|T047|AB|277.4|ICD9CM|Dis bilirubin excretion|Dis bilirubin excretion
C0012711|T047|PT|277.4|ICD9CM|Disorders of bilirubin excretion|Disorders of bilirubin excretion
C0026703|T047|AB|277.5|ICD9CM|Mucopolysaccharidosis|Mucopolysaccharidosis
C0026703|T047|PT|277.5|ICD9CM|Mucopolysaccharidosis|Mucopolysaccharidosis
C0029570|T047|AB|277.6|ICD9CM|Defic circul enzyme NEC|Defic circul enzyme NEC
C0029570|T047|PT|277.6|ICD9CM|Other deficiencies of circulating enzymes|Other deficiencies of circulating enzymes
C0524620|T047|PT|277.7|ICD9CM|Dysmetabolic syndrome X|Dysmetabolic syndrome X
C0524620|T047|AB|277.7|ICD9CM|Dysmetabolic syndrome x|Dysmetabolic syndrome x
C0494362|T047|HT|277.8|ICD9CM|Other specified disorders of metabolism|Other specified disorders of metabolism
C0342788|T047|PT|277.81|ICD9CM|Primary carnitine deficiency|Primary carnitine deficiency
C0342788|T047|AB|277.81|ICD9CM|Primary carnitine defncy|Primary carnitine defncy
C3875374|T047|PT|277.82|ICD9CM|Carnitine deficiency due to inborn errors of metabolism|Carnitine deficiency due to inborn errors of metabolism
C3875374|T047|AB|277.82|ICD9CM|Crnitne def d/t nb met|Crnitne def d/t nb met
C1260391|T046|AB|277.83|ICD9CM|Iatrogenic carnitine def|Iatrogenic carnitine def
C1260391|T046|PT|277.83|ICD9CM|Iatrogenic carnitine deficiency|Iatrogenic carnitine deficiency
C1260392|T047|PT|277.84|ICD9CM|Other secondary carnitine deficiency|Other secondary carnitine deficiency
C1260392|T047|AB|277.84|ICD9CM|Sec carnitine defncy NEC|Sec carnitine defncy NEC
C1456270|T047|AB|277.85|ICD9CM|Disorders acid oxidation|Disorders acid oxidation
C1456270|T047|PT|277.85|ICD9CM|Disorders of fatty acid oxidation|Disorders of fatty acid oxidation
C0282528|T047|AB|277.86|ICD9CM|Peroxisomal disorders|Peroxisomal disorders
C0282528|T047|PT|277.86|ICD9CM|Peroxisomal disorders|Peroxisomal disorders
C1456275|T047|AB|277.87|ICD9CM|Dis mitochondrial metab|Dis mitochondrial metab
C1456275|T047|PT|277.87|ICD9CM|Disorders of mitochondrial metabolism|Disorders of mitochondrial metabolism
C0041364|T047|PT|277.88|ICD9CM|Tumor lysis syndrome|Tumor lysis syndrome
C0041364|T047|AB|277.88|ICD9CM|Tumor lysis syndrome|Tumor lysis syndrome
C0494362|T047|AB|277.89|ICD9CM|Metabolism disorder NEC|Metabolism disorder NEC
C0494362|T047|PT|277.89|ICD9CM|Other specified disorders of metabolism|Other specified disorders of metabolism
C0025517|T047|AB|277.9|ICD9CM|Metabolism disorder NOS|Metabolism disorder NOS
C0025517|T047|PT|277.9|ICD9CM|Unspecified disorder of metabolism|Unspecified disorder of metabolism
C1561827|T047|HT|278|ICD9CM|Overweight, obesity and other hyperalimentation|Overweight, obesity and other hyperalimentation
C1561826|T047|HT|278.0|ICD9CM|Overweight and obesity|Overweight and obesity
C0028754|T047|AB|278.00|ICD9CM|Obesity NOS|Obesity NOS
C0028754|T047|PT|278.00|ICD9CM|Obesity, unspecified|Obesity, unspecified
C0028756|T047|AB|278.01|ICD9CM|Morbid obesity|Morbid obesity
C0028756|T047|PT|278.01|ICD9CM|Morbid obesity|Morbid obesity
C0497406|T033|AB|278.02|ICD9CM|Overweight|Overweight
C0497406|T033|PT|278.02|ICD9CM|Overweight|Overweight
C0031880|T047|AB|278.03|ICD9CM|Obesity hypovent synd|Obesity hypovent synd
C0031880|T047|PT|278.03|ICD9CM|Obesity hypoventilation syndrome|Obesity hypoventilation syndrome
C0154270|T033|AB|278.1|ICD9CM|Localized adiposity|Localized adiposity
C0154270|T033|PT|278.1|ICD9CM|Localized adiposity|Localized adiposity
C0020579|T047|PT|278.2|ICD9CM|Hypervitaminosis A|Hypervitaminosis A
C0020579|T047|AB|278.2|ICD9CM|Hypervitaminosis a|Hypervitaminosis a
C0154271|T047|AB|278.3|ICD9CM|Hypercarotinemia|Hypercarotinemia
C0154271|T047|PT|278.3|ICD9CM|Hypercarotinemia|Hypercarotinemia
C1442839|T047|PT|278.4|ICD9CM|Hypervitaminosis D|Hypervitaminosis D
C1442839|T047|AB|278.4|ICD9CM|Hypervitaminosis d|Hypervitaminosis d
C0029635|T047|AB|278.8|ICD9CM|Other hyperalimentation|Other hyperalimentation
C0029635|T047|PT|278.8|ICD9CM|Other hyperalimentation|Other hyperalimentation
C0041806|T047|HT|279|ICD9CM|Disorders involving the immune mechanism|Disorders involving the immune mechanism
C0522274|T047|HT|279.0|ICD9CM|Deficiency of humoral immunity|Deficiency of humoral immunity
C0086438|T047|AB|279.00|ICD9CM|Hypogammaglobulinem NOS|Hypogammaglobulinem NOS
C0086438|T047|PT|279.00|ICD9CM|Hypogammaglobulinemia, unspecified|Hypogammaglobulinemia, unspecified
C4049006|T047|AB|279.01|ICD9CM|Selective iga immunodef|Selective iga immunodef
C4049006|T047|PT|279.01|ICD9CM|Selective IgA immunodeficiency|Selective IgA immunodeficiency
C0154275|T046|AB|279.02|ICD9CM|Selective IgM immunodef|Selective IgM immunodef
C0154275|T046|PT|279.02|ICD9CM|Selective IgM immunodeficiency|Selective IgM immunodeficiency
C0154276|T047|PT|279.03|ICD9CM|Other selective immunoglobulin deficiencies|Other selective immunoglobulin deficiencies
C0154276|T047|AB|279.03|ICD9CM|Selective ig defic NEC|Selective ig defic NEC
C1457897|T047|AB|279.04|ICD9CM|Cong hypogammaglobulinem|Cong hypogammaglobulinem
C1457897|T047|PT|279.04|ICD9CM|Congenital hypogammaglobulinemia|Congenital hypogammaglobulinemia
C0740331|T047|AB|279.05|ICD9CM|Immunodefic w hyper-igm|Immunodefic w hyper-igm
C0740331|T047|PT|279.05|ICD9CM|Immunodeficiency with increased IgM|Immunodeficiency with increased IgM
C0009447|T047|AB|279.06|ICD9CM|Common variabl immunodef|Common variabl immunodef
C0009447|T047|PT|279.06|ICD9CM|Common variable immunodeficiency|Common variable immunodeficiency
C0522274|T047|AB|279.09|ICD9CM|Humoral immunity def NEC|Humoral immunity def NEC
C0522274|T047|PT|279.09|ICD9CM|Other deficiency of humoral immunity|Other deficiency of humoral immunity
C1533651|T046|HT|279.1|ICD9CM|Deficiency of cell-mediated immunity|Deficiency of cell-mediated immunity
C1608262|T046|AB|279.10|ICD9CM|Immundef t-cell def NOS|Immundef t-cell def NOS
C1608262|T046|PT|279.10|ICD9CM|Immunodeficiency with predominant T-cell defect, unspecified|Immunodeficiency with predominant T-cell defect, unspecified
C0012236|T047|AB|279.11|ICD9CM|Digeorge's syndrome|Digeorge's syndrome
C0012236|T047|PT|279.11|ICD9CM|Digeorge's syndrome|Digeorge's syndrome
C0043194|T047|AB|279.12|ICD9CM|Wiskott-aldrich syndrome|Wiskott-aldrich syndrome
C0043194|T047|PT|279.12|ICD9CM|Wiskott-aldrich syndrome|Wiskott-aldrich syndrome
C0152094|T047|AB|279.13|ICD9CM|Nezelof's syndrome|Nezelof's syndrome
C0152094|T047|PT|279.13|ICD9CM|Nezelof's syndrome|Nezelof's syndrome
C0154282|T047|AB|279.19|ICD9CM|Defic cell immunity NOS|Defic cell immunity NOS
C0154282|T047|PT|279.19|ICD9CM|Other deficiency of cell-mediated immunity|Other deficiency of cell-mediated immunity
C0494261|T047|AB|279.2|ICD9CM|Combined immunity defic|Combined immunity defic
C0494261|T047|PT|279.2|ICD9CM|Combined immunity deficiency|Combined immunity deficiency
C0021051|T047|AB|279.3|ICD9CM|Immunity deficiency NOS|Immunity deficiency NOS
C0021051|T047|PT|279.3|ICD9CM|Unspecified immunity deficiency|Unspecified immunity deficiency
C0687719|T047|HT|279.4|ICD9CM|Autoimmune disease, not elsewhere classified|Autoimmune disease, not elsewhere classified
C1328840|T047|AB|279.41|ICD9CM|Autoimmun lymphprof synd|Autoimmun lymphprof synd
C1328840|T047|PT|279.41|ICD9CM|Autoimmune lymphoproliferative syndrome|Autoimmune lymphoproliferative syndrome
C0687719|T047|AB|279.49|ICD9CM|Autoimmune disease NEC|Autoimmune disease NEC
C0687719|T047|PT|279.49|ICD9CM|Autoimmune disease, not elsewhere classified|Autoimmune disease, not elsewhere classified
C0018133|T047|HT|279.5|ICD9CM|Graft-versus-host disease|Graft-versus-host disease
C0018133|T047|PT|279.50|ICD9CM|Graft-versus-host disease, unspecified|Graft-versus-host disease, unspecified
C0018133|T047|AB|279.50|ICD9CM|Graft-versus-host NOS|Graft-versus-host NOS
C0856825|T047|AB|279.51|ICD9CM|Ac graft-versus-host dis|Ac graft-versus-host dis
C0856825|T047|PT|279.51|ICD9CM|Acute graft-versus-host disease|Acute graft-versus-host disease
C0867389|T047|AB|279.52|ICD9CM|Chronc graft-vs-host dis|Chronc graft-vs-host dis
C0867389|T047|PT|279.52|ICD9CM|Chronic graft-versus-host disease|Chronic graft-versus-host disease
C2349403|T047|AB|279.53|ICD9CM|Ac on chrn grft-vs-host|Ac on chrn grft-vs-host
C2349403|T047|PT|279.53|ICD9CM|Acute on chronic graft-versus-host disease|Acute on chronic graft-versus-host disease
C0398672|T047|AB|279.8|ICD9CM|Immune mechanism dis NEC|Immune mechanism dis NEC
C0398672|T047|PT|279.8|ICD9CM|Other specified disorders involving the immune mechanism|Other specified disorders involving the immune mechanism
C0041806|T047|AB|279.9|ICD9CM|Immune mechanism dis NOS|Immune mechanism dis NOS
C0041806|T047|PT|279.9|ICD9CM|Unspecified disorder of immune mechanism|Unspecified disorder of immune mechanism
C0162316|T047|HT|280|ICD9CM|Iron deficiency anemias|Iron deficiency anemias
C0018939|T047|HT|280-289.99|ICD9CM|DISEASES OF THE BLOOD AND BLOOD-FORMING ORGANS|DISEASES OF THE BLOOD AND BLOOD-FORMING ORGANS
C0154286|T047|AB|280.0|ICD9CM|Chr blood loss anemia|Chr blood loss anemia
C0154286|T047|PT|280.0|ICD9CM|Iron deficiency anemia secondary to blood loss (chronic)|Iron deficiency anemia secondary to blood loss (chronic)
C0154287|T047|AB|280.1|ICD9CM|Iron def anemia dietary|Iron def anemia dietary
C0154287|T047|PT|280.1|ICD9CM|Iron deficiency anemia secondary to inadequate dietary iron intake|Iron deficiency anemia secondary to inadequate dietary iron intake
C0029810|T047|AB|280.8|ICD9CM|Iron defic anemia NEC|Iron defic anemia NEC
C0029810|T047|PT|280.8|ICD9CM|Other specified iron deficiency anemias|Other specified iron deficiency anemias
C0162316|T047|AB|280.9|ICD9CM|Iron defic anemia NOS|Iron defic anemia NOS
C0162316|T047|PT|280.9|ICD9CM|Iron deficiency anemia, unspecified|Iron deficiency anemia, unspecified
C0154288|T047|HT|281|ICD9CM|Other deficiency anemias|Other deficiency anemias
C0002892|T047|AB|281.0|ICD9CM|Pernicious anemia|Pernicious anemia
C0002892|T047|PT|281.0|ICD9CM|Pernicious anemia|Pernicious anemia
C0154289|T047|AB|281.1|ICD9CM|B12 defic anemia NEC|B12 defic anemia NEC
C0154289|T047|PT|281.1|ICD9CM|Other vitamin B12 deficiency anemia|Other vitamin B12 deficiency anemia
C0151482|T047|AB|281.2|ICD9CM|Folate-deficiency anemia|Folate-deficiency anemia
C0151482|T047|PT|281.2|ICD9CM|Folate-deficiency anemia|Folate-deficiency anemia
C0302367|T047|AB|281.3|ICD9CM|Megaloblastic anemia NEC|Megaloblastic anemia NEC
C0302367|T047|PT|281.3|ICD9CM|Other specified megaloblastic anemias not elsewhere classified|Other specified megaloblastic anemias not elsewhere classified
C0154290|T047|AB|281.4|ICD9CM|Protein defic anemia|Protein defic anemia
C0154290|T047|PT|281.4|ICD9CM|Protein-deficiency anemia|Protein-deficiency anemia
C0154291|T047|PT|281.8|ICD9CM|Anemia associated with other specified nutritional deficiency|Anemia associated with other specified nutritional deficiency
C0154291|T047|AB|281.8|ICD9CM|Nutritional anemia NEC|Nutritional anemia NEC
C0041782|T047|AB|281.9|ICD9CM|Deficiency anemia NOS|Deficiency anemia NOS
C0041782|T047|PT|281.9|ICD9CM|Unspecified deficiency anemia|Unspecified deficiency anemia
C0002881|T047|HT|282|ICD9CM|Hereditary hemolytic anemias|Hereditary hemolytic anemias
C0037889|T047|AB|282.0|ICD9CM|Hereditary spherocytosis|Hereditary spherocytosis
C0037889|T047|PT|282.0|ICD9CM|Hereditary spherocytosis|Hereditary spherocytosis
C0013902|T047|AB|282.1|ICD9CM|Heredit elliptocytosis|Heredit elliptocytosis
C0013902|T047|PT|282.1|ICD9CM|Hereditary elliptocytosis|Hereditary elliptocytosis
C0002899|T047|PT|282.2|ICD9CM|Anemias due to disorders of glutathione metabolism|Anemias due to disorders of glutathione metabolism
C0002899|T047|AB|282.2|ICD9CM|Glutathione dis anemia|Glutathione dis anemia
C0154292|T047|AB|282.3|ICD9CM|Enzyme defic anemia NEC|Enzyme defic anemia NEC
C0154292|T047|PT|282.3|ICD9CM|Other hemolytic anemias due to enzyme deficiency|Other hemolytic anemias due to enzyme deficiency
C0039730|T047|HT|282.4|ICD9CM|Thalassemias|Thalassemias
C0039730|T047|AB|282.40|ICD9CM|Thalassemia, unspecified|Thalassemia, unspecified
C0039730|T047|PT|282.40|ICD9CM|Thalassemia, unspecified|Thalassemia, unspecified
C1260393|T047|PT|282.41|ICD9CM|Sickle-cell thalassemia without crisis|Sickle-cell thalassemia without crisis
C1260393|T047|AB|282.41|ICD9CM|Thlasema Hb-S w/o crisis|Thlasema Hb-S w/o crisis
C1260395|T047|PT|282.42|ICD9CM|Sickle-cell thalassemia with crisis|Sickle-cell thalassemia with crisis
C1260395|T047|AB|282.42|ICD9CM|Thlassemia Hb-S w crisis|Thlassemia Hb-S w crisis
C0002312|T047|PT|282.43|ICD9CM|Alpha thalassemia|Alpha thalassemia
C0002312|T047|AB|282.43|ICD9CM|Alpha thalassemia|Alpha thalassemia
C0005283|T047|PT|282.44|ICD9CM|Beta thalassemia|Beta thalassemia
C0005283|T047|AB|282.44|ICD9CM|Beta thalassemia|Beta thalassemia
C0271985|T047|AB|282.45|ICD9CM|Delta-beta thalassemia|Delta-beta thalassemia
C0271985|T047|PT|282.45|ICD9CM|Delta-beta thalassemia|Delta-beta thalassemia
C0085578|T047|PT|282.46|ICD9CM|Thalassemia minor|Thalassemia minor
C0085578|T047|AB|282.46|ICD9CM|Thalassemia minor|Thalassemia minor
C0472777|T047|PT|282.47|ICD9CM|Hemoglobin E-beta thalassemia|Hemoglobin E-beta thalassemia
C0472777|T047|AB|282.47|ICD9CM|Hgb E-beta thalassemia|Hgb E-beta thalassemia
C0477306|T047|PT|282.49|ICD9CM|Other thalassemia|Other thalassemia
C0477306|T047|AB|282.49|ICD9CM|Thalassemia NEC|Thalassemia NEC
C0037054|T047|AB|282.5|ICD9CM|Sickle-cell trait|Sickle-cell trait
C0037054|T047|PT|282.5|ICD9CM|Sickle-cell trait|Sickle-cell trait
C0002895|T047|HT|282.6|ICD9CM|Sickle-cell disease|Sickle-cell disease
C0002895|T047|AB|282.60|ICD9CM|Sickle cell disease NOS|Sickle cell disease NOS
C0002895|T047|PT|282.60|ICD9CM|Sickle-cell disease, unspecified|Sickle-cell disease, unspecified
C0272078|T047|AB|282.61|ICD9CM|Hb-SS disease w/o crisis|Hb-SS disease w/o crisis
C0272078|T047|PT|282.61|ICD9CM|Hb-SS disease without crisis|Hb-SS disease without crisis
C0238425|T047|AB|282.62|ICD9CM|Hb-SS disease w crisis|Hb-SS disease w crisis
C0238425|T047|PT|282.62|ICD9CM|Hb-SS disease with crisis|Hb-SS disease with crisis
C0019034|T047|AB|282.63|ICD9CM|Hb-SS/hb-C dis w/o crsis|Hb-SS/hb-C dis w/o crsis
C0019034|T047|PT|282.63|ICD9CM|Sickle-cell/Hb-C disease without crisis|Sickle-cell/Hb-C disease without crisis
C1260398|T047|AB|282.64|ICD9CM|Hb-S/Hb-C dis w crisis|Hb-S/Hb-C dis w crisis
C1260398|T047|PT|282.64|ICD9CM|Sickle-cell/Hb-C disease with crisis|Sickle-cell/Hb-C disease with crisis
C1260401|T047|AB|282.68|ICD9CM|Hb-S dis w/o crisis NEC|Hb-S dis w/o crisis NEC
C1260401|T047|PT|282.68|ICD9CM|Other sickle-cell disease without crisis|Other sickle-cell disease without crisis
C1260673|T047|AB|282.69|ICD9CM|Hb-SS dis NEC w crisis|Hb-SS dis NEC w crisis
C1260673|T047|PT|282.69|ICD9CM|Other sickle-cell disease with crisis|Other sickle-cell disease with crisis
C0029632|T047|AB|282.7|ICD9CM|Hemoglobinopathies NEC|Hemoglobinopathies NEC
C0029632|T047|PT|282.7|ICD9CM|Other hemoglobinopathies|Other hemoglobinopathies
C0154296|T047|AB|282.8|ICD9CM|Hered hemolytic anem NEC|Hered hemolytic anem NEC
C0154296|T047|PT|282.8|ICD9CM|Other specified hereditary hemolytic anemias|Other specified hereditary hemolytic anemias
C0002881|T047|AB|282.9|ICD9CM|Hered hemolytic anem NOS|Hered hemolytic anem NOS
C0002881|T047|PT|282.9|ICD9CM|Hereditary hemolytic anemia, unspecified|Hereditary hemolytic anemia, unspecified
C0002879|T047|HT|283|ICD9CM|Acquired hemolytic anemias|Acquired hemolytic anemias
C0002880|T047|AB|283.0|ICD9CM|Autoimmun hemolytic anem|Autoimmun hemolytic anem
C0002880|T047|PT|283.0|ICD9CM|Autoimmune hemolytic anemias|Autoimmune hemolytic anemias
C0028283|T047|HT|283.1|ICD9CM|Non-autoimmune hemolytic anemias|Non-autoimmune hemolytic anemias
C0028283|T047|PT|283.10|ICD9CM|Non-autoimmune hemolytic anemia, unspecified|Non-autoimmune hemolytic anemia, unspecified
C0028283|T047|AB|283.10|ICD9CM|Nonauto hem anemia NOS|Nonauto hem anemia NOS
C0019061|T047|AB|283.11|ICD9CM|Hemolytic uremic synd|Hemolytic uremic synd
C0019061|T047|PT|283.11|ICD9CM|Hemolytic-uremic syndrome|Hemolytic-uremic syndrome
C0375155|T047|AB|283.19|ICD9CM|Oth nonauto hem anemia|Oth nonauto hem anemia
C0375155|T047|PT|283.19|ICD9CM|Other non-autoimmune hemolytic anemias|Other non-autoimmune hemolytic anemias
C0019049|T047|PT|283.2|ICD9CM|Hemoglobinuria due to hemolysis from external causes|Hemoglobinuria due to hemolysis from external causes
C0019049|T047|AB|283.2|ICD9CM|Hemolytic hemoglobinuria|Hemolytic hemoglobinuria
C0002879|T047|AB|283.9|ICD9CM|Acq hemolytic anemia NOS|Acq hemolytic anemia NOS
C0002879|T047|PT|283.9|ICD9CM|Acquired hemolytic anemia, unspecified|Acquired hemolytic anemia, unspecified
C1719323|T047|HT|284|ICD9CM|Aplastic anemia and other bone marrow failure syndromes|Aplastic anemia and other bone marrow failure syndromes
C0702159|T047|HT|284.0|ICD9CM|Constitutional aplastic anemia|Constitutional aplastic anemia
C1719319|T047|AB|284.01|ICD9CM|Constitution RBC aplasia|Constitution RBC aplasia
C1719319|T047|PT|284.01|ICD9CM|Constitutional red blood cell aplasia|Constitutional red blood cell aplasia
C1719322|T047|AB|284.09|ICD9CM|Const aplastc anemia NEC|Const aplastc anemia NEC
C1719322|T047|PT|284.09|ICD9CM|Other constitutional aplastic anemia|Other constitutional aplastic anemia
C0030312|T047|HT|284.1|ICD9CM|Pancytopenia|Pancytopenia
C3161073|T046|AB|284.11|ICD9CM|Antin chemo indcd pancyt|Antin chemo indcd pancyt
C3161073|T046|PT|284.11|ICD9CM|Antineoplastic chemotherapy induced pancytopenia|Antineoplastic chemotherapy induced pancytopenia
C3161074|T046|AB|284.12|ICD9CM|Oth drg indcd pancytopna|Oth drg indcd pancytopna
C3161074|T046|PT|284.12|ICD9CM|Other drug-induced pancytopenia|Other drug-induced pancytopenia
C3161075|T047|PT|284.19|ICD9CM|Other pancytopenia|Other pancytopenia
C3161075|T047|AB|284.19|ICD9CM|Other pancytopenia|Other pancytopenia
C0302112|T047|PT|284.2|ICD9CM|Myelophthisis|Myelophthisis
C0302112|T047|AB|284.2|ICD9CM|Myelophthisis|Myelophthisis
C0029745|T047|HT|284.8|ICD9CM|Other specified aplastic anemias|Other specified aplastic anemias
C0865240|T047|AB|284.81|ICD9CM|Red cell aplasia|Red cell aplasia
C0865240|T047|PT|284.81|ICD9CM|Red cell aplasia (acquired)(adult)(with thymoma)|Red cell aplasia (acquired)(adult)(with thymoma)
C1955746|T047|AB|284.89|ICD9CM|Aplastic anemias NEC|Aplastic anemias NEC
C1955746|T047|PT|284.89|ICD9CM|Other specified aplastic anemias|Other specified aplastic anemias
C0002874|T047|AB|284.9|ICD9CM|Aplastic anemia NOS|Aplastic anemia NOS
C0002874|T047|PT|284.9|ICD9CM|Aplastic anemia, unspecified|Aplastic anemia, unspecified
C0472702|T047|HT|285|ICD9CM|Other and unspecified anemias|Other and unspecified anemias
C0002896|T047|AB|285.0|ICD9CM|Sideroblastic anemia|Sideroblastic anemia
C0002896|T047|PT|285.0|ICD9CM|Sideroblastic anemia|Sideroblastic anemia
C0154298|T047|AB|285.1|ICD9CM|Ac posthemorrhag anemia|Ac posthemorrhag anemia
C0154298|T047|PT|285.1|ICD9CM|Acute posthemorrhagic anemia|Acute posthemorrhagic anemia
C0002873|T047|HT|285.2|ICD9CM|Anemia of chronic disease|Anemia of chronic disease
C1561828|T047|AB|285.21|ICD9CM|Anemia in chr kidney dis|Anemia in chr kidney dis
C1561828|T047|PT|285.21|ICD9CM|Anemia in chronic kidney disease|Anemia in chronic kidney disease
C0475534|T047|AB|285.22|ICD9CM|Anemia in neoplastic dis|Anemia in neoplastic dis
C0475534|T047|PT|285.22|ICD9CM|Anemia in neoplastic disease|Anemia in neoplastic disease
C1719324|T047|PT|285.29|ICD9CM|Anemia of other chronic disease|Anemia of other chronic disease
C1719324|T047|AB|285.29|ICD9CM|Anemia-other chronic dis|Anemia-other chronic dis
C2712646|T047|AB|285.3|ICD9CM|Anemia d/t antineo chemo|Anemia d/t antineo chemo
C2712646|T047|PT|285.3|ICD9CM|Antineoplastic chemotherapy induced anemia|Antineoplastic chemotherapy induced anemia
C0029744|T047|AB|285.8|ICD9CM|Anemia NEC|Anemia NEC
C0029744|T047|PT|285.8|ICD9CM|Other specified anemias|Other specified anemias
C0002871|T047|AB|285.9|ICD9CM|Anemia NOS|Anemia NOS
C0002871|T047|PT|285.9|ICD9CM|Anemia, unspecified|Anemia, unspecified
C0005779|T047|HT|286|ICD9CM|Coagulation defects|Coagulation defects
C0019069|T047|AB|286.0|ICD9CM|Cong factor viii diord|Cong factor viii diord
C0019069|T047|PT|286.0|ICD9CM|Congenital factor VIII disorder|Congenital factor VIII disorder
C0008533|T047|AB|286.1|ICD9CM|Cong factor IX disorder|Cong factor IX disorder
C0008533|T047|PT|286.1|ICD9CM|Congenital factor IX disorder|Congenital factor IX disorder
C0015523|T047|AB|286.2|ICD9CM|Cong factor xi disorder|Cong factor xi disorder
C0015523|T047|PT|286.2|ICD9CM|Congenital factor XI deficiency|Congenital factor XI deficiency
C0009699|T047|AB|286.3|ICD9CM|Cong def clot factor NEC|Cong def clot factor NEC
C0009699|T047|PT|286.3|ICD9CM|Congenital deficiency of other clotting factors|Congenital deficiency of other clotting factors
C0042974|T047|PT|286.4|ICD9CM|Von Willebrand's disease|Von Willebrand's disease
C0042974|T047|AB|286.4|ICD9CM|Von willebrand's disease|Von willebrand's disease
C3648917|T047|HT|286.5|ICD9CM|Hemorrhagic disorder due to intrinsic circulating anticoagulants, antibodies, or inhibitors|Hemorrhagic disorder due to intrinsic circulating anticoagulants, antibodies, or inhibitors
C1096116|T047|AB|286.52|ICD9CM|Acquired hemophilia|Acquired hemophilia
C1096116|T047|PT|286.52|ICD9CM|Acquired hemophilia|Acquired hemophilia
C3161076|T047|PT|286.53|ICD9CM|Antiphospholipid antibody with hemorrhagic disorder|Antiphospholipid antibody with hemorrhagic disorder
C3161076|T047|AB|286.53|ICD9CM|Antiphospholipid w hemor|Antiphospholipid w hemor
C3161077|T047|AB|286.59|ICD9CM|Ot hem d/t circ anticoag|Ot hem d/t circ anticoag
C3161077|T047|PT|286.59|ICD9CM|Other hemorrhagic disorder due to intrinsic circulating anticoagulants, antibodies, or inhibitors|Other hemorrhagic disorder due to intrinsic circulating anticoagulants, antibodies, or inhibitors
C0012739|T047|AB|286.6|ICD9CM|Defibrination syndrome|Defibrination syndrome
C0012739|T047|PT|286.6|ICD9CM|Defibrination syndrome|Defibrination syndrome
C0001169|T047|AB|286.7|ICD9CM|Acq coagul factor defic|Acq coagul factor defic
C0001169|T047|PT|286.7|ICD9CM|Acquired coagulation factor deficiency|Acquired coagulation factor deficiency
C0029496|T047|AB|286.9|ICD9CM|Coagulat defect NEC/NOS|Coagulat defect NEC/NOS
C0029496|T047|PT|286.9|ICD9CM|Other and unspecified coagulation defects|Other and unspecified coagulation defects
C0154300|T047|HT|287|ICD9CM|Purpura and other hemorrhagic conditions|Purpura and other hemorrhagic conditions
C0034152|T047|AB|287.0|ICD9CM|Allergic purpura|Allergic purpura
C0034152|T047|PT|287.0|ICD9CM|Allergic purpura|Allergic purpura
C0235604|T047|PT|287.1|ICD9CM|Qualitative platelet defects|Qualitative platelet defects
C0235604|T047|AB|287.1|ICD9CM|Thrombocytopathy|Thrombocytopathy
C0029678|T047|PT|287.2|ICD9CM|Other nonthrombocytopenic purpuras|Other nonthrombocytopenic purpuras
C0029678|T047|AB|287.2|ICD9CM|Purpura NOS|Purpura NOS
C0701157|T047|HT|287.3|ICD9CM|Primary thrombocytopenia|Primary thrombocytopenia
C1561830|T047|AB|287.30|ICD9CM|Prim thrombocytopen NOS|Prim thrombocytopen NOS
C1561830|T047|PT|287.30|ICD9CM|Primary thrombocytopenia,unspecified|Primary thrombocytopenia,unspecified
C0398650|T047|AB|287.31|ICD9CM|Immune thrombocyt purpra|Immune thrombocyt purpra
C0398650|T047|PT|287.31|ICD9CM|Immune thrombocytopenic purpura|Immune thrombocytopenic purpura
C0272126|T047|AB|287.32|ICD9CM|Evans' syndrome|Evans' syndrome
C0272126|T047|PT|287.32|ICD9CM|Evans' syndrome|Evans' syndrome
C1561831|T047|AB|287.33|ICD9CM|Cong/herid thromb purpra|Cong/herid thromb purpra
C1561831|T047|PT|287.33|ICD9CM|Congenital and hereditary thrombocytopenic purpura|Congenital and hereditary thrombocytopenic purpura
C0477317|T047|PT|287.39|ICD9CM|Other primary thrombocytopenia|Other primary thrombocytopenia
C0477317|T047|AB|287.39|ICD9CM|Prim thrombocytopen NEC|Prim thrombocytopen NEC
C0154301|T047|HT|287.4|ICD9CM|Secondary thrombocytopenia|Secondary thrombocytopenia
C0398648|T046|PT|287.41|ICD9CM|Posttransfusion purpura|Posttransfusion purpura
C0398648|T046|AB|287.41|ICD9CM|Posttransfusion purpura|Posttransfusion purpura
C2921026|T047|PT|287.49|ICD9CM|Other secondary thrombocytopenia|Other secondary thrombocytopenia
C2921026|T047|AB|287.49|ICD9CM|Sec thrombocytpenia NEC|Sec thrombocytpenia NEC
C0040034|T047|AB|287.5|ICD9CM|Thrombocytopenia NOS|Thrombocytopenia NOS
C0040034|T047|PT|287.5|ICD9CM|Thrombocytopenia, unspecified|Thrombocytopenia, unspecified
C0029804|T046|AB|287.8|ICD9CM|Hemorrhagic cond NEC|Hemorrhagic cond NEC
C0029804|T046|PT|287.8|ICD9CM|Other specified hemorrhagic conditions|Other specified hemorrhagic conditions
C0019087|T047|AB|287.9|ICD9CM|Hemorrhagic cond NOS|Hemorrhagic cond NOS
C0019087|T047|PT|287.9|ICD9CM|Unspecified hemorrhagic conditions|Unspecified hemorrhagic conditions
C0023510|T047|HT|288|ICD9CM|Diseases of white blood cells|Diseases of white blood cells
C0027947|T047|HT|288.0|ICD9CM|Neutropenia|Neutropenia
C0027947|T047|AB|288.00|ICD9CM|Neutropenia NOS|Neutropenia NOS
C0027947|T047|PT|288.00|ICD9CM|Neutropenia, unspecified|Neutropenia, unspecified
C0340970|T019|PT|288.01|ICD9CM|Congenital neutropenia|Congenital neutropenia
C0340970|T019|AB|288.01|ICD9CM|Congenital neutropenia|Congenital neutropenia
C0221023|T047|PT|288.02|ICD9CM|Cyclic neutropenia|Cyclic neutropenia
C0221023|T047|AB|288.02|ICD9CM|Cyclic neutropenia|Cyclic neutropenia
C0272178|T047|PT|288.03|ICD9CM|Drug induced neutropenia|Drug induced neutropenia
C0272178|T047|AB|288.03|ICD9CM|Drug induced neutropenia|Drug induced neutropenia
C0272181|T047|AB|288.04|ICD9CM|Neutropenia d/t infectn|Neutropenia d/t infectn
C0272181|T047|PT|288.04|ICD9CM|Neutropenia due to infection|Neutropenia due to infection
C2873812|T047|AB|288.09|ICD9CM|Neutropenia NEC|Neutropenia NEC
C2873812|T047|PT|288.09|ICD9CM|Other neutropenia|Other neutropenia
C0016808|T047|AB|288.1|ICD9CM|Function dis neutrophils|Function dis neutrophils
C0016808|T047|PT|288.1|ICD9CM|Functional disorders of polymorphonuclear neutrophils|Functional disorders of polymorphonuclear neutrophils
C0017377|T047|PT|288.2|ICD9CM|Genetic anomalies of leukocytes|Genetic anomalies of leukocytes
C0017377|T047|AB|288.2|ICD9CM|Genetic anomaly leukocyt|Genetic anomaly leukocyt
C0014457|T047|AB|288.3|ICD9CM|Eosinophilia|Eosinophilia
C0014457|T047|PT|288.3|ICD9CM|Eosinophilia|Eosinophilia
C3887558|T047|AB|288.4|ICD9CM|Hemophagocytic syndromes|Hemophagocytic syndromes
C3887558|T047|PT|288.4|ICD9CM|Hemophagocytic syndromes|Hemophagocytic syndromes
C0750394|T033|HT|288.5|ICD9CM|Decreased white blood cell count|Decreased white blood cell count
C0023530|T047|AB|288.50|ICD9CM|Leukocytopenia NOS|Leukocytopenia NOS
C0023530|T047|PT|288.50|ICD9CM|Leukocytopenia, unspecified|Leukocytopenia, unspecified
C0024312|T047|PT|288.51|ICD9CM|Lymphocytopenia|Lymphocytopenia
C0024312|T047|AB|288.51|ICD9CM|Lymphocytopenia|Lymphocytopenia
C1719330|T047|AB|288.59|ICD9CM|Decreased WBC count NEC|Decreased WBC count NEC
C1719330|T047|PT|288.59|ICD9CM|Other decreased white blood cell count|Other decreased white blood cell count
C0750426|T033|HT|288.6|ICD9CM|Elevated white blood cell count|Elevated white blood cell count
C0023518|T047|AB|288.60|ICD9CM|Leukocytosis NOS|Leukocytosis NOS
C0023518|T047|PT|288.60|ICD9CM|Leukocytosis, unspecified|Leukocytosis, unspecified
C1719337|T047|PT|288.61|ICD9CM|Lymphocytosis (symptomatic)|Lymphocytosis (symptomatic)
C1719337|T047|AB|288.61|ICD9CM|Lymphocytosis-symptomatc|Lymphocytosis-symptomatc
C0023501|T047|PT|288.62|ICD9CM|Leukemoid reaction|Leukemoid reaction
C0023501|T047|AB|288.62|ICD9CM|Leukemoid reaction|Leukemoid reaction
C1719340|T047|PT|288.63|ICD9CM|Monocytosis (symptomatic)|Monocytosis (symptomatic)
C1719340|T047|AB|288.63|ICD9CM|Monocytosis-symptomatic|Monocytosis-symptomatic
C0085663|T047|PT|288.64|ICD9CM|Plasmacytosis|Plasmacytosis
C0085663|T047|AB|288.64|ICD9CM|Plasmacytosis|Plasmacytosis
C0702266|T047|PT|288.65|ICD9CM|Basophilia|Basophilia
C0702266|T047|AB|288.65|ICD9CM|Basophilia|Basophilia
C0741439|T047|PT|288.66|ICD9CM|Bandemia|Bandemia
C0741439|T047|AB|288.66|ICD9CM|Bandemia|Bandemia
C1719341|T047|AB|288.69|ICD9CM|Elevated WBC count NEC|Elevated WBC count NEC
C1719341|T047|PT|288.69|ICD9CM|Other elevated white blood cell count|Other elevated white blood cell count
C0477318|T047|PT|288.8|ICD9CM|Other specified disease of white blood cells|Other specified disease of white blood cells
C0477318|T047|AB|288.8|ICD9CM|Wbc disease NEC|Wbc disease NEC
C0023510|T047|PT|288.9|ICD9CM|Unspecified disease of white blood cells|Unspecified disease of white blood cells
C0023510|T047|AB|288.9|ICD9CM|Wbc disease NOS|Wbc disease NOS
C0451639|T047|HT|289|ICD9CM|Other diseases of blood and blood-forming organs|Other diseases of blood and blood-forming organs
C1318533|T047|PT|289.0|ICD9CM|Polycythemia, secondary|Polycythemia, secondary
C1318533|T047|AB|289.0|ICD9CM|Secondary polycythemia|Secondary polycythemia
C0154304|T047|AB|289.1|ICD9CM|Chronic lymphadenitis|Chronic lymphadenitis
C0154304|T047|PT|289.1|ICD9CM|Chronic lymphadenitis|Chronic lymphadenitis
C0025469|T047|AB|289.2|ICD9CM|Mesenteric lymphadenitis|Mesenteric lymphadenitis
C0025469|T047|PT|289.2|ICD9CM|Nonspecific mesenteric lymphadenitis|Nonspecific mesenteric lymphadenitis
C0024207|T047|AB|289.3|ICD9CM|Lymphadenitis NOS|Lymphadenitis NOS
C0024207|T047|PT|289.3|ICD9CM|Lymphadenitis, unspecified, except mesenteric|Lymphadenitis, unspecified, except mesenteric
C0020532|T047|AB|289.4|ICD9CM|Hypersplenism|Hypersplenism
C0020532|T047|PT|289.4|ICD9CM|Hypersplenism|Hypersplenism
C0154305|T047|HT|289.5|ICD9CM|Other diseases of spleen|Other diseases of spleen
C0037997|T047|PT|289.50|ICD9CM|Disease of spleen, unspecified|Disease of spleen, unspecified
C0037997|T047|AB|289.50|ICD9CM|Spleen disease NOS|Spleen disease NOS
C0398661|T047|AB|289.51|ICD9CM|Chr congest splenomegaly|Chr congest splenomegaly
C0398661|T047|PT|289.51|ICD9CM|Chronic congestive splenomegaly|Chronic congestive splenomegaly
C1260402|T047|AB|289.52|ICD9CM|Splenic sequestration|Splenic sequestration
C1260402|T047|PT|289.52|ICD9CM|Splenic sequestration|Splenic sequestration
C0398580|T047|PT|289.53|ICD9CM|Neutropenic splenomegaly|Neutropenic splenomegaly
C0398580|T047|AB|289.53|ICD9CM|Neutropenic splenomegaly|Neutropenic splenomegaly
C0154305|T047|PT|289.59|ICD9CM|Other diseases of spleen|Other diseases of spleen
C0154305|T047|AB|289.59|ICD9CM|Spleen disease NEC|Spleen disease NEC
C0152264|T047|AB|289.6|ICD9CM|Familial polycythemia|Familial polycythemia
C0152264|T047|PT|289.6|ICD9CM|Familial polycythemia|Familial polycythemia
C0025637|T047|AB|289.7|ICD9CM|Methemoglobinemia|Methemoglobinemia
C0025637|T047|PT|289.7|ICD9CM|Methemoglobinemia|Methemoglobinemia
C0029768|T047|HT|289.8|ICD9CM|Other specified diseases of blood and blood-forming organs|Other specified diseases of blood and blood-forming organs
C1260404|T047|AB|289.81|ICD9CM|Prim hypercoagulable st|Prim hypercoagulable st
C1260404|T047|PT|289.81|ICD9CM|Primary hypercoagulable state|Primary hypercoagulable state
C1456282|T047|AB|289.82|ICD9CM|Sec hypercoagulable st|Sec hypercoagulable st
C1456282|T047|PT|289.82|ICD9CM|Secondary hypercoagulable state|Secondary hypercoagulable state
C0026987|T191|PT|289.83|ICD9CM|Myelofibrosis|Myelofibrosis
C0026987|T191|AB|289.83|ICD9CM|Myelofibrosis|Myelofibrosis
C0272285|T047|AB|289.84|ICD9CM|Heparin-indu thrombocyto|Heparin-indu thrombocyto
C0272285|T047|PT|289.84|ICD9CM|Heparin-induced thrombocytopenia (HIT)|Heparin-induced thrombocytopenia (HIT)
C0029768|T047|AB|289.89|ICD9CM|Blood diseases NEC|Blood diseases NEC
C0029768|T047|PT|289.89|ICD9CM|Other specified diseases of blood and blood-forming organs|Other specified diseases of blood and blood-forming organs
C0018939|T047|AB|289.9|ICD9CM|Blood disease NOS|Blood disease NOS
C0018939|T047|PT|289.9|ICD9CM|Unspecified diseases of blood and blood-forming organs|Unspecified diseases of blood and blood-forming organs
C0497327|T048|HT|290|ICD9CM|Dementias|Dementias
C0520473|T048|HT|290-294.99|ICD9CM|ORGANIC PSYCHOTIC CONDITIONS|ORGANIC PSYCHOTIC CONDITIONS
C0033975|T048|HT|290-299.99|ICD9CM|PSYCHOSES|PSYCHOSES
C3161379|T048|HT|290-319.99|ICD9CM|MENTAL, BEHAVIORAL AND NEURODEVELOPMENTAL DISORDERS|MENTAL, BEHAVIORAL AND NEURODEVELOPMENTAL DISORDERS
C3665587|T048|AB|290.0|ICD9CM|Senile dementia uncomp|Senile dementia uncomp
C3665587|T048|PT|290.0|ICD9CM|Senile dementia, uncomplicated|Senile dementia, uncomplicated
C0011265|T048|HT|290.1|ICD9CM|Presenile dementia|Presenile dementia
C0677545|T048|AB|290.10|ICD9CM|Presenile dementia|Presenile dementia
C0677545|T048|PT|290.10|ICD9CM|Presenile dementia, uncomplicated|Presenile dementia, uncomplicated
C0154309|T048|AB|290.11|ICD9CM|Presenile delirium|Presenile delirium
C0154309|T048|PT|290.11|ICD9CM|Presenile dementia with delirium|Presenile dementia with delirium
C0154310|T048|AB|290.12|ICD9CM|Presenile delusion|Presenile delusion
C0154310|T048|PT|290.12|ICD9CM|Presenile dementia with delusional features|Presenile dementia with delusional features
C0338629|T048|PT|290.13|ICD9CM|Presenile dementia with depressive features|Presenile dementia with depressive features
C0338629|T048|AB|290.13|ICD9CM|Presenile depression|Presenile depression
C0859643|T048|HT|290.2|ICD9CM|Senile dementia with delusional or depressive features|Senile dementia with delusional or depressive features
C1269750|T048|AB|290.20|ICD9CM|Senile delusion|Senile delusion
C1269750|T048|PT|290.20|ICD9CM|Senile dementia with delusional features|Senile dementia with delusional features
C0338631|T048|PT|290.21|ICD9CM|Senile dementia with depressive features|Senile dementia with depressive features
C0338631|T048|AB|290.21|ICD9CM|Senile depressive|Senile depressive
C0154315|T048|AB|290.3|ICD9CM|Senile delirium|Senile delirium
C0154315|T048|PT|290.3|ICD9CM|Senile dementia with delirium|Senile dementia with delirium
C0011269|T047|HT|290.4|ICD9CM|Vascular dementia|Vascular dementia
C0236650|T048|PT|290.40|ICD9CM|Vascular dementia, uncomplicated|Vascular dementia, uncomplicated
C0236650|T048|AB|290.40|ICD9CM|Vascular dementia,uncomp|Vascular dementia,uncomp
C0236651|T048|AB|290.41|ICD9CM|Vasc dementia w delirium|Vasc dementia w delirium
C0236651|T048|PT|290.41|ICD9CM|Vascular dementia, with delirium|Vascular dementia, with delirium
C0236652|T048|AB|290.42|ICD9CM|Vasc dementia w delusion|Vasc dementia w delusion
C0236652|T048|PT|290.42|ICD9CM|Vascular dementia, with delusions|Vascular dementia, with delusions
C0236653|T048|AB|290.43|ICD9CM|Vasc dementia w depressn|Vasc dementia w depressn
C0236653|T048|PT|290.43|ICD9CM|Vascular dementia, with depressed mood|Vascular dementia, with depressed mood
C0154319|T048|PT|290.8|ICD9CM|Other specified senile psychotic conditions|Other specified senile psychotic conditions
C0154319|T048|AB|290.8|ICD9CM|Senile psychosis NEC|Senile psychosis NEC
C1457889|T048|AB|290.9|ICD9CM|Senile psychot cond NOS|Senile psychot cond NOS
C1457889|T048|PT|290.9|ICD9CM|Unspecified senile psychotic condition|Unspecified senile psychotic condition
C1456285|T048|HT|291|ICD9CM|Alcohol-induced mental disorders|Alcohol-induced mental disorders
C0001957|T047|PT|291.0|ICD9CM|Alcohol withdrawal delirium|Alcohol withdrawal delirium
C0001957|T047|AB|291.0|ICD9CM|Delirium tremens|Delirium tremens
C0001940|T048|AB|291.1|ICD9CM|Alcohol amnestic disordr|Alcohol amnestic disordr
C0001940|T048|PT|291.1|ICD9CM|Alcohol-induced persisting amnestic disorder|Alcohol-induced persisting amnestic disorder
C0236656|T048|AB|291.2|ICD9CM|Alcohol persist dementia|Alcohol persist dementia
C0236656|T048|PT|291.2|ICD9CM|Alcohol-induced persisting dementia|Alcohol-induced persisting dementia
C0302369|T047|AB|291.3|ICD9CM|Alcoh psy dis w hallucin|Alcoh psy dis w hallucin
C0302369|T047|PT|291.3|ICD9CM|Alcohol-induced psychotic disorder with hallucinations|Alcohol-induced psychotic disorder with hallucinations
C0001950|T048|PT|291.4|ICD9CM|Idiosyncratic alcohol intoxication|Idiosyncratic alcohol intoxication
C0001950|T048|AB|291.4|ICD9CM|Pathologic alcohol intox|Pathologic alcohol intox
C0236658|T048|AB|291.5|ICD9CM|Alcoh psych dis w delus|Alcoh psych dis w delus
C0236658|T048|PT|291.5|ICD9CM|Alcohol-induced psychotic disorder with delusions|Alcohol-induced psychotic disorder with delusions
C1456283|T048|HT|291.8|ICD9CM|Other specified alcohol-induced mental disorders|Other specified alcohol-induced mental disorders
C0236663|T047|AB|291.81|ICD9CM|Alcohol withdrawal|Alcohol withdrawal
C0236663|T047|PT|291.81|ICD9CM|Alcohol withdrawal|Alcohol withdrawal
C0236662|T048|AB|291.82|ICD9CM|Alcoh induce sleep disor|Alcoh induce sleep disor
C0236662|T048|PT|291.82|ICD9CM|Alcohol induced sleep disorders|Alcohol induced sleep disorders
C1456283|T048|AB|291.89|ICD9CM|Alcohol mental disor NEC|Alcohol mental disor NEC
C1456283|T048|PT|291.89|ICD9CM|Other alcohol-induced mental disorders|Other alcohol-induced mental disorders
C0033936|T048|AB|291.9|ICD9CM|Alcohol mental disor NOS|Alcohol mental disor NOS
C0033936|T048|PT|291.9|ICD9CM|Unspecified alcohol-induced mental disorders|Unspecified alcohol-induced mental disorders
C0154330|T048|HT|292|ICD9CM|Drug-induced mental disorders|Drug-induced mental disorders
C0152128|T047|AB|292.0|ICD9CM|Drug withdrawal|Drug withdrawal
C0152128|T047|PT|292.0|ICD9CM|Drug withdrawal|Drug withdrawal
C0033937|T048|HT|292.1|ICD9CM|Drug-induced psychotic disorders|Drug-induced psychotic disorders
C1456286|T048|AB|292.11|ICD9CM|Drug psych disor w delus|Drug psych disor w delus
C1456286|T048|PT|292.11|ICD9CM|Drug-induced psychotic disorder with delusions|Drug-induced psychotic disorder with delusions
C1456732|T048|AB|292.12|ICD9CM|Drug psy dis w hallucin|Drug psy dis w hallucin
C1456732|T048|PT|292.12|ICD9CM|Drug-induced psychotic disorder with hallucinations|Drug-induced psychotic disorder with hallucinations
C0152129|T037|AB|292.2|ICD9CM|Pathologic drug intox|Pathologic drug intox
C0152129|T037|PT|292.2|ICD9CM|Pathological drug intoxication|Pathological drug intoxication
C0154325|T048|HT|292.8|ICD9CM|Other specified drug-induced mental disorders|Other specified drug-induced mental disorders
C0154326|T048|AB|292.81|ICD9CM|Drug-induced delirium|Drug-induced delirium
C0154326|T048|PT|292.81|ICD9CM|Drug-induced delirium|Drug-induced delirium
C1456288|T048|AB|292.82|ICD9CM|Drug persisting dementia|Drug persisting dementia
C1456288|T048|PT|292.82|ICD9CM|Drug-induced persisting dementia|Drug-induced persisting dementia
C1456289|T047|AB|292.83|ICD9CM|Drug persist amnestc dis|Drug persist amnestc dis
C1456289|T047|PT|292.83|ICD9CM|Drug-induced persisting amnestic disorder|Drug-induced persisting amnestic disorder
C1998428|T048|AB|292.84|ICD9CM|Drug-induced mood disord|Drug-induced mood disord
C1998428|T048|PT|292.84|ICD9CM|Drug-induced mood disorder|Drug-induced mood disorder
C1456292|T048|AB|292.85|ICD9CM|Drug induced sleep disor|Drug induced sleep disor
C1456292|T048|PT|292.85|ICD9CM|Drug induced sleep disorders|Drug induced sleep disorders
C0154325|T048|AB|292.89|ICD9CM|Drug mental disorder NEC|Drug mental disorder NEC
C0154325|T048|PT|292.89|ICD9CM|Other specified drug-induced mental disorders|Other specified drug-induced mental disorders
C0154330|T048|AB|292.9|ICD9CM|Drug mental disorder NOS|Drug mental disorder NOS
C0154330|T048|PT|292.9|ICD9CM|Unspecified drug-induced mental disorder|Unspecified drug-induced mental disorder
C1456303|T048|HT|293|ICD9CM|Transient mental disorders due to conditions classified elsewhere|Transient mental disorders due to conditions classified elsewhere
C1456296|T048|AB|293.0|ICD9CM|Delirium d/t other cond|Delirium d/t other cond
C1456296|T048|PT|293.0|ICD9CM|Delirium due to conditions classified elsewhere|Delirium due to conditions classified elsewhere
C0154333|T048|AB|293.1|ICD9CM|Subacute delirium|Subacute delirium
C0154333|T048|PT|293.1|ICD9CM|Subacute delirium|Subacute delirium
C1456301|T048|HT|293.8|ICD9CM|Other specified transient mental disorders due to conditions classified elsewhere|Other specified transient mental disorders due to conditions classified elsewhere
C1456297|T048|AB|293.81|ICD9CM|Psy dis w delus oth dis|Psy dis w delus oth dis
C1456297|T048|PT|293.81|ICD9CM|Psychotic disorder with delusions in conditions classified elsewhere|Psychotic disorder with delusions in conditions classified elsewhere
C0029226|T048|AB|293.82|ICD9CM|Psy dis w halluc oth dis|Psy dis w halluc oth dis
C0029226|T048|PT|293.82|ICD9CM|Psychotic disorder with hallucinations in conditions classified elsewhere|Psychotic disorder with hallucinations in conditions classified elsewhere
C1456298|T048|PT|293.83|ICD9CM|Mood disorder in conditions classified elsewhere|Mood disorder in conditions classified elsewhere
C1456298|T048|AB|293.83|ICD9CM|Mood disorder other dis|Mood disorder other dis
C1456299|T048|PT|293.84|ICD9CM|Anxiety disorder in conditions classified elsewhere|Anxiety disorder in conditions classified elsewhere
C1456299|T048|AB|293.84|ICD9CM|Anxiety disorder oth dis|Anxiety disorder oth dis
C0154334|T048|PT|293.89|ICD9CM|Other specified transient mental disorders due to conditions classified elsewhere, other|Other specified transient mental disorders due to conditions classified elsewhere, other
C0154334|T048|AB|293.89|ICD9CM|Transient mental dis NEC|Transient mental dis NEC
C1456302|T048|AB|293.9|ICD9CM|Transient mental dis NOS|Transient mental dis NOS
C1456302|T048|PT|293.9|ICD9CM|Unspecified transient mental disorder in conditions classified elsewhere|Unspecified transient mental disorder in conditions classified elsewhere
C0154336|T048|HT|294|ICD9CM|Persistent mental disorders due to conditions classified elsewhere|Persistent mental disorders due to conditions classified elsewhere
C0002625|T048|AB|294.0|ICD9CM|Amnestic disord oth dis|Amnestic disord oth dis
C0002625|T048|PT|294.0|ICD9CM|Amnestic disorder in conditions classified elsewhere|Amnestic disorder in conditions classified elsewhere
C0338632|T048|HT|294.1|ICD9CM|Dementia in conditions classified elsewhere|Dementia in conditions classified elsewhere
C0878691|T047|PT|294.10|ICD9CM|Dementia in conditions classified elsewhere without behavioral disturbance|Dementia in conditions classified elsewhere without behavioral disturbance
C0878691|T047|AB|294.10|ICD9CM|Dementia w/o behav dist|Dementia w/o behav dist
C0878692|T047|PT|294.11|ICD9CM|Dementia in conditions classified elsewhere with behavioral disturbance|Dementia in conditions classified elsewhere with behavioral disturbance
C0878692|T047|AB|294.11|ICD9CM|Dementia w behavior dist|Dementia w behavior dist
C0497327|T048|HT|294.2|ICD9CM|Dementia, unspecified|Dementia, unspecified
C3161078|T048|AB|294.20|ICD9CM|Demen NOS w/o behv dstrb|Demen NOS w/o behv dstrb
C3161078|T048|PT|294.20|ICD9CM|Dementia, unspecified, without behavioral disturbance|Dementia, unspecified, without behavioral disturbance
C3161079|T048|AB|294.21|ICD9CM|Demen NOS w behav distrb|Demen NOS w behav distrb
C3161079|T048|PT|294.21|ICD9CM|Dementia, unspecified, with behavioral disturbance|Dementia, unspecified, with behavioral disturbance
C0154338|T048|AB|294.8|ICD9CM|Mental disor NEC oth dis|Mental disor NEC oth dis
C0154338|T048|PT|294.8|ICD9CM|Other persistent mental disorders due to conditions classified elsewhere|Other persistent mental disorders due to conditions classified elsewhere
C1456428|T048|AB|294.9|ICD9CM|Mental disor NOS oth dis|Mental disor NOS oth dis
C1456428|T048|PT|294.9|ICD9CM|Unspecified persistent mental disorders due to conditions classified elsewhere|Unspecified persistent mental disorders due to conditions classified elsewhere
C0036341|T048|HT|295|ICD9CM|Schizophrenic disorders|Schizophrenic disorders
C0497333|T048|HT|295-299.99|ICD9CM|OTHER PSYCHOSES|OTHER PSYCHOSES
C0221520|T048|HT|295.0|ICD9CM|Simple type schizophrenia|Simple type schizophrenia
C0221520|T048|AB|295.00|ICD9CM|Simpl schizophren-unspec|Simpl schizophren-unspec
C0221520|T048|PT|295.00|ICD9CM|Simple type schizophrenia, unspecified|Simple type schizophrenia, unspecified
C0154339|T048|AB|295.01|ICD9CM|Simpl schizophren-subchr|Simpl schizophren-subchr
C0154339|T048|PT|295.01|ICD9CM|Simple type schizophrenia, subchronic|Simple type schizophrenia, subchronic
C0154340|T048|AB|295.02|ICD9CM|Simple schizophren-chr|Simple schizophren-chr
C0154340|T048|PT|295.02|ICD9CM|Simple type schizophrenia, chronic|Simple type schizophrenia, chronic
C0154341|T048|AB|295.03|ICD9CM|Simp schiz-subchr/exacer|Simp schiz-subchr/exacer
C0154341|T048|PT|295.03|ICD9CM|Simple type schizophrenia, subchronic with acute exacerbation|Simple type schizophrenia, subchronic with acute exacerbation
C0154342|T048|AB|295.04|ICD9CM|Simpl schizo-chr/exacerb|Simpl schizo-chr/exacerb
C0154342|T048|PT|295.04|ICD9CM|Simple type schizophrenia, chronic with acute exacerbation|Simple type schizophrenia, chronic with acute exacerbation
C0154343|T048|AB|295.05|ICD9CM|Simpl schizophren-remiss|Simpl schizophren-remiss
C0154343|T048|PT|295.05|ICD9CM|Simple type schizophrenia, in remission|Simple type schizophrenia, in remission
C0036347|T048|HT|295.1|ICD9CM|Disorganized type schizophrenia|Disorganized type schizophrenia
C0375157|T048|PT|295.10|ICD9CM|Disorganized type schizophrenia, unspecified|Disorganized type schizophrenia, unspecified
C0375157|T048|AB|295.10|ICD9CM|Hebephrenia-unspec|Hebephrenia-unspec
C0154344|T048|PT|295.11|ICD9CM|Disorganized type schizophrenia, subchronic|Disorganized type schizophrenia, subchronic
C0154344|T048|AB|295.11|ICD9CM|Hebephrenia-subchronic|Hebephrenia-subchronic
C0154345|T048|PT|295.12|ICD9CM|Disorganized type schizophrenia, chronic|Disorganized type schizophrenia, chronic
C0154345|T048|AB|295.12|ICD9CM|Hebephrenia-chronic|Hebephrenia-chronic
C0154346|T048|PT|295.13|ICD9CM|Disorganized type schizophrenia, subchronic with acute exacerbation|Disorganized type schizophrenia, subchronic with acute exacerbation
C0154346|T048|AB|295.13|ICD9CM|Hebephren-subchr/exacerb|Hebephren-subchr/exacerb
C0154347|T048|PT|295.14|ICD9CM|Disorganized type schizophrenia, chronic with acute exacerbation|Disorganized type schizophrenia, chronic with acute exacerbation
C0154347|T048|AB|295.14|ICD9CM|Hebephrenia-chr/exacerb|Hebephrenia-chr/exacerb
C0270395|T048|PT|295.15|ICD9CM|Disorganized type schizophrenia, in remission|Disorganized type schizophrenia, in remission
C0270395|T048|AB|295.15|ICD9CM|Hebephrenia-remission|Hebephrenia-remission
C0036344|T048|HT|295.2|ICD9CM|Catatonic type schizophrenia|Catatonic type schizophrenia
C0375158|T048|AB|295.20|ICD9CM|Catatonia-unspec|Catatonia-unspec
C0375158|T048|PT|295.20|ICD9CM|Catatonic type schizophrenia, unspecified|Catatonic type schizophrenia, unspecified
C0154349|T048|AB|295.21|ICD9CM|Catatonia-subchronic|Catatonia-subchronic
C0154349|T048|PT|295.21|ICD9CM|Catatonic type schizophrenia, subchronic|Catatonic type schizophrenia, subchronic
C0154350|T048|AB|295.22|ICD9CM|Catatonia-chronic|Catatonia-chronic
C0154350|T048|PT|295.22|ICD9CM|Catatonic type schizophrenia, chronic|Catatonic type schizophrenia, chronic
C0154351|T048|AB|295.23|ICD9CM|Catatonia-subchr/exacerb|Catatonia-subchr/exacerb
C0154351|T048|PT|295.23|ICD9CM|Catatonic type schizophrenia, subchronic with acute exacerbation|Catatonic type schizophrenia, subchronic with acute exacerbation
C0154352|T048|AB|295.24|ICD9CM|Catatonia-chr/exacerb|Catatonia-chr/exacerb
C0154352|T048|PT|295.24|ICD9CM|Catatonic type schizophrenia, chronic with acute exacerbation|Catatonic type schizophrenia, chronic with acute exacerbation
C0270390|T048|AB|295.25|ICD9CM|Catatonia-remission|Catatonia-remission
C0270390|T048|PT|295.25|ICD9CM|Catatonic type schizophrenia, in remission|Catatonic type schizophrenia, in remission
C0036349|T048|HT|295.3|ICD9CM|Paranoid type schizophrenia|Paranoid type schizophrenia
C0036349|T048|AB|295.30|ICD9CM|Paranoid schizo-unspec|Paranoid schizo-unspec
C0036349|T048|PT|295.30|ICD9CM|Paranoid type schizophrenia, unspecified|Paranoid type schizophrenia, unspecified
C0154354|T048|AB|295.31|ICD9CM|Paranoid schizo-subchr|Paranoid schizo-subchr
C0154354|T048|PT|295.31|ICD9CM|Paranoid type schizophrenia, subchronic|Paranoid type schizophrenia, subchronic
C0270398|T048|AB|295.32|ICD9CM|Paranoid schizo-chronic|Paranoid schizo-chronic
C0270398|T048|PT|295.32|ICD9CM|Paranoid type schizophrenia, chronic|Paranoid type schizophrenia, chronic
C0154356|T048|AB|295.33|ICD9CM|Paran schizo-subchr/exac|Paran schizo-subchr/exac
C0154356|T048|PT|295.33|ICD9CM|Paranoid type schizophrenia, subchronic with acute exacerbation|Paranoid type schizophrenia, subchronic with acute exacerbation
C0154357|T048|AB|295.34|ICD9CM|Paran schizo-chr/exacerb|Paran schizo-chr/exacerb
C0154357|T048|PT|295.34|ICD9CM|Paranoid type schizophrenia, chronic with acute exacerbation|Paranoid type schizophrenia, chronic with acute exacerbation
C0154358|T048|AB|295.35|ICD9CM|Paranoid schizo-remiss|Paranoid schizo-remiss
C0154358|T048|PT|295.35|ICD9CM|Paranoid type schizophrenia, in remission|Paranoid type schizophrenia, in remission
C0036358|T048|HT|295.4|ICD9CM|Schizophreniform disorder|Schizophreniform disorder
C0813173|T048|AB|295.40|ICD9CM|Schizophreniform dis NOS|Schizophreniform dis NOS
C0813173|T048|PT|295.40|ICD9CM|Schizophreniform disorder, unspecified|Schizophreniform disorder, unspecified
C0154360|T048|AB|295.41|ICD9CM|Schizophrenic dis-subchr|Schizophrenic dis-subchr
C0154360|T048|PT|295.41|ICD9CM|Schizophreniform disorder, subchronic|Schizophreniform disorder, subchronic
C0154361|T048|AB|295.42|ICD9CM|Schizophren dis-chronic|Schizophren dis-chronic
C0154361|T048|PT|295.42|ICD9CM|Schizophreniform disorder, chronic|Schizophreniform disorder, chronic
C0154362|T048|AB|295.43|ICD9CM|Schizo dis-subchr/exacer|Schizo dis-subchr/exacer
C0154362|T048|PT|295.43|ICD9CM|Schizophreniform disorder, subchronic with acute exacerbation|Schizophreniform disorder, subchronic with acute exacerbation
C0154363|T048|AB|295.44|ICD9CM|Schizophr dis-chr/exacer|Schizophr dis-chr/exacer
C0154363|T048|PT|295.44|ICD9CM|Schizophreniform disorder, chronic with acute exacerbation|Schizophreniform disorder, chronic with acute exacerbation
C0154364|T048|AB|295.45|ICD9CM|Schizophrenic dis-remiss|Schizophrenic dis-remiss
C0154364|T048|PT|295.45|ICD9CM|Schizophreniform disorder, in remission|Schizophreniform disorder, in remission
C0023105|T048|HT|295.5|ICD9CM|Latent schizophrenia|Latent schizophrenia
C0023105|T048|AB|295.50|ICD9CM|Latent schizophren-unsp|Latent schizophren-unsp
C0023105|T048|PT|295.50|ICD9CM|Latent schizophrenia, unspecified|Latent schizophrenia, unspecified
C0338810|T048|AB|295.51|ICD9CM|Lat schizophren-subchr|Lat schizophren-subchr
C0338810|T048|PT|295.51|ICD9CM|Latent schizophrenia, subchronic|Latent schizophrenia, subchronic
C0338811|T047|AB|295.52|ICD9CM|Latent schizophren-chr|Latent schizophren-chr
C0338811|T047|PT|295.52|ICD9CM|Latent schizophrenia, chronic|Latent schizophrenia, chronic
C0338812|T048|AB|295.53|ICD9CM|Lat schizo-subchr/exacer|Lat schizo-subchr/exacer
C0338812|T048|PT|295.53|ICD9CM|Latent schizophrenia, subchronic with acute exacerbation|Latent schizophrenia, subchronic with acute exacerbation
C0338813|T048|AB|295.54|ICD9CM|Latent schizo-chr/exacer|Latent schizo-chr/exacer
C0338813|T048|PT|295.54|ICD9CM|Latent schizophrenia, chronic with acute exacerbation|Latent schizophrenia, chronic with acute exacerbation
C0154369|T048|AB|295.55|ICD9CM|Lat schizophren-remiss|Lat schizophren-remiss
C0154369|T048|PT|295.55|ICD9CM|Latent schizophrenia, in remission|Latent schizophrenia, in remission
C0036351|T048|HT|295.6|ICD9CM|Residual type schizophrenic disorders|Residual type schizophrenic disorders
C0036351|T048|AB|295.60|ICD9CM|Schizophr dis resid NOS|Schizophr dis resid NOS
C0036351|T048|PT|295.60|ICD9CM|Schizophrenic disorders, residual type, unspecified|Schizophrenic disorders, residual type, unspecified
C0270406|T048|AB|295.61|ICD9CM|Schizoph dis resid-subch|Schizoph dis resid-subch
C0270406|T048|PT|295.61|ICD9CM|Schizophrenic disorders, residual type, subchronic|Schizophrenic disorders, residual type, subchronic
C0270408|T048|AB|295.62|ICD9CM|Schizophr dis resid-chr|Schizophr dis resid-chr
C0270408|T048|PT|295.62|ICD9CM|Schizophrenic disorders, residual type, chronic|Schizophrenic disorders, residual type, chronic
C0154372|T048|AB|295.63|ICD9CM|Schizo resid subchr/exac|Schizo resid subchr/exac
C0154372|T048|PT|295.63|ICD9CM|Schizophrenic disorders, residual type, subchronic with acute exacerbation|Schizophrenic disorders, residual type, subchronic with acute exacerbation
C0154373|T048|AB|295.64|ICD9CM|Schizoph resid-chro/exac|Schizoph resid-chro/exac
C0154373|T048|PT|295.64|ICD9CM|Schizophrenic disorders, residual type, chronic with acute exacerbation|Schizophrenic disorders, residual type, chronic with acute exacerbation
C0154374|T048|AB|295.65|ICD9CM|Schizoph dis resid-remis|Schizoph dis resid-remis
C0154374|T048|PT|295.65|ICD9CM|Schizophrenic disorders, residual type, in remission|Schizophrenic disorders, residual type, in remission
C0036337|T048|HT|295.7|ICD9CM|Schizoaffective disorder|Schizoaffective disorder
C0375162|T048|AB|295.70|ICD9CM|Schizoaffective dis NOS|Schizoaffective dis NOS
C0375162|T048|PT|295.70|ICD9CM|Schizoaffective disorder, unspecified|Schizoaffective disorder, unspecified
C0154375|T048|PT|295.71|ICD9CM|Schizoaffective disorder, subchronic|Schizoaffective disorder, subchronic
C0154375|T048|AB|295.71|ICD9CM|Schizoaffectv dis-subchr|Schizoaffectv dis-subchr
C0154376|T048|AB|295.72|ICD9CM|Schizoaffective dis-chr|Schizoaffective dis-chr
C0154376|T048|PT|295.72|ICD9CM|Schizoaffective disorder, chronic|Schizoaffective disorder, chronic
C0154377|T048|AB|295.73|ICD9CM|Schizoaff dis-subch/exac|Schizoaff dis-subch/exac
C0154377|T048|PT|295.73|ICD9CM|Schizoaffective disorder, subchronic with acute exacerbation|Schizoaffective disorder, subchronic with acute exacerbation
C0154378|T048|PT|295.74|ICD9CM|Schizoaffective disorder, chronic with acute exacerbation|Schizoaffective disorder, chronic with acute exacerbation
C0154378|T048|AB|295.74|ICD9CM|Schizoafftv dis-chr/exac|Schizoafftv dis-chr/exac
C0338828|T048|PT|295.75|ICD9CM|Schizoaffective disorder, in remission|Schizoaffective disorder, in remission
C0338828|T048|AB|295.75|ICD9CM|Schizoaffectve dis-remis|Schizoaffectve dis-remis
C0029838|T048|HT|295.8|ICD9CM|Other specified types of schizophrenia|Other specified types of schizophrenia
C0029838|T048|PT|295.80|ICD9CM|Other specified types of schizophrenia, unspecified|Other specified types of schizophrenia, unspecified
C0029838|T048|AB|295.80|ICD9CM|Schizophrenia NEC-unspec|Schizophrenia NEC-unspec
C0154380|T048|PT|295.81|ICD9CM|Other specified types of schizophrenia, subchronic|Other specified types of schizophrenia, subchronic
C0154380|T048|AB|295.81|ICD9CM|Schizophrenia NEC-subchr|Schizophrenia NEC-subchr
C0154381|T048|PT|295.82|ICD9CM|Other specified types of schizophrenia, chronic|Other specified types of schizophrenia, chronic
C0154381|T048|AB|295.82|ICD9CM|Schizophrenia NEC-chr|Schizophrenia NEC-chr
C0154382|T048|PT|295.83|ICD9CM|Other specified types of schizophrenia, subchronic with acute exacerbation|Other specified types of schizophrenia, subchronic with acute exacerbation
C0154382|T048|AB|295.83|ICD9CM|Schizo NEC-subchr/exacer|Schizo NEC-subchr/exacer
C0154383|T048|PT|295.84|ICD9CM|Other specified types of schizophrenia, chronic with acute exacerbation|Other specified types of schizophrenia, chronic with acute exacerbation
C0154383|T048|AB|295.84|ICD9CM|Schizo NEC-chr/exacerb|Schizo NEC-chr/exacerb
C0154384|T048|PT|295.85|ICD9CM|Other specified types of schizophrenia, in remission|Other specified types of schizophrenia, in remission
C0154384|T048|AB|295.85|ICD9CM|Schizophrenia NEC-remiss|Schizophrenia NEC-remiss
C0036341|T048|HT|295.9|ICD9CM|Unspecified schizophrenia|Unspecified schizophrenia
C0036341|T048|AB|295.90|ICD9CM|Schizophrenia NOS-unspec|Schizophrenia NOS-unspec
C0036341|T048|PT|295.90|ICD9CM|Unspecified schizophrenia, unspecified|Unspecified schizophrenia, unspecified
C0270381|T048|AB|295.91|ICD9CM|Schizophrenia NOS-subchr|Schizophrenia NOS-subchr
C0270381|T048|PT|295.91|ICD9CM|Unspecified schizophrenia, subchronic|Unspecified schizophrenia, subchronic
C0270403|T048|AB|295.92|ICD9CM|Schizophrenia NOS-chr|Schizophrenia NOS-chr
C0270403|T048|PT|295.92|ICD9CM|Unspecified schizophrenia, chronic|Unspecified schizophrenia, chronic
C0154387|T048|AB|295.93|ICD9CM|Schizo NOS-subchr/exacer|Schizo NOS-subchr/exacer
C0154387|T048|PT|295.93|ICD9CM|Unspecified schizophrenia, subchronic with acute exacerbation|Unspecified schizophrenia, subchronic with acute exacerbation
C0154388|T048|AB|295.94|ICD9CM|Schizo NOS-chr/exacerb|Schizo NOS-chr/exacerb
C0154388|T048|PT|295.94|ICD9CM|Unspecified schizophrenia, chronic with acute exacerbation|Unspecified schizophrenia, chronic with acute exacerbation
C0270384|T048|AB|295.95|ICD9CM|Schizophrenia NOS-remiss|Schizophrenia NOS-remiss
C0270384|T048|PT|295.95|ICD9CM|Unspecified schizophrenia, in remission|Unspecified schizophrenia, in remission
C1456434|T048|HT|296|ICD9CM|Episodic mood disorders|Episodic mood disorders
C0236756|T048|HT|296.0|ICD9CM|Bipolar I disorder, single manic episode|Bipolar I disorder, single manic episode
C0236756|T048|AB|296.00|ICD9CM|Bipol I single manic NOS|Bipol I single manic NOS
C0236756|T048|PT|296.00|ICD9CM|Bipolar I disorder, single manic episode, unspecified|Bipolar I disorder, single manic episode, unspecified
C0236757|T048|AB|296.01|ICD9CM|Bipol I single manc-mild|Bipol I single manc-mild
C0236757|T048|PT|296.01|ICD9CM|Bipolar I disorder, single manic episode, mild|Bipolar I disorder, single manic episode, mild
C0236758|T048|AB|296.02|ICD9CM|Bipol I single manic-mod|Bipol I single manic-mod
C0236758|T048|PT|296.02|ICD9CM|Bipolar I disorder, single manic episode, moderate|Bipolar I disorder, single manic episode, moderate
C0154392|T048|AB|296.03|ICD9CM|Bipol I sing-sev w/o psy|Bipol I sing-sev w/o psy
C0154392|T048|PT|296.03|ICD9CM|Bipolar I disorder, single manic episode, severe, without mention of psychotic behavior|Bipolar I disorder, single manic episode, severe, without mention of psychotic behavior
C0154393|T048|AB|296.04|ICD9CM|Bipo I sin man-sev w psy|Bipo I sin man-sev w psy
C0154393|T048|PT|296.04|ICD9CM|Bipolar I disorder, single manic episode, severe, specified as with psychotic behavior|Bipolar I disorder, single manic episode, severe, specified as with psychotic behavior
C0338843|T048|AB|296.05|ICD9CM|Bipol I sing man rem NOS|Bipol I sing man rem NOS
C0338843|T048|PT|296.05|ICD9CM|Bipolar I disorder, single manic episode, in partial or unspecified remission|Bipolar I disorder, single manic episode, in partial or unspecified remission
C0236762|T048|AB|296.06|ICD9CM|Bipol I single manic rem|Bipol I single manic rem
C0236762|T048|PT|296.06|ICD9CM|Bipolar I disorder, single manic episode, in full remission|Bipolar I disorder, single manic episode, in full remission
C0338832|T048|HT|296.1|ICD9CM|Manic disorder, recurrent episode|Manic disorder, recurrent episode
C0375164|T048|PT|296.10|ICD9CM|Manic affective disorder, recurrent episode, unspecified|Manic affective disorder, recurrent episode, unspecified
C0375164|T048|AB|296.10|ICD9CM|Recur manic dis-unspec|Recur manic dis-unspec
C0154397|T048|PT|296.11|ICD9CM|Manic affective disorder, recurrent episode, mild|Manic affective disorder, recurrent episode, mild
C0154397|T048|AB|296.11|ICD9CM|Recur manic dis-mild|Recur manic dis-mild
C0154398|T048|PT|296.12|ICD9CM|Manic affective disorder, recurrent episode, moderate|Manic affective disorder, recurrent episode, moderate
C0154398|T048|AB|296.12|ICD9CM|Recur manic dis-mod|Recur manic dis-mod
C0154399|T048|PT|296.13|ICD9CM|Manic affective disorder, recurrent episode, severe, without mention of psychotic behavior|Manic affective disorder, recurrent episode, severe, without mention of psychotic behavior
C0154399|T048|AB|296.13|ICD9CM|Recur manic dis-severe|Recur manic dis-severe
C0154400|T048|PT|296.14|ICD9CM|Manic affective disorder, recurrent episode, severe, specified as with psychotic behavior|Manic affective disorder, recurrent episode, severe, specified as with psychotic behavior
C0154400|T048|AB|296.14|ICD9CM|Recur manic-sev w psycho|Recur manic-sev w psycho
C0338838|T048|PT|296.15|ICD9CM|Manic affective disorder, recurrent episode, in partial or unspecified remission|Manic affective disorder, recurrent episode, in partial or unspecified remission
C0338838|T048|AB|296.15|ICD9CM|Recur manic-part remiss|Recur manic-part remiss
C0338839|T048|PT|296.16|ICD9CM|Manic affective disorder, recurrent episode, in full remission|Manic affective disorder, recurrent episode, in full remission
C0338839|T048|AB|296.16|ICD9CM|Recur manic-full remiss|Recur manic-full remiss
C0024517|T048|HT|296.2|ICD9CM|Major depressive disorder, single episode|Major depressive disorder, single episode
C0024517|T048|AB|296.20|ICD9CM|Depress psychosis-unspec|Depress psychosis-unspec
C0024517|T048|PT|296.20|ICD9CM|Major depressive affective disorder, single episode, unspecified|Major depressive affective disorder, single episode, unspecified
C0154403|T048|AB|296.21|ICD9CM|Depress psychosis-mild|Depress psychosis-mild
C0154403|T048|PT|296.21|ICD9CM|Major depressive affective disorder, single episode, mild|Major depressive affective disorder, single episode, mild
C0154404|T048|AB|296.22|ICD9CM|Depressive psychosis-mod|Depressive psychosis-mod
C0154404|T048|PT|296.22|ICD9CM|Major depressive affective disorder, single episode, moderate|Major depressive affective disorder, single episode, moderate
C0154405|T048|AB|296.23|ICD9CM|Depress psychosis-severe|Depress psychosis-severe
C0154405|T048|PT|296.23|ICD9CM|Major depressive affective disorder, single episode, severe, without mention of psychotic behavior|Major depressive affective disorder, single episode, severe, without mention of psychotic behavior
C0154406|T048|AB|296.24|ICD9CM|Depr psychos-sev w psych|Depr psychos-sev w psych
C0154406|T048|PT|296.24|ICD9CM|Major depressive affective disorder, single episode, severe, specified as with psychotic behavior|Major depressive affective disorder, single episode, severe, specified as with psychotic behavior
C0338886|T048|AB|296.25|ICD9CM|Depr psychos-part remiss|Depr psychos-part remiss
C0338886|T048|PT|296.25|ICD9CM|Major depressive affective disorder, single episode, in partial or unspecified remission|Major depressive affective disorder, single episode, in partial or unspecified remission
C0154408|T048|AB|296.26|ICD9CM|Depr psychos-full remiss|Depr psychos-full remiss
C0154408|T048|PT|296.26|ICD9CM|Major depressive affective disorder, single episode, in full remission|Major depressive affective disorder, single episode, in full remission
C0154409|T048|HT|296.3|ICD9CM|Major depressive disorder, recurrent episode|Major depressive disorder, recurrent episode
C0154409|T048|PT|296.30|ICD9CM|Major depressive affective disorder, recurrent episode, unspecified|Major depressive affective disorder, recurrent episode, unspecified
C0154409|T048|AB|296.30|ICD9CM|Recurr depr psychos-unsp|Recurr depr psychos-unsp
C3665435|T048|PT|296.31|ICD9CM|Major depressive affective disorder, recurrent episode, mild|Major depressive affective disorder, recurrent episode, mild
C3665435|T048|AB|296.31|ICD9CM|Recurr depr psychos-mild|Recurr depr psychos-mild
C0154411|T048|PT|296.32|ICD9CM|Major depressive affective disorder, recurrent episode, moderate|Major depressive affective disorder, recurrent episode, moderate
C0154411|T048|AB|296.32|ICD9CM|Recurr depr psychos-mod|Recurr depr psychos-mod
C0154412|T048|AB|296.33|ICD9CM|Recur depr psych-severe|Recur depr psych-severe
C0154413|T048|PT|296.34|ICD9CM|Major depressive affective disorder, recurrent episode, severe, specified as with psychotic behavior|Major depressive affective disorder, recurrent episode, severe, specified as with psychotic behavior
C0154413|T048|AB|296.34|ICD9CM|Rec depr psych-psychotic|Rec depr psych-psychotic
C0338893|T048|PT|296.35|ICD9CM|Major depressive affective disorder, recurrent episode, in partial or unspecified remission|Major depressive affective disorder, recurrent episode, in partial or unspecified remission
C0338893|T048|AB|296.35|ICD9CM|Recur depr psyc-part rem|Recur depr psyc-part rem
C3665667|T048|PT|296.36|ICD9CM|Major depressive affective disorder, recurrent episode, in full remission|Major depressive affective disorder, recurrent episode, in full remission
C3665667|T048|AB|296.36|ICD9CM|Recur depr psyc-full rem|Recur depr psyc-full rem
C1456304|T048|HT|296.4|ICD9CM|Bipolar I disorder, most recent episode (or current) manic|Bipolar I disorder, most recent episode (or current) manic
C0024713|T048|AB|296.40|ICD9CM|Bipol I currnt manic NOS|Bipol I currnt manic NOS
C0024713|T048|PT|296.40|ICD9CM|Bipolar I disorder, most recent episode (or current) manic, unspecified|Bipolar I disorder, most recent episode (or current) manic, unspecified
C0154417|T048|AB|296.41|ICD9CM|Bipol I curnt manic-mild|Bipol I curnt manic-mild
C0154417|T048|PT|296.41|ICD9CM|Bipolar I disorder, most recent episode (or current) manic, mild|Bipolar I disorder, most recent episode (or current) manic, mild
C0154418|T048|AB|296.42|ICD9CM|Bipol I currnt manic-mod|Bipol I currnt manic-mod
C0154418|T048|PT|296.42|ICD9CM|Bipolar I disorder, most recent episode (or current) manic, moderate|Bipolar I disorder, most recent episode (or current) manic, moderate
C0154419|T048|AB|296.43|ICD9CM|Bipol I manc-sev w/o psy|Bipol I manc-sev w/o psy
C0154420|T048|AB|296.44|ICD9CM|Bipol I manic-sev w psy|Bipol I manic-sev w psy
C0154421|T048|AB|296.45|ICD9CM|Bipol I cur man part rem|Bipol I cur man part rem
C0154421|T048|PT|296.45|ICD9CM|Bipolar I disorder, most recent episode (or current) manic, in partial or unspecified remission|Bipolar I disorder, most recent episode (or current) manic, in partial or unspecified remission
C0154422|T048|AB|296.46|ICD9CM|Bipol I cur man full rem|Bipol I cur man full rem
C0154422|T048|PT|296.46|ICD9CM|Bipolar I disorder, most recent episode (or current) manic, in full remission|Bipolar I disorder, most recent episode (or current) manic, in full remission
C1456305|T048|HT|296.5|ICD9CM|Bipolar I disorder, most recent episode (or current) depressed|Bipolar I disorder, most recent episode (or current) depressed
C0236773|T048|AB|296.50|ICD9CM|Bipol I cur depres NOS|Bipol I cur depres NOS
C0236773|T048|PT|296.50|ICD9CM|Bipolar I disorder, most recent episode (or current) depressed, unspecified|Bipolar I disorder, most recent episode (or current) depressed, unspecified
C0154424|T048|AB|296.51|ICD9CM|Bipol I cur depress-mild|Bipol I cur depress-mild
C0154424|T048|PT|296.51|ICD9CM|Bipolar I disorder, most recent episode (or current) depressed, mild|Bipolar I disorder, most recent episode (or current) depressed, mild
C0154425|T048|AB|296.52|ICD9CM|Bipol I cur depress-mod|Bipol I cur depress-mod
C0154425|T048|PT|296.52|ICD9CM|Bipolar I disorder, most recent episode (or current) depressed, moderate|Bipolar I disorder, most recent episode (or current) depressed, moderate
C0154426|T048|AB|296.53|ICD9CM|Bipol I curr dep w/o psy|Bipol I curr dep w/o psy
C0154427|T048|AB|296.54|ICD9CM|Bipol I currnt dep w psy|Bipol I currnt dep w psy
C0154428|T048|AB|296.55|ICD9CM|Bipol I cur dep rem NOS|Bipol I cur dep rem NOS
C0154428|T048|PT|296.55|ICD9CM|Bipolar I disorder, most recent episode (or current) depressed, in partial or unspecified remission|Bipolar I disorder, most recent episode (or current) depressed, in partial or unspecified remission
C0154429|T048|AB|296.56|ICD9CM|Bipol I currnt dep remis|Bipol I currnt dep remis
C0154429|T048|PT|296.56|ICD9CM|Bipolar I disorder, most recent episode (or current) depressed, in full remission|Bipolar I disorder, most recent episode (or current) depressed, in full remission
C1456306|T048|HT|296.6|ICD9CM|Bipolar I disorder, most recent episode (or current) mixed|Bipolar I disorder, most recent episode (or current) mixed
C0236780|T048|AB|296.60|ICD9CM|Bipol I currnt mixed NOS|Bipol I currnt mixed NOS
C0236780|T048|PT|296.60|ICD9CM|Bipolar I disorder, most recent episode (or current) mixed, unspecified|Bipolar I disorder, most recent episode (or current) mixed, unspecified
C2874891|T048|AB|296.61|ICD9CM|Bipol I currnt mix-mild|Bipol I currnt mix-mild
C2874891|T048|PT|296.61|ICD9CM|Bipolar I disorder, most recent episode (or current) mixed, mild|Bipolar I disorder, most recent episode (or current) mixed, mild
C2874892|T048|AB|296.62|ICD9CM|Bipol I currnt mixed-mod|Bipol I currnt mixed-mod
C2874892|T048|PT|296.62|ICD9CM|Bipolar I disorder, most recent episode (or current) mixed, moderate|Bipolar I disorder, most recent episode (or current) mixed, moderate
C0154432|T048|AB|296.63|ICD9CM|Bipol I cur mix w/o psy|Bipol I cur mix w/o psy
C0154433|T048|AB|296.64|ICD9CM|Bipol I cur mixed w psy|Bipol I cur mixed w psy
C0154434|T048|AB|296.65|ICD9CM|Bipol I cur mix-part rem|Bipol I cur mix-part rem
C0154434|T048|PT|296.65|ICD9CM|Bipolar I disorder, most recent episode (or current) mixed, in partial or unspecified remission|Bipolar I disorder, most recent episode (or current) mixed, in partial or unspecified remission
C0270434|T048|AB|296.66|ICD9CM|Bipol I cur mixed remiss|Bipol I cur mixed remiss
C0270434|T048|PT|296.66|ICD9CM|Bipolar I disorder, most recent episode (or current) mixed, in full remission|Bipolar I disorder, most recent episode (or current) mixed, in full remission
C1456307|T048|PT|296.7|ICD9CM|Bipolar I disorder, most recent episode (or current) unspecified|Bipolar I disorder, most recent episode (or current) unspecified
C1456307|T048|AB|296.7|ICD9CM|Bipolor I current NOS|Bipolor I current NOS
C1456309|T048|HT|296.8|ICD9CM|Other and unspecified bipolar disorders|Other and unspecified bipolar disorders
C0005586|T048|AB|296.80|ICD9CM|Bipolar disorder NOS|Bipolar disorder NOS
C0005586|T048|PT|296.80|ICD9CM|Bipolar disorder, unspecified|Bipolar disorder, unspecified
C0154436|T048|AB|296.81|ICD9CM|Atypical manic disorder|Atypical manic disorder
C0154436|T048|PT|296.81|ICD9CM|Atypical manic disorder|Atypical manic disorder
C0154437|T048|AB|296.82|ICD9CM|Atypical depressive dis|Atypical depressive dis
C0154437|T048|PT|296.82|ICD9CM|Atypical depressive disorder|Atypical depressive disorder
C1456308|T048|AB|296.89|ICD9CM|Bipolar disorder NEC|Bipolar disorder NEC
C1456308|T048|PT|296.89|ICD9CM|Other bipolar disorders|Other bipolar disorders
C1456311|T048|HT|296.9|ICD9CM|Other and unspecified episodic mood disorder|Other and unspecified episodic mood disorder
C1456434|T048|AB|296.90|ICD9CM|Episodic mood disord NOS|Episodic mood disord NOS
C1456434|T048|PT|296.90|ICD9CM|Unspecified episodic mood disorder|Unspecified episodic mood disorder
C1456310|T048|AB|296.99|ICD9CM|Episodic mood disord NEC|Episodic mood disord NEC
C1456310|T048|PT|296.99|ICD9CM|Other specified episodic mood disorder|Other specified episodic mood disorder
C1456783|T048|HT|297|ICD9CM|Paranoid states (Delusional disorders)|Paranoid states (Delusional disorders)
C0154440|T048|AB|297.0|ICD9CM|Paranoid state, simple|Paranoid state, simple
C0154440|T048|PT|297.0|ICD9CM|Paranoid state, simple|Paranoid state, simple
C0011251|T048|AB|297.1|ICD9CM|Delusional disorder|Delusional disorder
C0011251|T048|PT|297.1|ICD9CM|Delusional disorder|Delusional disorder
C0030484|T048|AB|297.2|ICD9CM|Paraphrenia|Paraphrenia
C0030484|T048|PT|297.2|ICD9CM|Paraphrenia|Paraphrenia
C0036939|T048|AB|297.3|ICD9CM|Shared psychotic disord|Shared psychotic disord
C0036939|T048|PT|297.3|ICD9CM|Shared psychotic disorder|Shared psychotic disorder
C0154441|T048|PT|297.8|ICD9CM|Other specified paranoid states|Other specified paranoid states
C0154441|T048|AB|297.8|ICD9CM|Paranoid states NEC|Paranoid states NEC
C1456786|T048|AB|297.9|ICD9CM|Paranoid state NOS|Paranoid state NOS
C1456786|T048|PT|297.9|ICD9CM|Unspecified paranoid state|Unspecified paranoid state
C0154442|T048|HT|298|ICD9CM|Other nonorganic psychoses|Other nonorganic psychoses
C3665340|T048|PT|298.0|ICD9CM|Depressive type psychosis|Depressive type psychosis
C3665340|T048|AB|298.0|ICD9CM|React depress psychosis|React depress psychosis
C0338930|T048|AB|298.1|ICD9CM|Excitativ type psychosis|Excitativ type psychosis
C0338930|T048|PT|298.1|ICD9CM|Excitative type psychosis|Excitative type psychosis
C0152124|T048|AB|298.2|ICD9CM|Reactive confusion|Reactive confusion
C0152124|T048|PT|298.2|ICD9CM|Reactive confusion|Reactive confusion
C0152125|T048|AB|298.3|ICD9CM|Acute paranoid reaction|Acute paranoid reaction
C0152125|T048|PT|298.3|ICD9CM|Acute paranoid reaction|Acute paranoid reaction
C0152126|T048|AB|298.4|ICD9CM|Psychogen paranoid psych|Psychogen paranoid psych
C0152126|T048|PT|298.4|ICD9CM|Psychogenic paranoid psychosis|Psychogenic paranoid psychosis
C0029516|T048|PT|298.8|ICD9CM|Other and unspecified reactive psychosis|Other and unspecified reactive psychosis
C0029516|T048|AB|298.8|ICD9CM|React psychosis NEC/NOS|React psychosis NEC/NOS
C0033975|T048|AB|298.9|ICD9CM|Psychosis NOS|Psychosis NOS
C0033975|T048|PT|298.9|ICD9CM|Unspecified psychosis|Unspecified psychosis
C0524528|T048|HT|299|ICD9CM|Pervasive developmental disorders|Pervasive developmental disorders
C0004352|T048|HT|299.0|ICD9CM|Autistic disorder|Autistic disorder
C0154446|T048|AB|299.00|ICD9CM|Autistic disord-current|Autistic disord-current
C0154446|T048|PT|299.00|ICD9CM|Autistic disorder, current or active state|Autistic disorder, current or active state
C0338984|T048|AB|299.01|ICD9CM|Autistic disord-residual|Autistic disord-residual
C0338984|T048|PT|299.01|ICD9CM|Autistic disorder, residual state|Autistic disorder, residual state
C0236791|T048|HT|299.1|ICD9CM|Childhood disintegrative disorder|Childhood disintegrative disorder
C0154448|T048|AB|299.10|ICD9CM|Childhd disintegr-active|Childhd disintegr-active
C0154448|T048|PT|299.10|ICD9CM|Childhood disintegrative disorder, current or active state|Childhood disintegrative disorder, current or active state
C0154449|T048|AB|299.11|ICD9CM|Childhd disintegr-resid|Childhd disintegr-resid
C0154449|T048|PT|299.11|ICD9CM|Childhood disintegrative disorder, residual state|Childhood disintegrative disorder, residual state
C1456313|T048|HT|299.8|ICD9CM|Other specified pervasive developmental disorders|Other specified pervasive developmental disorders
C0154451|T048|PT|299.80|ICD9CM|Other specified pervasive developmental disorders, current or active state|Other specified pervasive developmental disorders, current or active state
C0154451|T048|AB|299.80|ICD9CM|Pervasv dev dis-cur NEC|Pervasv dev dis-cur NEC
C0154452|T048|PT|299.81|ICD9CM|Other specified pervasive developmental disorders, residual state|Other specified pervasive developmental disorders, residual state
C0154452|T048|AB|299.81|ICD9CM|Pervasv dev dis-res NEC|Pervasv dev dis-res NEC
C0524528|T048|HT|299.9|ICD9CM|Unspecified pervasive developmental disorder|Unspecified pervasive developmental disorder
C0154453|T048|AB|299.90|ICD9CM|Pervasv dev dis-cur NOS|Pervasv dev dis-cur NOS
C0154453|T048|PT|299.90|ICD9CM|Unspecified pervasive developmental disorder, current or active state|Unspecified pervasive developmental disorder, current or active state
C0154454|T048|AB|299.91|ICD9CM|Pervasv dev dis-res NOS|Pervasv dev dis-res NOS
C0154454|T048|PT|299.91|ICD9CM|Unspecified pervasive developmental disorder, residual state|Unspecified pervasive developmental disorder, residual state
C1456316|T048|HT|300|ICD9CM|Anxiety, dissociative and somatoform disorders|Anxiety, dissociative and somatoform disorders
C0338608|T048|HT|300-316.99|ICD9CM|NEUROTIC DISORDERS, PERSONALITY DISORDERS, AND OTHER NONPSYCHOTIC MENTAL DISORDERS|NEUROTIC DISORDERS, PERSONALITY DISORDERS, AND OTHER NONPSYCHOTIC MENTAL DISORDERS
C0700613|T048|HT|300.0|ICD9CM|Anxiety states|Anxiety states
C0700613|T048|AB|300.00|ICD9CM|Anxiety state NOS|Anxiety state NOS
C0700613|T048|PT|300.00|ICD9CM|Anxiety state, unspecified|Anxiety state, unspecified
C0236794|T048|AB|300.01|ICD9CM|Panic dis w/o agorphobia|Panic dis w/o agorphobia
C0236794|T048|PT|300.01|ICD9CM|Panic disorder without agoraphobia|Panic disorder without agoraphobia
C0270549|T048|AB|300.02|ICD9CM|Generalized anxiety dis|Generalized anxiety dis
C0270549|T048|PT|300.02|ICD9CM|Generalized anxiety disorder|Generalized anxiety disorder
C0154455|T048|AB|300.09|ICD9CM|Anxiety state NEC|Anxiety state NEC
C0154455|T048|PT|300.09|ICD9CM|Other anxiety states|Other anxiety states
C1456314|T048|HT|300.1|ICD9CM|Dissociative, conversion and factitious disorders|Dissociative, conversion and factitious disorders
C0020701|T048|AB|300.10|ICD9CM|Hysteria NOS|Hysteria NOS
C0020701|T048|PT|300.10|ICD9CM|Hysteria, unspecified|Hysteria, unspecified
C0009946|T048|AB|300.11|ICD9CM|Conversion disorder|Conversion disorder
C0009946|T048|PT|300.11|ICD9CM|Conversion disorder|Conversion disorder
C0236795|T048|AB|300.12|ICD9CM|Dissociative amnesia|Dissociative amnesia
C0236795|T048|PT|300.12|ICD9CM|Dissociative amnesia|Dissociative amnesia
C0020703|T048|AB|300.13|ICD9CM|Dissociative fugue|Dissociative fugue
C0020703|T048|PT|300.13|ICD9CM|Dissociative fugue|Dissociative fugue
C0026773|T048|PT|300.14|ICD9CM|Dissociative identity disorder|Dissociative identity disorder
C0026773|T048|AB|300.14|ICD9CM|Dissociatve identity dis|Dissociatve identity dis
C0012746|T048|PT|300.15|ICD9CM|Dissociative disorder or reaction, unspecified|Dissociative disorder or reaction, unspecified
C0012746|T048|AB|300.15|ICD9CM|Dissociative react NOS|Dissociative react NOS
C0015481|T048|AB|300.16|ICD9CM|Factitious dis w symptom|Factitious dis w symptom
C0015481|T048|PT|300.16|ICD9CM|Factitious disorder with predominantly psychological signs and symptoms|Factitious disorder with predominantly psychological signs and symptoms
C0154456|T048|AB|300.19|ICD9CM|Factitious ill NEC/NOS|Factitious ill NEC/NOS
C0154456|T048|PT|300.19|ICD9CM|Other and unspecified factitious illness|Other and unspecified factitious illness
C0349231|T048|HT|300.2|ICD9CM|Phobic disorders|Phobic disorders
C0349231|T048|AB|300.20|ICD9CM|Phobia NOS|Phobia NOS
C0349231|T048|PT|300.20|ICD9CM|Phobia, unspecified|Phobia, unspecified
C0236800|T048|AB|300.21|ICD9CM|Agoraphobia w panic dis|Agoraphobia w panic dis
C0236800|T048|PT|300.21|ICD9CM|Agoraphobia with panic disorder|Agoraphobia with panic disorder
C0001819|T048|AB|300.22|ICD9CM|Agoraphobia w/o panic|Agoraphobia w/o panic
C0001819|T048|PT|300.22|ICD9CM|Agoraphobia without mention of panic attacks|Agoraphobia without mention of panic attacks
C0031572|T048|AB|300.23|ICD9CM|Social phobia|Social phobia
C0031572|T048|PT|300.23|ICD9CM|Social phobia|Social phobia
C1456315|T048|AB|300.29|ICD9CM|Isolated/spec phobia NEC|Isolated/spec phobia NEC
C1456315|T048|PT|300.29|ICD9CM|Other isolated or specific phobias|Other isolated or specific phobias
C0028768|T048|AB|300.3|ICD9CM|Obsessive-compulsive dis|Obsessive-compulsive dis
C0028768|T048|PT|300.3|ICD9CM|Obsessive-compulsive disorders|Obsessive-compulsive disorders
C0013415|T048|AB|300.4|ICD9CM|Dysthymic disorder|Dysthymic disorder
C0013415|T048|PT|300.4|ICD9CM|Dysthymic disorder|Dysthymic disorder
C0027804|T048|AB|300.5|ICD9CM|Neurasthenia|Neurasthenia
C0027804|T048|PT|300.5|ICD9CM|Neurasthenia|Neurasthenia
C0683416|T048|AB|300.6|ICD9CM|Depersonalization disord|Depersonalization disord
C0683416|T048|PT|300.6|ICD9CM|Depersonalization disorder|Depersonalization disorder
C0020604|T048|AB|300.7|ICD9CM|Hypochondriasis|Hypochondriasis
C0020604|T048|PT|300.7|ICD9CM|Hypochondriasis|Hypochondriasis
C0037650|T048|HT|300.8|ICD9CM|Somatoform disorders|Somatoform disorders
C0520482|T048|AB|300.81|ICD9CM|Somatization disorder|Somatization disorder
C0520482|T048|PT|300.81|ICD9CM|Somatization disorder|Somatization disorder
C0041672|T048|AB|300.82|ICD9CM|Undiff somatoform disrdr|Undiff somatoform disrdr
C0041672|T048|PT|300.82|ICD9CM|Undifferentiated somatoform disorder|Undifferentiated somatoform disorder
C0349249|T048|PT|300.89|ICD9CM|Other somatoform disorders|Other somatoform disorders
C0349249|T048|AB|300.89|ICD9CM|Somatoform disorders NEC|Somatoform disorders NEC
C0041857|T048|AB|300.9|ICD9CM|Nonpsychotic disord NOS|Nonpsychotic disord NOS
C0041857|T048|PT|300.9|ICD9CM|Unspecified nonpsychotic mental disorder|Unspecified nonpsychotic mental disorder
C0031212|T048|HT|301|ICD9CM|Personality disorders|Personality disorders
C0030477|T048|AB|301.0|ICD9CM|Paranoid personality|Paranoid personality
C0030477|T048|PT|301.0|ICD9CM|Paranoid personality disorder|Paranoid personality disorder
C0010598|T048|HT|301.1|ICD9CM|Affective personality disorder|Affective personality disorder
C0010598|T048|AB|301.10|ICD9CM|Affectiv personality NOS|Affectiv personality NOS
C0010598|T048|PT|301.10|ICD9CM|Affective personality disorder, unspecified|Affective personality disorder, unspecified
C0154459|T048|AB|301.11|ICD9CM|Chronic hypomanic person|Chronic hypomanic person
C0154459|T048|PT|301.11|ICD9CM|Chronic hypomanic personality disorder|Chronic hypomanic personality disorder
C3665457|T048|AB|301.12|ICD9CM|Chr depressive person|Chr depressive person
C3665457|T048|PT|301.12|ICD9CM|Chronic depressive personality disorder|Chronic depressive personality disorder
C0010598|T048|AB|301.13|ICD9CM|Cyclothymic disorder|Cyclothymic disorder
C0010598|T048|PT|301.13|ICD9CM|Cyclothymic disorder|Cyclothymic disorder
C0036339|T048|HT|301.2|ICD9CM|Schizoid personality disorder|Schizoid personality disorder
C0036339|T048|PT|301.20|ICD9CM|Schizoid personality disorder, unspecified|Schizoid personality disorder, unspecified
C0036339|T048|AB|301.20|ICD9CM|Schizoid personality NOS|Schizoid personality NOS
C0338969|T048|AB|301.21|ICD9CM|Introverted personality|Introverted personality
C0338969|T048|PT|301.21|ICD9CM|Introverted personality|Introverted personality
C0036363|T048|AB|301.22|ICD9CM|Schizotypal person dis|Schizotypal person dis
C0036363|T048|PT|301.22|ICD9CM|Schizotypal personality disorder|Schizotypal personality disorder
C0152183|T048|AB|301.3|ICD9CM|Explosive personality|Explosive personality
C0152183|T048|PT|301.3|ICD9CM|Explosive personality disorder|Explosive personality disorder
C0009595|T048|AB|301.4|ICD9CM|Obsessive-compulsive dis|Obsessive-compulsive dis
C0009595|T048|PT|301.4|ICD9CM|Obsessive-compulsive personality disorder|Obsessive-compulsive personality disorder
C0019681|T048|HT|301.5|ICD9CM|Histrionic personality disorder|Histrionic personality disorder
C0019681|T048|AB|301.50|ICD9CM|Histrionic person NOS|Histrionic person NOS
C0019681|T048|PT|301.50|ICD9CM|Histrionic personality disorder, unspecified|Histrionic personality disorder, unspecified
C0008682|T048|AB|301.51|ICD9CM|Chr factitious illness|Chr factitious illness
C0008682|T048|PT|301.51|ICD9CM|Chronic factitious illness with physical symptoms|Chronic factitious illness with physical symptoms
C0029633|T048|AB|301.59|ICD9CM|Histrionic person NEC|Histrionic person NEC
C0029633|T048|PT|301.59|ICD9CM|Other histrionic personality disorder|Other histrionic personality disorder
C0011548|T048|AB|301.6|ICD9CM|Dependent personality|Dependent personality
C0011548|T048|PT|301.6|ICD9CM|Dependent personality disorder|Dependent personality disorder
C0003431|T048|AB|301.7|ICD9CM|Antisocial personality|Antisocial personality
C0003431|T048|PT|301.7|ICD9CM|Antisocial personality disorder|Antisocial personality disorder
C0029707|T048|HT|301.8|ICD9CM|Other personality disorders|Other personality disorders
C0027402|T048|AB|301.81|ICD9CM|Narcissistic personality|Narcissistic personality
C0027402|T048|PT|301.81|ICD9CM|Narcissistic personality disorder|Narcissistic personality disorder
C0004444|T048|AB|301.82|ICD9CM|Avoidant personality dis|Avoidant personality dis
C0004444|T048|PT|301.82|ICD9CM|Avoidant personality disorder|Avoidant personality disorder
C0006012|T048|AB|301.83|ICD9CM|Borderline personality|Borderline personality
C0006012|T048|PT|301.83|ICD9CM|Borderline personality disorder|Borderline personality disorder
C0030631|T048|AB|301.84|ICD9CM|Passive-aggressiv person|Passive-aggressiv person
C0030631|T048|PT|301.84|ICD9CM|Passive-aggressive personality|Passive-aggressive personality
C0029707|T048|PT|301.89|ICD9CM|Other personality disorders|Other personality disorders
C0029707|T048|AB|301.89|ICD9CM|Personality disorder NEC|Personality disorder NEC
C0031212|T048|AB|301.9|ICD9CM|Personality disorder NOS|Personality disorder NOS
C0031212|T048|PT|301.9|ICD9CM|Unspecified personality disorder|Unspecified personality disorder
C0236989|T048|HT|302|ICD9CM|Sexual and gender identity disorders|Sexual and gender identity disorders
C0233880|T048|AB|302.0|ICD9CM|Ego-dystonic sex orient|Ego-dystonic sex orient
C0233880|T048|PT|302.0|ICD9CM|Ego-dystonic sexual orientation|Ego-dystonic sexual orientation
C0152186|T048|AB|302.1|ICD9CM|Zoophilia|Zoophilia
C0152186|T048|PT|302.1|ICD9CM|Zoophilia|Zoophilia
C0030764|T048|AB|302.2|ICD9CM|Pedophilia|Pedophilia
C0030764|T048|PT|302.2|ICD9CM|Pedophilia|Pedophilia
C0015269|T048|AB|302.4|ICD9CM|Exhibitionism|Exhibitionism
C0015269|T048|PT|302.4|ICD9CM|Exhibitionism|Exhibitionism
C0236802|T048|PT|302.6|ICD9CM|Gender identity disorder in children|Gender identity disorder in children
C0236802|T048|AB|302.6|ICD9CM|Gendr identity dis-child|Gendr identity dis-child
C3714744|T048|HT|302.7|ICD9CM|Psychosexual dysfunction|Psychosexual dysfunction
C3714744|T048|AB|302.70|ICD9CM|Psychosexual dysfunc NOS|Psychosexual dysfunc NOS
C3714744|T048|PT|302.70|ICD9CM|Psychosexual dysfunction, unspecified|Psychosexual dysfunction, unspecified
C0020594|T048|AB|302.71|ICD9CM|Hypoactive sex desire|Hypoactive sex desire
C0020594|T048|PT|302.71|ICD9CM|Hypoactive sexual desire disorder|Hypoactive sexual desire disorder
C0033950|T048|AB|302.72|ICD9CM|Inhibited sex excitement|Inhibited sex excitement
C0033950|T048|PT|302.72|ICD9CM|Psychosexual dysfunction with inhibited sexual excitement|Psychosexual dysfunction with inhibited sexual excitement
C0033948|T048|AB|302.73|ICD9CM|Female orgasmic disorder|Female orgasmic disorder
C0033948|T048|PT|302.73|ICD9CM|Female orgasmic disorder|Female orgasmic disorder
C1456319|T048|AB|302.74|ICD9CM|Male orgasmic disorder|Male orgasmic disorder
C1456319|T048|PT|302.74|ICD9CM|Male orgasmic disorder|Male orgasmic disorder
C0033038|T048|AB|302.75|ICD9CM|Premature ejaculation|Premature ejaculation
C0033038|T048|PT|302.75|ICD9CM|Premature ejaculation|Premature ejaculation
C0154466|T048|PT|302.76|ICD9CM|Dyspareunia, psychogenic|Dyspareunia, psychogenic
C0154466|T048|AB|302.76|ICD9CM|Dyspareunia,psychogenic|Dyspareunia,psychogenic
C0033951|T048|AB|302.79|ICD9CM|Psychosexual dysfunc NEC|Psychosexual dysfunc NEC
C0033951|T048|PT|302.79|ICD9CM|Psychosexual dysfunction with other specified psychosexual dysfunctions|Psychosexual dysfunction with other specified psychosexual dysfunctions
C0029825|T048|HT|302.8|ICD9CM|Other specified psychosexual disorders|Other specified psychosexual disorders
C0015957|T048|AB|302.81|ICD9CM|Fetishism|Fetishism
C0015957|T048|PT|302.81|ICD9CM|Fetishism|Fetishism
C0042979|T048|AB|302.82|ICD9CM|Voyeurism|Voyeurism
C0042979|T048|PT|302.82|ICD9CM|Voyeurism|Voyeurism
C0036908|T048|AB|302.83|ICD9CM|Sexual masochism|Sexual masochism
C0036908|T048|PT|302.83|ICD9CM|Sexual masochism|Sexual masochism
C0036913|T048|AB|302.84|ICD9CM|Sexual sadism|Sexual sadism
C0036913|T048|PT|302.84|ICD9CM|Sexual sadism|Sexual sadism
C0154467|T048|AB|302.85|ICD9CM|Gend iden dis,adol/adult|Gend iden dis,adol/adult
C0154467|T048|PT|302.85|ICD9CM|Gender identity disorder in adolescents or adults|Gender identity disorder in adolescents or adults
C0029825|T048|PT|302.89|ICD9CM|Other specified psychosexual disorders|Other specified psychosexual disorders
C0029825|T048|AB|302.89|ICD9CM|Psychosexual dis NEC|Psychosexual dis NEC
C0033953|T048|AB|302.9|ICD9CM|Psychosexual dis NOS|Psychosexual dis NOS
C0033953|T048|PT|302.9|ICD9CM|Unspecified psychosexual disorder|Unspecified psychosexual disorder
C0001973|T048|HT|303|ICD9CM|Alcohol dependence syndrome|Alcohol dependence syndrome
C0394996|T048|HT|303.0|ICD9CM|Acute alcoholic intoxication|Acute alcoholic intoxication
C0812429|T048|AB|303.00|ICD9CM|Ac alcohol intox-unspec|Ac alcohol intox-unspec
C0812429|T048|PT|303.00|ICD9CM|Acute alcoholic intoxication in alcoholism, unspecified|Acute alcoholic intoxication in alcoholism, unspecified
C0338787|T048|AB|303.01|ICD9CM|Ac alcohol intox-contin|Ac alcohol intox-contin
C0338787|T048|PT|303.01|ICD9CM|Acute alcoholic intoxication in alcoholism, continuous|Acute alcoholic intoxication in alcoholism, continuous
C0338788|T048|AB|303.02|ICD9CM|Ac alcohol intox-episod|Ac alcohol intox-episod
C0338788|T048|PT|303.02|ICD9CM|Acute alcoholic intoxication in alcoholism, episodic|Acute alcoholic intoxication in alcoholism, episodic
C0154473|T048|AB|303.03|ICD9CM|Ac alcohol intox-remiss|Ac alcohol intox-remiss
C0154473|T048|PT|303.03|ICD9CM|Acute alcoholic intoxication in alcoholism, in remission|Acute alcoholic intoxication in alcoholism, in remission
C0154474|T048|HT|303.9|ICD9CM|Other and unspecified alcohol dependence|Other and unspecified alcohol dependence
C0154474|T048|AB|303.90|ICD9CM|Alcoh dep NEC/NOS-unspec|Alcoh dep NEC/NOS-unspec
C0154474|T048|PT|303.90|ICD9CM|Other and unspecified alcohol dependence, unspecified|Other and unspecified alcohol dependence, unspecified
C0154475|T048|AB|303.91|ICD9CM|Alcoh dep NEC/NOS-contin|Alcoh dep NEC/NOS-contin
C0154475|T048|PT|303.91|ICD9CM|Other and unspecified alcohol dependence, continuous|Other and unspecified alcohol dependence, continuous
C0154476|T048|AB|303.92|ICD9CM|Alcoh dep NEC/NOS-episod|Alcoh dep NEC/NOS-episod
C0154476|T048|PT|303.92|ICD9CM|Other and unspecified alcohol dependence, episodic|Other and unspecified alcohol dependence, episodic
C0154477|T048|AB|303.93|ICD9CM|Alcoh dep NEC/NOS-remiss|Alcoh dep NEC/NOS-remiss
C0154477|T048|PT|303.93|ICD9CM|Other and unspecified alcohol dependence, in remission|Other and unspecified alcohol dependence, in remission
C1510472|T048|HT|304|ICD9CM|Drug dependence|Drug dependence
C0524662|T048|HT|304.0|ICD9CM|Opioid type dependence|Opioid type dependence
C0524662|T048|AB|304.00|ICD9CM|Opioid dependence-unspec|Opioid dependence-unspec
C0524662|T048|PT|304.00|ICD9CM|Opioid type dependence, unspecified|Opioid type dependence, unspecified
C0154478|T048|AB|304.01|ICD9CM|Opioid dependence-contin|Opioid dependence-contin
C0154478|T048|PT|304.01|ICD9CM|Opioid type dependence, continuous|Opioid type dependence, continuous
C0154479|T048|AB|304.02|ICD9CM|Opioid dependence-episod|Opioid dependence-episod
C0154479|T048|PT|304.02|ICD9CM|Opioid type dependence, episodic|Opioid type dependence, episodic
C0154480|T048|AB|304.03|ICD9CM|Opioid dependence-remiss|Opioid dependence-remiss
C0154480|T048|PT|304.03|ICD9CM|Opioid type dependence, in remission|Opioid type dependence, in remission
C0036552|T048|HT|304.1|ICD9CM|Sedative, hypnotic or anxiolytic dependence|Sedative, hypnotic or anxiolytic dependence
C0375172|T048|AB|304.10|ICD9CM|Sed,hyp,anxiolyt dep-NOS|Sed,hyp,anxiolyt dep-NOS
C0375172|T048|PT|304.10|ICD9CM|Sedative, hypnotic or anxiolytic dependence, unspecified|Sedative, hypnotic or anxiolytic dependence, unspecified
C0154482|T048|AB|304.11|ICD9CM|Sed,hyp,anxiolyt dep-con|Sed,hyp,anxiolyt dep-con
C0154482|T048|PT|304.11|ICD9CM|Sedative, hypnotic or anxiolytic dependence, continuous|Sedative, hypnotic or anxiolytic dependence, continuous
C0154483|T048|AB|304.12|ICD9CM|Sed,hyp,anxiolyt dep-epi|Sed,hyp,anxiolyt dep-epi
C0154483|T048|PT|304.12|ICD9CM|Sedative, hypnotic or anxiolytic dependence, episodic|Sedative, hypnotic or anxiolytic dependence, episodic
C2874528|T048|AB|304.13|ICD9CM|Sed,hyp,anxiolyt dep-rem|Sed,hyp,anxiolyt dep-rem
C2874528|T048|PT|304.13|ICD9CM|Sedative, hypnotic or anxiolytic dependence, in remission|Sedative, hypnotic or anxiolytic dependence, in remission
C0600427|T048|HT|304.2|ICD9CM|Cocaine dependence|Cocaine dependence
C0600427|T048|AB|304.20|ICD9CM|Cocaine depend-unspec|Cocaine depend-unspec
C0600427|T048|PT|304.20|ICD9CM|Cocaine dependence, unspecified|Cocaine dependence, unspecified
C0338762|T048|AB|304.21|ICD9CM|Cocaine depend-contin|Cocaine depend-contin
C0338762|T048|PT|304.21|ICD9CM|Cocaine dependence, continuous|Cocaine dependence, continuous
C0338763|T048|AB|304.22|ICD9CM|Cocaine depend-episodic|Cocaine depend-episodic
C0338763|T048|PT|304.22|ICD9CM|Cocaine dependence, episodic|Cocaine dependence, episodic
C0154487|T048|AB|304.23|ICD9CM|Cocaine depend-remiss|Cocaine depend-remiss
C0154487|T048|PT|304.23|ICD9CM|Cocaine dependence, in remission|Cocaine dependence, in remission
C0006870|T048|HT|304.3|ICD9CM|Cannabis dependence|Cannabis dependence
C0375174|T048|AB|304.30|ICD9CM|Cannabis depend-unspec|Cannabis depend-unspec
C0375174|T048|PT|304.30|ICD9CM|Cannabis dependence, unspecified|Cannabis dependence, unspecified
C0338757|T048|AB|304.31|ICD9CM|Cannabis depend-contin|Cannabis depend-contin
C0338757|T048|PT|304.31|ICD9CM|Cannabis dependence, continuous|Cannabis dependence, continuous
C0338758|T048|AB|304.32|ICD9CM|Cannabis depend-episodic|Cannabis depend-episodic
C0338758|T048|PT|304.32|ICD9CM|Cannabis dependence, episodic|Cannabis dependence, episodic
C0154490|T047|AB|304.33|ICD9CM|Cannabis depend-remiss|Cannabis depend-remiss
C0154490|T047|PT|304.33|ICD9CM|Cannabis dependence, in remission|Cannabis dependence, in remission
C0375175|T048|HT|304.4|ICD9CM|Amphetamine and other psychostimulant dependence|Amphetamine and other psychostimulant dependence
C0375175|T048|AB|304.40|ICD9CM|Amphetamin depend-unspec|Amphetamin depend-unspec
C0375175|T048|PT|304.40|ICD9CM|Amphetamine and other psychostimulant dependence, unspecified|Amphetamine and other psychostimulant dependence, unspecified
C0154492|T048|AB|304.41|ICD9CM|Amphetamin depend-contin|Amphetamin depend-contin
C0154492|T048|PT|304.41|ICD9CM|Amphetamine and other psychostimulant dependence, continuous|Amphetamine and other psychostimulant dependence, continuous
C0154493|T048|AB|304.42|ICD9CM|Amphetamin depend-episod|Amphetamin depend-episod
C0154493|T048|PT|304.42|ICD9CM|Amphetamine and other psychostimulant dependence, episodic|Amphetamine and other psychostimulant dependence, episodic
C0154494|T048|AB|304.43|ICD9CM|Amphetamin depend-remiss|Amphetamin depend-remiss
C0154494|T048|PT|304.43|ICD9CM|Amphetamine and other psychostimulant dependence, in remission|Amphetamine and other psychostimulant dependence, in remission
C0018528|T048|HT|304.5|ICD9CM|Hallucinogen dependence|Hallucinogen dependence
C0018528|T048|AB|304.50|ICD9CM|Hallucinogen dep-unspec|Hallucinogen dep-unspec
C0018528|T048|PT|304.50|ICD9CM|Hallucinogen dependence, unspecified|Hallucinogen dependence, unspecified
C0338749|T048|AB|304.51|ICD9CM|Hallucinogen dep-contin|Hallucinogen dep-contin
C0338749|T048|PT|304.51|ICD9CM|Hallucinogen dependence, continuous|Hallucinogen dependence, continuous
C0338750|T048|AB|304.52|ICD9CM|Hallucinogen dep-episod|Hallucinogen dep-episod
C0338750|T048|PT|304.52|ICD9CM|Hallucinogen dependence, episodic|Hallucinogen dependence, episodic
C0154497|T047|AB|304.53|ICD9CM|Hallucinogen dep-remiss|Hallucinogen dep-remiss
C0154497|T047|PT|304.53|ICD9CM|Hallucinogen dependence, in remission|Hallucinogen dependence, in remission
C0029792|T048|HT|304.6|ICD9CM|Other specified drug dependence|Other specified drug dependence
C0029792|T048|AB|304.60|ICD9CM|Drug depend NEC-unspec|Drug depend NEC-unspec
C0029792|T048|PT|304.60|ICD9CM|Other specified drug dependence, unspecified|Other specified drug dependence, unspecified
C0338738|T048|AB|304.61|ICD9CM|Drug depend NEC-contin|Drug depend NEC-contin
C0338738|T048|PT|304.61|ICD9CM|Other specified drug dependence, continuous|Other specified drug dependence, continuous
C0338739|T048|AB|304.62|ICD9CM|Drug depend NEC-episodic|Drug depend NEC-episodic
C0338739|T048|PT|304.62|ICD9CM|Other specified drug dependence, episodic|Other specified drug dependence, episodic
C0154500|T048|AB|304.63|ICD9CM|Drug depend NEC-in rem|Drug depend NEC-in rem
C0154500|T048|PT|304.63|ICD9CM|Other specified drug dependence, in remission|Other specified drug dependence, in remission
C0154501|T048|HT|304.7|ICD9CM|Combinations of opioid type drug with any other drug dependence|Combinations of opioid type drug with any other drug dependence
C0375176|T048|PT|304.70|ICD9CM|Combinations of opioid type drug with any other drug dependence, unspecified|Combinations of opioid type drug with any other drug dependence, unspecified
C0375176|T048|AB|304.70|ICD9CM|Opioid/other dep-unspec|Opioid/other dep-unspec
C0154502|T048|PT|304.71|ICD9CM|Combinations of opioid type drug with any other drug dependence, continuous|Combinations of opioid type drug with any other drug dependence, continuous
C0154502|T048|AB|304.71|ICD9CM|Opioid/other dep-contin|Opioid/other dep-contin
C0154503|T048|PT|304.72|ICD9CM|Combinations of opioid type drug with any other drug dependence, episodic|Combinations of opioid type drug with any other drug dependence, episodic
C0154503|T048|AB|304.72|ICD9CM|Opioid/other dep-episod|Opioid/other dep-episod
C0154504|T048|PT|304.73|ICD9CM|Combinations of opioid type drug with any other drug dependence, in remission|Combinations of opioid type drug with any other drug dependence, in remission
C0154504|T048|AB|304.73|ICD9CM|Opioid/other dep-remiss|Opioid/other dep-remiss
C0154505|T048|HT|304.8|ICD9CM|Combinations of drug dependence excluding opioid type drug|Combinations of drug dependence excluding opioid type drug
C0375177|T048|AB|304.80|ICD9CM|Comb drug dep NEC-unspec|Comb drug dep NEC-unspec
C0375177|T048|PT|304.80|ICD9CM|Combinations of drug dependence excluding opioid type drug, unspecified|Combinations of drug dependence excluding opioid type drug, unspecified
C0154506|T048|AB|304.81|ICD9CM|Comb drug dep NEC-contin|Comb drug dep NEC-contin
C0154506|T048|PT|304.81|ICD9CM|Combinations of drug dependence excluding opioid type drug, continuous|Combinations of drug dependence excluding opioid type drug, continuous
C0154507|T048|AB|304.82|ICD9CM|Comb drug dep NEC-episod|Comb drug dep NEC-episod
C0154507|T048|PT|304.82|ICD9CM|Combinations of drug dependence excluding opioid type drug, episodic|Combinations of drug dependence excluding opioid type drug, episodic
C0154508|T048|AB|304.83|ICD9CM|Comb drug dep NEC-remiss|Comb drug dep NEC-remiss
C0154508|T048|PT|304.83|ICD9CM|Combinations of drug dependence excluding opioid type drug, in remission|Combinations of drug dependence excluding opioid type drug, in remission
C1510472|T048|HT|304.9|ICD9CM|Unspecified drug dependence|Unspecified drug dependence
C0375178|T048|AB|304.90|ICD9CM|Drug depend NOS-unspec|Drug depend NOS-unspec
C0375178|T048|PT|304.90|ICD9CM|Unspecified drug dependence, unspecified|Unspecified drug dependence, unspecified
C0154509|T048|AB|304.91|ICD9CM|Drug depend NOS-contin|Drug depend NOS-contin
C0154509|T048|PT|304.91|ICD9CM|Unspecified drug dependence, continuous|Unspecified drug dependence, continuous
C0154510|T048|AB|304.92|ICD9CM|Drug depend NOS-episodic|Drug depend NOS-episodic
C0154510|T048|PT|304.92|ICD9CM|Unspecified drug dependence, episodic|Unspecified drug dependence, episodic
C0154511|T048|AB|304.93|ICD9CM|Drug depend NOS-remiss|Drug depend NOS-remiss
C0154511|T048|PT|304.93|ICD9CM|Unspecified drug dependence, in remission|Unspecified drug dependence, in remission
C3665497|T048|HT|305|ICD9CM|Nondependent abuse of drugs|Nondependent abuse of drugs
C0085762|T048|HT|305.0|ICD9CM|Alcohol abuse|Alcohol abuse
C0085762|T048|AB|305.00|ICD9CM|Alcohol abuse-unspec|Alcohol abuse-unspec
C0085762|T048|PT|305.00|ICD9CM|Alcohol abuse, unspecified|Alcohol abuse, unspecified
C1812624|T048|AB|305.01|ICD9CM|Alcohol abuse-continuous|Alcohol abuse-continuous
C1812624|T048|PT|305.01|ICD9CM|Alcohol abuse, continuous|Alcohol abuse, continuous
C0154515|T048|AB|305.02|ICD9CM|Alcohol abuse-episodic|Alcohol abuse-episodic
C0154515|T048|PT|305.02|ICD9CM|Alcohol abuse, episodic|Alcohol abuse, episodic
C0154516|T048|AB|305.03|ICD9CM|Alcohol abuse-in remiss|Alcohol abuse-in remiss
C0154516|T048|PT|305.03|ICD9CM|Alcohol abuse, in remission|Alcohol abuse, in remission
C0040336|T048|AB|305.1|ICD9CM|Tobacco use disorder|Tobacco use disorder
C0040336|T048|PT|305.1|ICD9CM|Tobacco use disorder|Tobacco use disorder
C0006868|T048|HT|305.2|ICD9CM|Cannabis abuse|Cannabis abuse
C0375179|T048|AB|305.20|ICD9CM|Cannabis abuse-unspec|Cannabis abuse-unspec
C0375179|T048|PT|305.20|ICD9CM|Cannabis abuse, unspecified|Cannabis abuse, unspecified
C0154520|T048|AB|305.21|ICD9CM|Cannabis abuse-contin|Cannabis abuse-contin
C0154520|T048|PT|305.21|ICD9CM|Cannabis abuse, continuous|Cannabis abuse, continuous
C0154521|T048|AB|305.22|ICD9CM|Cannabis abuse-episodic|Cannabis abuse-episodic
C0154521|T048|PT|305.22|ICD9CM|Cannabis abuse, episodic|Cannabis abuse, episodic
C0154522|T048|AB|305.23|ICD9CM|Cannabis abuse-in remiss|Cannabis abuse-in remiss
C0154522|T048|PT|305.23|ICD9CM|Cannabis abuse, in remission|Cannabis abuse, in remission
C0018526|T048|HT|305.3|ICD9CM|Hallucinogen abuse|Hallucinogen abuse
C0375180|T048|AB|305.30|ICD9CM|Hallucinog abuse-unspec|Hallucinog abuse-unspec
C0375180|T048|PT|305.30|ICD9CM|Hallucinogen abuse, unspecified|Hallucinogen abuse, unspecified
C0154523|T048|AB|305.31|ICD9CM|Hallucinog abuse-contin|Hallucinog abuse-contin
C0154523|T048|PT|305.31|ICD9CM|Hallucinogen abuse, continuous|Hallucinogen abuse, continuous
C0154524|T048|AB|305.32|ICD9CM|Hallucinog abuse-episod|Hallucinog abuse-episod
C0154524|T048|PT|305.32|ICD9CM|Hallucinogen abuse, episodic|Hallucinogen abuse, episodic
C0154525|T048|AB|305.33|ICD9CM|Hallucinog abuse-remiss|Hallucinog abuse-remiss
C0154525|T048|PT|305.33|ICD9CM|Hallucinogen abuse, in remission|Hallucinogen abuse, in remission
C0036550|T048|HT|305.4|ICD9CM|Sedative, hypnotic or anxiolytic abuse|Sedative, hypnotic or anxiolytic abuse
C0375181|T048|AB|305.40|ICD9CM|Sed,hyp,anxiolytc ab-NOS|Sed,hyp,anxiolytc ab-NOS
C0375181|T048|PT|305.40|ICD9CM|Sedative, hypnotic or anxiolytic abuse, unspecified|Sedative, hypnotic or anxiolytic abuse, unspecified
C0154527|T048|AB|305.41|ICD9CM|Sed,hyp,anxiolytc ab-con|Sed,hyp,anxiolytc ab-con
C0154527|T048|PT|305.41|ICD9CM|Sedative, hypnotic or anxiolytic abuse, continuous|Sedative, hypnotic or anxiolytic abuse, continuous
C0154528|T048|AB|305.42|ICD9CM|Sed,hyp,anxiolytc ab-epi|Sed,hyp,anxiolytc ab-epi
C0154528|T048|PT|305.42|ICD9CM|Sedative, hypnotic or anxiolytic abuse, episodic|Sedative, hypnotic or anxiolytic abuse, episodic
C0154529|T048|AB|305.43|ICD9CM|Sed,hyp,anxiolytc ab-rem|Sed,hyp,anxiolytc ab-rem
C0154529|T048|PT|305.43|ICD9CM|Sedative, hypnotic or anxiolytic abuse, in remission|Sedative, hypnotic or anxiolytic abuse, in remission
C0029095|T048|HT|305.5|ICD9CM|Opioid abuse|Opioid abuse
C0375182|T048|AB|305.50|ICD9CM|Opioid abuse-unspec|Opioid abuse-unspec
C0375182|T048|PT|305.50|ICD9CM|Opioid abuse, unspecified|Opioid abuse, unspecified
C0154530|T048|AB|305.51|ICD9CM|Opioid abuse-continuous|Opioid abuse-continuous
C0154530|T048|PT|305.51|ICD9CM|Opioid abuse, continuous|Opioid abuse, continuous
C0154531|T048|AB|305.52|ICD9CM|Opioid abuse-episodic|Opioid abuse-episodic
C0154531|T048|PT|305.52|ICD9CM|Opioid abuse, episodic|Opioid abuse, episodic
C0154532|T048|AB|305.53|ICD9CM|Opioid abuse-in remiss|Opioid abuse-in remiss
C0154532|T048|PT|305.53|ICD9CM|Opioid abuse, in remission|Opioid abuse, in remission
C0009171|T048|HT|305.6|ICD9CM|Cocaine abuse|Cocaine abuse
C0009171|T048|AB|305.60|ICD9CM|Cocaine abuse-unspec|Cocaine abuse-unspec
C0009171|T048|PT|305.60|ICD9CM|Cocaine abuse, unspecified|Cocaine abuse, unspecified
C0154533|T048|AB|305.61|ICD9CM|Cocaine abuse-continuous|Cocaine abuse-continuous
C0154533|T048|PT|305.61|ICD9CM|Cocaine abuse, continuous|Cocaine abuse, continuous
C0154534|T048|AB|305.62|ICD9CM|Cocaine abuse-episodic|Cocaine abuse-episodic
C0154534|T048|PT|305.62|ICD9CM|Cocaine abuse, episodic|Cocaine abuse, episodic
C0154535|T048|AB|305.63|ICD9CM|Cocaine abuse-in remiss|Cocaine abuse-in remiss
C0154535|T048|PT|305.63|ICD9CM|Cocaine abuse, in remission|Cocaine abuse, in remission
C0154536|T048|HT|305.7|ICD9CM|Amphetamine or related acting sympathomimetic abuse|Amphetamine or related acting sympathomimetic abuse
C0375184|T048|AB|305.70|ICD9CM|Amphetamine abuse-unspec|Amphetamine abuse-unspec
C0375184|T048|PT|305.70|ICD9CM|Amphetamine or related acting sympathomimetic abuse, unspecified|Amphetamine or related acting sympathomimetic abuse, unspecified
C0154537|T048|AB|305.71|ICD9CM|Amphetamine abuse-contin|Amphetamine abuse-contin
C0154537|T048|PT|305.71|ICD9CM|Amphetamine or related acting sympathomimetic abuse, continuous|Amphetamine or related acting sympathomimetic abuse, continuous
C0154538|T048|AB|305.72|ICD9CM|Amphetamine abuse-episod|Amphetamine abuse-episod
C0154538|T048|PT|305.72|ICD9CM|Amphetamine or related acting sympathomimetic abuse, episodic|Amphetamine or related acting sympathomimetic abuse, episodic
C0154539|T048|AB|305.73|ICD9CM|Amphetamine abuse-remiss|Amphetamine abuse-remiss
C0154539|T048|PT|305.73|ICD9CM|Amphetamine or related acting sympathomimetic abuse, in remission|Amphetamine or related acting sympathomimetic abuse, in remission
C0154540|T048|HT|305.8|ICD9CM|Antidepressant type abuse|Antidepressant type abuse
C0375185|T048|AB|305.80|ICD9CM|Antidepress abuse-unspec|Antidepress abuse-unspec
C0375185|T048|PT|305.80|ICD9CM|Antidepressant type abuse, unspecified|Antidepressant type abuse, unspecified
C0154541|T048|AB|305.81|ICD9CM|Antidepress abuse-contin|Antidepress abuse-contin
C0154541|T048|PT|305.81|ICD9CM|Antidepressant type abuse, continuous|Antidepressant type abuse, continuous
C0154542|T048|AB|305.82|ICD9CM|Antidepress abuse-episod|Antidepress abuse-episod
C0154542|T048|PT|305.82|ICD9CM|Antidepressant type abuse, episodic|Antidepressant type abuse, episodic
C0154543|T048|AB|305.83|ICD9CM|Antidepress abuse-remiss|Antidepress abuse-remiss
C0154543|T048|PT|305.83|ICD9CM|Antidepressant type abuse, in remission|Antidepressant type abuse, in remission
C0154544|T048|HT|305.9|ICD9CM|Other, mixed, or unspecified drug abuse|Other, mixed, or unspecified drug abuse
C0154544|T048|AB|305.90|ICD9CM|Drug abuse NEC-unspec|Drug abuse NEC-unspec
C0154544|T048|PT|305.90|ICD9CM|Other, mixed, or unspecified drug abuse, unspecified|Other, mixed, or unspecified drug abuse, unspecified
C0154545|T048|AB|305.91|ICD9CM|Drug abuse NEC-contin|Drug abuse NEC-contin
C0154545|T048|PT|305.91|ICD9CM|Other, mixed, or unspecified drug abuse, continuous|Other, mixed, or unspecified drug abuse, continuous
C0154546|T048|AB|305.92|ICD9CM|Drug abuse NEC-episodic|Drug abuse NEC-episodic
C0154546|T048|PT|305.92|ICD9CM|Other, mixed, or unspecified drug abuse, episodic|Other, mixed, or unspecified drug abuse, episodic
C0154547|T048|AB|305.93|ICD9CM|Drug abuse NEC-in remiss|Drug abuse NEC-in remiss
C0154547|T048|PT|305.93|ICD9CM|Other, mixed, or unspecified drug abuse, in remission|Other, mixed, or unspecified drug abuse, in remission
C0154548|T047|HT|306|ICD9CM|Physiological malfunction arising from mental factors|Physiological malfunction arising from mental factors
C0154549|T048|PT|306.0|ICD9CM|Musculoskeletal malfunction arising from mental factors|Musculoskeletal malfunction arising from mental factors
C0154549|T048|AB|306.0|ICD9CM|Psychogen musculskel dis|Psychogen musculskel dis
C0338945|T048|AB|306.1|ICD9CM|Psychogenic respir dis|Psychogenic respir dis
C0338945|T048|PT|306.1|ICD9CM|Respiratory malfunction arising from mental factors|Respiratory malfunction arising from mental factors
C0027821|T047|PT|306.2|ICD9CM|Cardiovascular malfunction arising from mental factors|Cardiovascular malfunction arising from mental factors
C0027821|T047|AB|306.2|ICD9CM|Psychogen cardiovasc dis|Psychogen cardiovasc dis
C0154551|T048|AB|306.3|ICD9CM|Psychogenic skin disease|Psychogenic skin disease
C0154551|T048|PT|306.3|ICD9CM|Skin disorder arising from mental factors|Skin disorder arising from mental factors
C0017183|T048|PT|306.4|ICD9CM|Gastrointestinal malfunction arising from mental factors|Gastrointestinal malfunction arising from mental factors
C0017183|T048|AB|306.4|ICD9CM|Psychogenic GI disease|Psychogenic GI disease
C0154552|T047|HT|306.5|ICD9CM|Genitourinary malfunction arising from mental factors|Genitourinary malfunction arising from mental factors
C0837158|T048|PT|306.50|ICD9CM|Psychogenic genitourinary malfunction, unspecified|Psychogenic genitourinary malfunction, unspecified
C0837158|T048|AB|306.50|ICD9CM|Psychogenic gu dis NOS|Psychogenic gu dis NOS
C0042266|T048|AB|306.51|ICD9CM|Psychogenic vaginismus|Psychogenic vaginismus
C0042266|T048|PT|306.51|ICD9CM|Psychogenic vaginismus|Psychogenic vaginismus
C0154555|T048|AB|306.52|ICD9CM|Psychogenic dysmenorrhea|Psychogenic dysmenorrhea
C0154555|T048|PT|306.52|ICD9CM|Psychogenic dysmenorrhea|Psychogenic dysmenorrhea
C0232857|T184|AB|306.53|ICD9CM|Psychogenic dysuria|Psychogenic dysuria
C0232857|T184|PT|306.53|ICD9CM|Psychogenic dysuria|Psychogenic dysuria
C0154557|T047|PT|306.59|ICD9CM|Other genitourinary malfunction arising from mental factors|Other genitourinary malfunction arising from mental factors
C0154557|T047|AB|306.59|ICD9CM|Psychogenic gu dis NEC|Psychogenic gu dis NEC
C0154558|T047|PT|306.6|ICD9CM|Endocrine disorder arising from mental factors|Endocrine disorder arising from mental factors
C0154558|T047|AB|306.6|ICD9CM|Psychogen endocrine dis|Psychogen endocrine dis
C0154559|T047|PT|306.7|ICD9CM|Disorder of organs of special sense arising from mental factors|Disorder of organs of special sense arising from mental factors
C0154559|T047|AB|306.7|ICD9CM|Psychogenic sensory dis|Psychogenic sensory dis
C0029824|T048|PT|306.8|ICD9CM|Other specified psychophysiological malfunction|Other specified psychophysiological malfunction
C0029824|T048|AB|306.8|ICD9CM|Psychogenic disorder NEC|Psychogenic disorder NEC
C0041876|T048|AB|306.9|ICD9CM|Psychogenic disorder NOS|Psychogenic disorder NOS
C0041876|T048|PT|306.9|ICD9CM|Unspecified psychophysiological malfunction|Unspecified psychophysiological malfunction
C0302370|T047|HT|307|ICD9CM|Special symptoms or syndromes, not elsewhere classified|Special symptoms or syndromes, not elsewhere classified
C2921027|T048|AB|307.0|ICD9CM|Adult onset flncy disord|Adult onset flncy disord
C2921027|T048|PT|307.0|ICD9CM|Adult onset fluency disorder|Adult onset fluency disorder
C0003125|T048|AB|307.1|ICD9CM|Anorexia nervosa|Anorexia nervosa
C0003125|T048|PT|307.1|ICD9CM|Anorexia nervosa|Anorexia nervosa
C0040188|T048|HT|307.2|ICD9CM|Tics|Tics
C0040188|T048|AB|307.20|ICD9CM|Tic disorder NOS|Tic disorder NOS
C0040188|T048|PT|307.20|ICD9CM|Tic disorder, unspecified|Tic disorder, unspecified
C0040702|T048|AB|307.21|ICD9CM|Transient tic disorder|Transient tic disorder
C0040702|T048|PT|307.21|ICD9CM|Transient tic disorder|Transient tic disorder
C0008701|T048|AB|307.22|ICD9CM|Chr motor/vocal tic dis|Chr motor/vocal tic dis
C0008701|T048|PT|307.22|ICD9CM|Chronic motor or vocal tic disorder|Chronic motor or vocal tic disorder
C0040517|T047|AB|307.23|ICD9CM|Tourette's disorder|Tourette's disorder
C0040517|T047|PT|307.23|ICD9CM|Tourette's disorder|Tourette's disorder
C0038273|T048|AB|307.3|ICD9CM|Stereotypic movement dis|Stereotypic movement dis
C0038273|T048|PT|307.3|ICD9CM|Stereotypic movement disorder|Stereotypic movement disorder
C0154564|T048|HT|307.4|ICD9CM|Specific disorders of sleep of nonorganic origin|Specific disorders of sleep of nonorganic origin
C0154565|T048|AB|307.40|ICD9CM|Nonorganic sleep dis NOS|Nonorganic sleep dis NOS
C0154565|T048|PT|307.40|ICD9CM|Nonorganic sleep disorder, unspecified|Nonorganic sleep disorder, unspecified
C0154566|T048|PT|307.41|ICD9CM|Transient disorder of initiating or maintaining sleep|Transient disorder of initiating or maintaining sleep
C0154566|T048|AB|307.41|ICD9CM|Transient insomnia|Transient insomnia
C0868777|T048|PT|307.42|ICD9CM|Persistent disorder of initiating or maintaining sleep|Persistent disorder of initiating or maintaining sleep
C0868777|T048|AB|307.42|ICD9CM|Persistent insomnia|Persistent insomnia
C0154568|T048|PT|307.43|ICD9CM|Transient disorder of initiating or maintaining wakefulness|Transient disorder of initiating or maintaining wakefulness
C0154568|T048|AB|307.43|ICD9CM|Transient hypersomnia|Transient hypersomnia
C0154569|T048|PT|307.44|ICD9CM|Persistent disorder of initiating or maintaining wakefulness|Persistent disorder of initiating or maintaining wakefulness
C0154569|T048|AB|307.44|ICD9CM|Persistent hypersomnia|Persistent hypersomnia
C1561844|T048|PT|307.45|ICD9CM|Circadian rhythm sleep disorder of nonorganic origin|Circadian rhythm sleep disorder of nonorganic origin
C1561844|T048|AB|307.45|ICD9CM|Nonorganic circadian rhy|Nonorganic circadian rhy
C0752294|T047|AB|307.46|ICD9CM|Sleep arousal disorder|Sleep arousal disorder
C0752294|T047|PT|307.46|ICD9CM|Sleep arousal disorder|Sleep arousal disorder
C0154571|T048|PT|307.47|ICD9CM|Other dysfunctions of sleep stages or arousal from sleep|Other dysfunctions of sleep stages or arousal from sleep
C0154571|T048|AB|307.47|ICD9CM|Sleep stage dysfunc NEC|Sleep stage dysfunc NEC
C0154572|T048|AB|307.48|ICD9CM|Repetit sleep intrusion|Repetit sleep intrusion
C0154572|T048|PT|307.48|ICD9CM|Repetitive intrusions of sleep|Repetitive intrusions of sleep
C0154573|T048|AB|307.49|ICD9CM|Nonorganic sleep dis NEC|Nonorganic sleep dis NEC
C0154573|T048|PT|307.49|ICD9CM|Other specific disorders of sleep of nonorganic origin|Other specific disorders of sleep of nonorganic origin
C0029587|T048|HT|307.5|ICD9CM|Other and unspecified disorders of eating|Other and unspecified disorders of eating
C0013473|T048|AB|307.50|ICD9CM|Eating disorder NOS|Eating disorder NOS
C0013473|T048|PT|307.50|ICD9CM|Eating disorder, unspecified|Eating disorder, unspecified
C2267227|T048|AB|307.51|ICD9CM|Bulimia nervosa|Bulimia nervosa
C2267227|T048|PT|307.51|ICD9CM|Bulimia nervosa|Bulimia nervosa
C0031873|T048|AB|307.52|ICD9CM|Pica|Pica
C0031873|T048|PT|307.52|ICD9CM|Pica|Pica
C0154575|T048|AB|307.53|ICD9CM|Rumination disorder|Rumination disorder
C0154575|T048|PT|307.53|ICD9CM|Rumination disorder|Rumination disorder
C0233757|T048|AB|307.54|ICD9CM|Psychogenic vomiting|Psychogenic vomiting
C0233757|T048|PT|307.54|ICD9CM|Psychogenic vomiting|Psychogenic vomiting
C0029587|T048|AB|307.59|ICD9CM|Eating disorder NEC|Eating disorder NEC
C0029587|T048|PT|307.59|ICD9CM|Other disorders of eating|Other disorders of eating
C0014394|T047|AB|307.6|ICD9CM|Enuresis|Enuresis
C0014394|T047|PT|307.6|ICD9CM|Enuresis|Enuresis
C0014089|T048|AB|307.7|ICD9CM|Encopresis|Encopresis
C0014089|T048|PT|307.7|ICD9CM|Encopresis|Encopresis
C1456322|T048|HT|307.8|ICD9CM|Pain disorders related to psychological factors|Pain disorders related to psychological factors
C0152174|T048|AB|307.80|ICD9CM|Psychogenic pain NOS|Psychogenic pain NOS
C0152174|T048|PT|307.80|ICD9CM|Psychogenic pain, site unspecified|Psychogenic pain, site unspecified
C0033893|T047|AB|307.81|ICD9CM|Tension headache|Tension headache
C0033893|T047|PT|307.81|ICD9CM|Tension headache|Tension headache
C1456321|T048|PT|307.89|ICD9CM|Other pain disorders related to psychological factors|Other pain disorders related to psychological factors
C1456321|T048|AB|307.89|ICD9CM|Psychogenic pain NEC|Psychogenic pain NEC
C0302371|T048|PT|307.9|ICD9CM|Other and unspecified special symptoms or syndromes, not elsewhere classified|Other and unspecified special symptoms or syndromes, not elsewhere classified
C0302371|T048|AB|307.9|ICD9CM|Special symptom NEC/NOS|Special symptom NEC/NOS
C0236816|T048|HT|308|ICD9CM|Acute reaction to stress|Acute reaction to stress
C0154578|T048|PT|308.0|ICD9CM|Predominant disturbance of emotions|Predominant disturbance of emotions
C0154578|T048|AB|308.0|ICD9CM|Stress react, emotional|Stress react, emotional
C0154579|T048|PT|308.1|ICD9CM|Predominant disturbance of consciousness|Predominant disturbance of consciousness
C0154579|T048|AB|308.1|ICD9CM|Stress reaction, fugue|Stress reaction, fugue
C0154580|T048|PT|308.2|ICD9CM|Predominant psychomotor disturbance|Predominant psychomotor disturbance
C0154580|T048|AB|308.2|ICD9CM|Stress react, psychomot|Stress react, psychomot
C0029488|T048|AB|308.3|ICD9CM|Acute stress react NEC|Acute stress react NEC
C0029488|T048|PT|308.3|ICD9CM|Other acute reactions to stress|Other acute reactions to stress
C0154581|T048|PT|308.4|ICD9CM|Mixed disorders as reaction to stress|Mixed disorders as reaction to stress
C0154581|T048|AB|308.4|ICD9CM|Stress react, mixed dis|Stress react, mixed dis
C0236816|T048|AB|308.9|ICD9CM|Acute stress react NOS|Acute stress react NOS
C0236816|T048|PT|308.9|ICD9CM|Unspecified acute reaction to stress|Unspecified acute reaction to stress
C0040701|T048|HT|309|ICD9CM|Adjustment reaction|Adjustment reaction
C0001539|T048|PT|309.0|ICD9CM|Adjustment disorder with depressed mood|Adjustment disorder with depressed mood
C0001539|T048|AB|309.0|ICD9CM|Adjustmnt dis w depressn|Adjustmnt dis w depressn
C0154583|T048|AB|309.1|ICD9CM|Prolong depressive react|Prolong depressive react
C0154583|T048|PT|309.1|ICD9CM|Prolonged depressive reaction|Prolonged depressive reaction
C0154584|T048|HT|309.2|ICD9CM|Adjustment reaction with predominant disturbance of other emotions|Adjustment reaction with predominant disturbance of other emotions
C0003477|T048|AB|309.21|ICD9CM|Separation anxiety|Separation anxiety
C0003477|T048|PT|309.21|ICD9CM|Separation anxiety disorder|Separation anxiety disorder
C0154585|T048|AB|309.22|ICD9CM|Emancipation disorder|Emancipation disorder
C0154585|T048|PT|309.22|ICD9CM|Emancipation disorder of adolescence and early adult life|Emancipation disorder of adolescence and early adult life
C0154586|T048|AB|309.23|ICD9CM|Academic/work inhibition|Academic/work inhibition
C0154586|T048|PT|309.23|ICD9CM|Specific academic or work inhibition|Specific academic or work inhibition
C0154587|T048|AB|309.24|ICD9CM|Adjustment dis w anxiety|Adjustment dis w anxiety
C0154587|T048|PT|309.24|ICD9CM|Adjustment disorder with anxiety|Adjustment disorder with anxiety
C0154588|T048|AB|309.28|ICD9CM|Adjust dis w anxiety/dep|Adjust dis w anxiety/dep
C0154588|T048|PT|309.28|ICD9CM|Adjustment disorder with mixed anxiety and depressed mood|Adjustment disorder with mixed anxiety and depressed mood
C0154589|T048|AB|309.29|ICD9CM|Adj react-emotion NEC|Adj react-emotion NEC
C0154589|T048|PT|309.29|ICD9CM|Other adjustment reactions with predominant disturbance of other emotions|Other adjustment reactions with predominant disturbance of other emotions
C0001540|T048|AB|309.3|ICD9CM|Adjust disor/dis conduct|Adjust disor/dis conduct
C0001540|T048|PT|309.3|ICD9CM|Adjustment disorder with disturbance of conduct|Adjustment disorder with disturbance of conduct
C0001541|T048|AB|309.4|ICD9CM|Adj dis-emotion/conduct|Adj dis-emotion/conduct
C0001541|T048|PT|309.4|ICD9CM|Adjustment disorder with mixed disturbance of emotions and conduct|Adjustment disorder with mixed disturbance of emotions and conduct
C0154592|T048|HT|309.8|ICD9CM|Other specified adjustment reactions|Other specified adjustment reactions
C0038436|T048|AB|309.81|ICD9CM|Posttraumatic stress dis|Posttraumatic stress dis
C0038436|T048|PT|309.81|ICD9CM|Posttraumatic stress disorder|Posttraumatic stress disorder
C0154594|T048|AB|309.82|ICD9CM|Adjust react-phys sympt|Adjust react-phys sympt
C0154594|T048|PT|309.82|ICD9CM|Adjustment reaction with physical symptoms|Adjustment reaction with physical symptoms
C0154595|T048|AB|309.83|ICD9CM|Adjust react-withdrawal|Adjust react-withdrawal
C0154595|T048|PT|309.83|ICD9CM|Adjustment reaction with withdrawal|Adjustment reaction with withdrawal
C0154592|T048|AB|309.89|ICD9CM|Adjustment reaction NEC|Adjustment reaction NEC
C0154592|T048|PT|309.89|ICD9CM|Other specified adjustment reactions|Other specified adjustment reactions
C0040701|T048|AB|309.9|ICD9CM|Adjustment reaction NOS|Adjustment reaction NOS
C0040701|T048|PT|309.9|ICD9CM|Unspecified adjustment reaction|Unspecified adjustment reaction
C1456324|T048|HT|310|ICD9CM|Specific nonpsychotic mental disorders due to brain damage|Specific nonpsychotic mental disorders due to brain damage
C0549117|T047|AB|310.0|ICD9CM|Frontal lobe syndrome|Frontal lobe syndrome
C0549117|T047|PT|310.0|ICD9CM|Frontal lobe syndrome|Frontal lobe syndrome
C1456323|T048|PT|310.1|ICD9CM|Personality change due to conditions classified elsewhere|Personality change due to conditions classified elsewhere
C1456323|T048|AB|310.1|ICD9CM|Personality chg oth dis|Personality chg oth dis
C0546983|T047|AB|310.2|ICD9CM|Postconcussion syndrome|Postconcussion syndrome
C0546983|T047|PT|310.2|ICD9CM|Postconcussion syndrome|Postconcussion syndrome
C0154598|T048|HT|310.8|ICD9CM|Other specified nonpsychotic mental disorders following organic brain damage|Other specified nonpsychotic mental disorders following organic brain damage
C2316460|T048|AB|310.81|ICD9CM|Pseudobulbar affect|Pseudobulbar affect
C2316460|T048|PT|310.81|ICD9CM|Pseudobulbar affect|Pseudobulbar affect
C0154598|T048|AB|310.89|ICD9CM|Nonpsych mntl disord NEC|Nonpsych mntl disord NEC
C0154598|T048|PT|310.89|ICD9CM|Other specified nonpsychotic mental disorders following organic brain damage|Other specified nonpsychotic mental disorders following organic brain damage
C0041862|T048|AB|310.9|ICD9CM|Nonpsychot brain syn NOS|Nonpsychot brain syn NOS
C0041862|T048|PT|310.9|ICD9CM|Unspecified nonpsychotic mental disorder following organic brain damage|Unspecified nonpsychotic mental disorder following organic brain damage
C0868892|T048|AB|311|ICD9CM|Depressive disorder NEC|Depressive disorder NEC
C0868892|T048|PT|311|ICD9CM|Depressive disorder, not elsewhere classified|Depressive disorder, not elsewhere classified
C0869273|T048|HT|312|ICD9CM|Disturbance of conduct, not elsewhere classified|Disturbance of conduct, not elsewhere classified
C0041665|T048|HT|312.0|ICD9CM|Undersocialized conduct disorder, aggressive type|Undersocialized conduct disorder, aggressive type
C0375189|T048|PT|312.00|ICD9CM|Undersocialized conduct disorder, aggressive type, unspecified|Undersocialized conduct disorder, aggressive type, unspecified
C0375189|T048|AB|312.00|ICD9CM|Unsocial aggress-unspec|Unsocial aggress-unspec
C0154600|T048|PT|312.01|ICD9CM|Undersocialized conduct disorder, aggressive type, mild|Undersocialized conduct disorder, aggressive type, mild
C0154600|T048|AB|312.01|ICD9CM|Unsocial aggression-mild|Unsocial aggression-mild
C0154601|T048|PT|312.02|ICD9CM|Undersocialized conduct disorder, aggressive type, moderate|Undersocialized conduct disorder, aggressive type, moderate
C0154601|T048|AB|312.02|ICD9CM|Unsocial aggression-mod|Unsocial aggression-mod
C0154602|T048|PT|312.03|ICD9CM|Undersocialized conduct disorder, aggressive type, severe|Undersocialized conduct disorder, aggressive type, severe
C0154602|T048|AB|312.03|ICD9CM|Unsocial aggress-severe|Unsocial aggress-severe
C0154603|T048|HT|312.1|ICD9CM|Undersocialized conduct disorder, unaggressive type|Undersocialized conduct disorder, unaggressive type
C0375190|T048|PT|312.10|ICD9CM|Undersocialized conduct disorder, unaggressive type, unspecified|Undersocialized conduct disorder, unaggressive type, unspecified
C0375190|T048|AB|312.10|ICD9CM|Unsocial unaggress-unsp|Unsocial unaggress-unsp
C0154604|T048|PT|312.11|ICD9CM|Undersocialized conduct disorder, unaggressive type, mild|Undersocialized conduct disorder, unaggressive type, mild
C0154604|T048|AB|312.11|ICD9CM|Unsocial unaggress-mild|Unsocial unaggress-mild
C0154605|T048|PT|312.12|ICD9CM|Undersocialized conduct disorder, unaggressive type, moderate|Undersocialized conduct disorder, unaggressive type, moderate
C0154605|T048|AB|312.12|ICD9CM|Unsocial unaggress-mod|Unsocial unaggress-mod
C0154606|T048|PT|312.13|ICD9CM|Undersocialized conduct disorder, unaggressive type, severe|Undersocialized conduct disorder, unaggressive type, severe
C0154606|T048|AB|312.13|ICD9CM|Unsocial unaggr-severe|Unsocial unaggr-severe
C0037448|T048|HT|312.2|ICD9CM|Socialized conduct disorder|Socialized conduct disorder
C0037448|T048|AB|312.20|ICD9CM|Social conduct dis-unsp|Social conduct dis-unsp
C0037448|T048|PT|312.20|ICD9CM|Socialized conduct disorder, unspecified|Socialized conduct disorder, unspecified
C2231357|T048|AB|312.21|ICD9CM|Social conduct dis-mild|Social conduct dis-mild
C2231357|T048|PT|312.21|ICD9CM|Socialized conduct disorder, mild|Socialized conduct disorder, mild
C2197988|T048|AB|312.22|ICD9CM|Social conduct dis-mod|Social conduct dis-mod
C2197988|T048|PT|312.22|ICD9CM|Socialized conduct disorder, moderate|Socialized conduct disorder, moderate
C2231358|T048|AB|312.23|ICD9CM|Social conduct dis-sev|Social conduct dis-sev
C2231358|T048|PT|312.23|ICD9CM|Socialized conduct disorder, severe|Socialized conduct disorder, severe
C0868739|T048|HT|312.3|ICD9CM|Disorders of impulse control, not elsewhere classified|Disorders of impulse control, not elsewhere classified
C0021122|T048|AB|312.30|ICD9CM|Impulse control dis NOS|Impulse control dis NOS
C0021122|T048|PT|312.30|ICD9CM|Impulse control disorder, unspecified|Impulse control disorder, unspecified
C0030662|T048|AB|312.31|ICD9CM|Pathological gambling|Pathological gambling
C0030662|T048|PT|312.31|ICD9CM|Pathological gambling|Pathological gambling
C0022734|T048|AB|312.32|ICD9CM|Kleptomania|Kleptomania
C0022734|T048|PT|312.32|ICD9CM|Kleptomania|Kleptomania
C0016142|T048|AB|312.33|ICD9CM|Pyromania|Pyromania
C0016142|T048|PT|312.33|ICD9CM|Pyromania|Pyromania
C0021776|T048|AB|312.34|ICD9CM|Intermitt explosive dis|Intermitt explosive dis
C0021776|T048|PT|312.34|ICD9CM|Intermittent explosive disorder|Intermittent explosive disorder
C0154610|T048|AB|312.35|ICD9CM|Isolated explosive dis|Isolated explosive dis
C0154610|T048|PT|312.35|ICD9CM|Isolated explosive disorder|Isolated explosive disorder
C0029588|T048|AB|312.39|ICD9CM|Impulse control dis NEC|Impulse control dis NEC
C0029588|T048|PT|312.39|ICD9CM|Other disorders of impulse control|Other disorders of impulse control
C0494432|T048|AB|312.4|ICD9CM|Mix dis conduct/emotion|Mix dis conduct/emotion
C0494432|T048|PT|312.4|ICD9CM|Mixed disturbance of conduct and emotions|Mixed disturbance of conduct and emotions
C0302373|T048|HT|312.8|ICD9CM|Other specified disturbances of conduct, not elsewhere classified|Other specified disturbances of conduct, not elsewhere classified
C0339005|T048|AB|312.81|ICD9CM|Cndct dsrdr chldhd onst|Cndct dsrdr chldhd onst
C0339005|T048|PT|312.81|ICD9CM|Conduct disorder, childhood onset type|Conduct disorder, childhood onset type
C0375192|T048|AB|312.82|ICD9CM|Cndct dsrdr adlscnt onst|Cndct dsrdr adlscnt onst
C0375192|T048|PT|312.82|ICD9CM|Conduct disorder, adolescent onset type|Conduct disorder, adolescent onset type
C0375193|T048|AB|312.89|ICD9CM|Other conduct disorder|Other conduct disorder
C0375193|T048|PT|312.89|ICD9CM|Other conduct disorder|Other conduct disorder
C0149654|T048|AB|312.9|ICD9CM|Conduct disturbance NOS|Conduct disturbance NOS
C0149654|T048|PT|312.9|ICD9CM|Unspecified disturbance of conduct|Unspecified disturbance of conduct
C0154613|T048|HT|313|ICD9CM|Disturbance of emotions specific to childhood and adolescence|Disturbance of emotions specific to childhood and adolescence
C0270307|T048|AB|313.0|ICD9CM|Overanxious disorder|Overanxious disorder
C0270307|T048|PT|313.0|ICD9CM|Overanxious disorder specific to childhood and adolescence|Overanxious disorder specific to childhood and adolescence
C0154614|T048|AB|313.1|ICD9CM|Misery & unhappiness dis|Misery & unhappiness dis
C0154614|T048|PT|313.1|ICD9CM|Misery and unhappiness disorder specific to childhood and adolescence|Misery and unhappiness disorder specific to childhood and adolescence
C0154615|T048|HT|313.2|ICD9CM|Sensitivity, shyness, and social withdrawal disorder specific to childhood and adolescence|Sensitivity, shyness, and social withdrawal disorder specific to childhood and adolescence
C0154616|T048|PT|313.21|ICD9CM|Shyness disorder of childhood|Shyness disorder of childhood
C0154616|T048|AB|313.21|ICD9CM|Shyness disorder-child|Shyness disorder-child
C0546819|T048|AB|313.22|ICD9CM|Introverted dis-child|Introverted dis-child
C0546819|T048|PT|313.22|ICD9CM|Introverted disorder of childhood|Introverted disorder of childhood
C1456326|T048|AB|313.23|ICD9CM|Selective mutism|Selective mutism
C1456326|T048|PT|313.23|ICD9CM|Selective mutism|Selective mutism
C0154618|T048|AB|313.3|ICD9CM|Relationship problems|Relationship problems
C0154618|T048|PT|313.3|ICD9CM|Relationship problems specific to childhood and adolescence|Relationship problems specific to childhood and adolescence
C0154619|T048|HT|313.8|ICD9CM|Other or mixed emotional disturbances of childhood or adolescence|Other or mixed emotional disturbances of childhood or adolescence
C0029121|T048|AB|313.81|ICD9CM|Opposition defiant disor|Opposition defiant disor
C0029121|T048|PT|313.81|ICD9CM|Oppositional defiant disorder|Oppositional defiant disorder
C0020795|T048|AB|313.82|ICD9CM|Identity disorder|Identity disorder
C0020795|T048|PT|313.82|ICD9CM|Identity disorder of childhood or adolescence|Identity disorder of childhood or adolescence
C0154621|T048|PT|313.83|ICD9CM|Academic underachievement disorder of childhood or adolescence|Academic underachievement disorder of childhood or adolescence
C0154621|T048|AB|313.83|ICD9CM|Academic underachievment|Academic underachievment
C0154622|T048|AB|313.89|ICD9CM|Emotional dis child NEC|Emotional dis child NEC
C0154622|T048|PT|313.89|ICD9CM|Other emotional disturbances of childhood or adolescence|Other emotional disturbances of childhood or adolescence
C0154623|T048|AB|313.9|ICD9CM|Emotional dis child NOS|Emotional dis child NOS
C0154623|T048|PT|313.9|ICD9CM|Unspecified emotional disturbance of childhood or adolescence|Unspecified emotional disturbance of childhood or adolescence
C1263846|T048|HT|314|ICD9CM|Hyperkinetic syndrome of childhood|Hyperkinetic syndrome of childhood
C0004269|T047|HT|314.0|ICD9CM|Attention deficit disorder of childhood|Attention deficit disorder of childhood
C0339002|T048|PT|314.00|ICD9CM|Attention deficit disorder without mention of hyperactivity|Attention deficit disorder without mention of hyperactivity
C0339002|T048|AB|314.00|ICD9CM|Attn defic nonhyperact|Attn defic nonhyperact
C1263846|T048|PT|314.01|ICD9CM|Attention deficit disorder with hyperactivity|Attention deficit disorder with hyperactivity
C1263846|T048|AB|314.01|ICD9CM|Attn deficit w hyperact|Attn deficit w hyperact
C0154627|T048|PT|314.1|ICD9CM|Hyperkinesis with developmental delay|Hyperkinesis with developmental delay
C0154627|T048|AB|314.1|ICD9CM|Hyperkinet w devel delay|Hyperkinet w devel delay
C0154628|T048|AB|314.2|ICD9CM|Hyperkinetic conduct dis|Hyperkinetic conduct dis
C0154628|T048|PT|314.2|ICD9CM|Hyperkinetic conduct disorder|Hyperkinetic conduct disorder
C0154629|T048|AB|314.8|ICD9CM|Other hyperkinetic synd|Other hyperkinetic synd
C0154629|T048|PT|314.8|ICD9CM|Other specified manifestations of hyperkinetic syndrome|Other specified manifestations of hyperkinetic syndrome
C1263846|T048|AB|314.9|ICD9CM|Hyperkinetic synd NOS|Hyperkinetic synd NOS
C1263846|T048|PT|314.9|ICD9CM|Unspecified hyperkinetic syndrome|Unspecified hyperkinetic syndrome
C0037785|T048|HT|315|ICD9CM|Specific delays in development|Specific delays in development
C0920296|T048|HT|315.0|ICD9CM|Developmental reading disorder|Developmental reading disorder
C0920296|T048|PT|315.00|ICD9CM|Developmental reading disorder, unspecified|Developmental reading disorder, unspecified
C0920296|T048|AB|315.00|ICD9CM|Reading disorder NOS|Reading disorder NOS
C0002018|T048|AB|315.01|ICD9CM|Alexia|Alexia
C0002018|T048|PT|315.01|ICD9CM|Alexia|Alexia
C0920296|T048|AB|315.02|ICD9CM|Developmental dyslexia|Developmental dyslexia
C0920296|T048|PT|315.02|ICD9CM|Developmental dyslexia|Developmental dyslexia
C0154631|T048|PT|315.09|ICD9CM|Other specific developmental reading disorder|Other specific developmental reading disorder
C0154631|T048|AB|315.09|ICD9CM|Reading disorder NEC|Reading disorder NEC
C1411876|T048|AB|315.1|ICD9CM|Mathematics disorder|Mathematics disorder
C1411876|T048|PT|315.1|ICD9CM|Mathematics disorder|Mathematics disorder
C0338982|T048|AB|315.2|ICD9CM|Oth learning difficulty|Oth learning difficulty
C0338982|T048|PT|315.2|ICD9CM|Other specific developmental learning difficulties|Other specific developmental learning difficulties
C0154632|T048|HT|315.3|ICD9CM|Developmental speech or language disorder|Developmental speech or language disorder
C0236826|T048|AB|315.31|ICD9CM|Expressive language dis|Expressive language dis
C0236826|T048|PT|315.31|ICD9CM|Expressive language disorder|Expressive language disorder
C0236827|T048|PT|315.32|ICD9CM|Mixed receptive-expressive language disorder|Mixed receptive-expressive language disorder
C0236827|T048|AB|315.32|ICD9CM|Recp-expres language dis|Recp-expres language dis
C1955750|T048|PT|315.34|ICD9CM|Speech and language developmental delay due to hearing loss|Speech and language developmental delay due to hearing loss
C1955750|T048|AB|315.34|ICD9CM|Speech del d/t hear loss|Speech del d/t hear loss
C2921028|T048|PT|315.35|ICD9CM|Childhood onset fluency disorder|Childhood onset fluency disorder
C2921028|T048|AB|315.35|ICD9CM|Chldhd onset flncy disor|Chldhd onset flncy disor
C0154633|T048|PT|315.39|ICD9CM|Other developmental speech or language disorder|Other developmental speech or language disorder
C0154633|T048|AB|315.39|ICD9CM|Speech/language dis NEC|Speech/language dis NEC
C0011757|T048|AB|315.4|ICD9CM|Devel coordination dis|Devel coordination dis
C0011757|T048|PT|315.4|ICD9CM|Developmental coordination disorder|Developmental coordination disorder
C0154634|T048|AB|315.5|ICD9CM|Mixed development dis|Mixed development dis
C0154634|T048|PT|315.5|ICD9CM|Mixed development disorder|Mixed development disorder
C0154635|T048|AB|315.8|ICD9CM|Development delays NEC|Development delays NEC
C0154635|T048|PT|315.8|ICD9CM|Other specified delays in development|Other specified delays in development
C0424605|T048|AB|315.9|ICD9CM|Development delay NOS|Development delay NOS
C0424605|T048|PT|315.9|ICD9CM|Unspecified delay in development|Unspecified delay in development
C0154637|T048|AB|316|ICD9CM|Psychic factor w oth dis|Psychic factor w oth dis
C0154637|T048|PT|316|ICD9CM|Psychic factors associated with diseases classified elsewhere|Psychic factors associated with diseases classified elsewhere
C0026106|T048|AB|317|ICD9CM|Mild intellect disabilty|Mild intellect disabilty
C0026106|T048|PT|317|ICD9CM|Mild intellectual disabilities|Mild intellectual disabilities
C3714756|T048|HT|317-319.99|ICD9CM|INTELLECTUAL DISABILITIES|INTELLECTUAL DISABILITIES
C3161382|T048|HT|318|ICD9CM|Other specified intellectual disabilities|Other specified intellectual disabilities
C0026351|T048|AB|318.0|ICD9CM|Mod intellect disability|Mod intellect disability
C0026351|T048|PT|318.0|ICD9CM|Moderate intellectual disabilities|Moderate intellectual disabilities
C0036857|T048|AB|318.1|ICD9CM|Sev intellect disability|Sev intellect disability
C0036857|T048|PT|318.1|ICD9CM|Severe intellectual disabilities|Severe intellectual disabilities
C3161330|T048|AB|318.2|ICD9CM|Profnd intellct disablty|Profnd intellct disablty
C3161330|T048|PT|318.2|ICD9CM|Profound intellectual disabilities|Profound intellectual disabilities
C3161331|T048|AB|319|ICD9CM|Intellect disability NOS|Intellect disability NOS
C3161331|T048|PT|319|ICD9CM|Unspecified intellectual disabilities|Unspecified intellectual disabilities
C0085437|T047|HT|320|ICD9CM|Bacterial meningitis|Bacterial meningitis
C0178264|T047|HT|320-326.99|ICD9CM|INFLAMMATORY DISEASES OF THE CENTRAL NERVOUS SYSTEM|INFLAMMATORY DISEASES OF THE CENTRAL NERVOUS SYSTEM
C0338381|T047|HT|320-389.99|ICD9CM|DISEASES OF THE NERVOUS SYSTEM AND SENSE ORGANS|DISEASES OF THE NERVOUS SYSTEM AND SENSE ORGANS
C0025292|T047|AB|320.0|ICD9CM|Hemophilus meningitis|Hemophilus meningitis
C0025292|T047|PT|320.0|ICD9CM|Hemophilus meningitis|Hemophilus meningitis
C0025295|T047|AB|320.1|ICD9CM|Pneumococcal meningitis|Pneumococcal meningitis
C0025295|T047|PT|320.1|ICD9CM|Pneumococcal meningitis|Pneumococcal meningitis
C0154639|T047|AB|320.2|ICD9CM|Streptococcal meningitis|Streptococcal meningitis
C0154639|T047|PT|320.2|ICD9CM|Streptococcal meningitis|Streptococcal meningitis
C0154640|T047|AB|320.3|ICD9CM|Staphylococc meningitis|Staphylococc meningitis
C0154640|T047|PT|320.3|ICD9CM|Staphylococcal meningitis|Staphylococcal meningitis
C0154641|T047|AB|320.7|ICD9CM|Mening in oth bact dis|Mening in oth bact dis
C0154641|T047|PT|320.7|ICD9CM|Meningitis in other bacterial diseases classified elsewhere|Meningitis in other bacterial diseases classified elsewhere
C0154642|T047|HT|320.8|ICD9CM|Meningitis due to other specified bacteria|Meningitis due to other specified bacteria
C0375197|T047|AB|320.81|ICD9CM|Anaerobic meningitis|Anaerobic meningitis
C0375197|T047|PT|320.81|ICD9CM|Anaerobic meningitis|Anaerobic meningitis
C0375198|T047|PT|320.82|ICD9CM|Meningitis due to gram-negative bacteria, not elsewhere classified|Meningitis due to gram-negative bacteria, not elsewhere classified
C0375198|T047|AB|320.82|ICD9CM|Mningts gram-neg bct NEC|Mningts gram-neg bct NEC
C0154642|T047|PT|320.89|ICD9CM|Meningitis due to other specified bacteria|Meningitis due to other specified bacteria
C0154642|T047|AB|320.89|ICD9CM|Meningitis oth spcf bact|Meningitis oth spcf bact
C0085437|T047|AB|320.9|ICD9CM|Bacterial meningitis NOS|Bacterial meningitis NOS
C0085437|T047|PT|320.9|ICD9CM|Meningitis due to unspecified bacterium|Meningitis due to unspecified bacterium
C0154644|T047|HT|321|ICD9CM|Meningitis due to other organisms|Meningitis due to other organisms
C0085436|T047|AB|321.0|ICD9CM|Cryptococcal meningitis|Cryptococcal meningitis
C0085436|T047|PT|321.0|ICD9CM|Cryptococcal meningitis|Cryptococcal meningitis
C0154645|T047|AB|321.1|ICD9CM|Mening in oth fungal dis|Mening in oth fungal dis
C0154645|T047|PT|321.1|ICD9CM|Meningitis in other fungal diseases|Meningitis in other fungal diseases
C0868783|T047|AB|321.2|ICD9CM|Mening in oth viral dis|Mening in oth viral dis
C0868783|T047|PT|321.2|ICD9CM|Meningitis due to viruses not elsewhere classified|Meningitis due to viruses not elsewhere classified
C0795686|T047|PT|321.3|ICD9CM|Meningitis due to trypanosomiasis|Meningitis due to trypanosomiasis
C0795686|T047|AB|321.3|ICD9CM|Trypanosomiasis meningit|Trypanosomiasis meningit
C0154648|T047|AB|321.4|ICD9CM|Meningit d/t sarcoidosis|Meningit d/t sarcoidosis
C0154648|T047|PT|321.4|ICD9CM|Meningitis in sarcoidosis|Meningitis in sarcoidosis
C0154649|T047|AB|321.8|ICD9CM|Mening in oth nonbac dis|Mening in oth nonbac dis
C0154649|T047|PT|321.8|ICD9CM|Meningitis due to other nonbacterial organisms classified elsewhere|Meningitis due to other nonbacterial organisms classified elsewhere
C0025289|T047|HT|322|ICD9CM|Meningitis of unspecified cause|Meningitis of unspecified cause
C0154651|T047|AB|322.0|ICD9CM|Nonpyogenic meningitis|Nonpyogenic meningitis
C0154651|T047|PT|322.0|ICD9CM|Nonpyogenic meningitis|Nonpyogenic meningitis
C0154652|T047|AB|322.1|ICD9CM|Eosinophilic meningitis|Eosinophilic meningitis
C0154652|T047|PT|322.1|ICD9CM|Eosinophilic meningitis|Eosinophilic meningitis
C0154653|T047|AB|322.2|ICD9CM|Chronic meningitis|Chronic meningitis
C0154653|T047|PT|322.2|ICD9CM|Chronic meningitis|Chronic meningitis
C0025289|T047|AB|322.9|ICD9CM|Meningitis NOS|Meningitis NOS
C0025289|T047|PT|322.9|ICD9CM|Meningitis, unspecified|Meningitis, unspecified
C0014058|T047|HT|323|ICD9CM|Encephalitis, myelitis, and encephalomyelitis|Encephalitis, myelitis, and encephalomyelitis
C0477341|T047|HT|323.0|ICD9CM|Encephalitis, myelitis, and encephalomyelitis in viral diseases classified elsewhere|Encephalitis, myelitis, and encephalomyelitis in viral diseases classified elsewhere
C1719346|T047|AB|323.01|ICD9CM|Enceph/encephmye oth dis|Enceph/encephmye oth dis
C1719346|T047|PT|323.01|ICD9CM|Encephalitis and encephalomyelitis in viral diseases classified elsewhere|Encephalitis and encephalomyelitis in viral diseases classified elsewhere
C1719347|T047|PT|323.02|ICD9CM|Myelitis in viral diseases classified elsewhere|Myelitis in viral diseases classified elsewhere
C1719347|T047|AB|323.02|ICD9CM|Myelitis-oth viral dis|Myelitis-oth viral dis
C1719348|T047|PT|323.1|ICD9CM|Encephalitis, myelitis, and encephalomyelitis in rickettsial diseases classified elsewhere|Encephalitis, myelitis, and encephalomyelitis in rickettsial diseases classified elsewhere
C1719348|T047|AB|323.1|ICD9CM|Rickettsial encephalitis|Rickettsial encephalitis
C1719349|T047|PT|323.2|ICD9CM|Encephalitis, myelitis, and encephalomyelitis in protozoal diseases classified elsewhere|Encephalitis, myelitis, and encephalomyelitis in protozoal diseases classified elsewhere
C1719349|T047|AB|323.2|ICD9CM|Protozoal encephalitis|Protozoal encephalitis
C1719352|T047|HT|323.4|ICD9CM|Other encephalitis, myelitis, and encephalomyelitis due to other infections classified elsewhere|Other encephalitis, myelitis, and encephalomyelitis due to other infections classified elsewhere
C1719350|T047|AB|323.41|ICD9CM|Ot encph/mye ot inf else|Ot encph/mye ot inf else
C1719350|T047|PT|323.41|ICD9CM|Other encephalitis and encephalomyelitis due to other infections classified elsewhere|Other encephalitis and encephalomyelitis due to other infections classified elsewhere
C1719351|T047|AB|323.42|ICD9CM|Oth myelitis ot inf else|Oth myelitis ot inf else
C1719351|T047|PT|323.42|ICD9CM|Other myelitis due to other infections classified elsewhere|Other myelitis due to other infections classified elsewhere
C1719358|T046|HT|323.5|ICD9CM|Encephalitis, myelitis, and encephalomyelitis following immunization procedures|Encephalitis, myelitis, and encephalomyelitis following immunization procedures
C1719353|T046|AB|323.51|ICD9CM|Enceph/myel folwg immune|Enceph/myel folwg immune
C1719353|T046|PT|323.51|ICD9CM|Encephalitis and encephalomyelitis following immunization procedures|Encephalitis and encephalomyelitis following immunization procedures
C1997588|T047|PT|323.52|ICD9CM|Myelitis following immunization procedures|Myelitis following immunization procedures
C1997588|T047|AB|323.52|ICD9CM|Myelitis follwg immune|Myelitis follwg immune
C1719361|T047|HT|323.6|ICD9CM|Postinfectious encephalitis, myelitis, and encephalomyelitis|Postinfectious encephalitis, myelitis, and encephalomyelitis
C1719722|T047|AB|323.61|ICD9CM|Inf ac dis encephalomyel|Inf ac dis encephalomyel
C1719722|T047|PT|323.61|ICD9CM|Infectious acute disseminated encephalomyelitis (ADEM)|Infectious acute disseminated encephalomyelitis (ADEM)
C1719360|T047|PT|323.62|ICD9CM|Other postinfectious encephalitis and encephalomyelitis|Other postinfectious encephalitis and encephalomyelitis
C1719360|T047|AB|323.62|ICD9CM|Postinf encephalitis NEC|Postinf encephalitis NEC
C0751343|T047|AB|323.63|ICD9CM|Postinfectious myelitis|Postinfectious myelitis
C0751343|T047|PT|323.63|ICD9CM|Postinfectious myelitis|Postinfectious myelitis
C1719364|T037|HT|323.7|ICD9CM|Toxic encephalitis, myelitis, and encephalomyelitis|Toxic encephalitis, myelitis, and encephalomyelitis
C1719362|T047|PT|323.71|ICD9CM|Toxic encephalitis and encephalomyelitis|Toxic encephalitis and encephalomyelitis
C1719362|T047|AB|323.71|ICD9CM|Toxic encph & encephlomy|Toxic encph & encephlomy
C2316057|T047|PT|323.72|ICD9CM|Toxic myelitis|Toxic myelitis
C2316057|T047|AB|323.72|ICD9CM|Toxic myelitis|Toxic myelitis
C1719368|T047|HT|323.8|ICD9CM|Other causes of encephalitis, myelitis, and encephalomyelitis|Other causes of encephalitis, myelitis, and encephalomyelitis
C1719365|T047|AB|323.81|ICD9CM|Enceph & encephlalo NEC|Enceph & encephlalo NEC
C1719365|T047|PT|323.81|ICD9CM|Other causes of encephalitis and encephalomyelitis|Other causes of encephalitis and encephalomyelitis
C1719367|T047|AB|323.82|ICD9CM|Myelitis cause NEC|Myelitis cause NEC
C1719367|T047|PT|323.82|ICD9CM|Other causes of myelitis|Other causes of myelitis
C1719369|T033|AB|323.9|ICD9CM|Encephalitis NOS|Encephalitis NOS
C1719369|T033|PT|323.9|ICD9CM|Unspecified causes of encephalitis, myelitis, and encephalomyelitis|Unspecified causes of encephalitis, myelitis, and encephalomyelitis
C0154660|T047|HT|324|ICD9CM|Intracranial and intraspinal abscess|Intracranial and intraspinal abscess
C0021874|T047|AB|324.0|ICD9CM|Intracranial abscess|Intracranial abscess
C0021874|T047|PT|324.0|ICD9CM|Intracranial abscess|Intracranial abscess
C0154661|T020|AB|324.1|ICD9CM|Intraspinal abscess|Intraspinal abscess
C0154661|T020|PT|324.1|ICD9CM|Intraspinal abscess|Intraspinal abscess
C0154660|T047|AB|324.9|ICD9CM|Cns abscess NOS|Cns abscess NOS
C0154660|T047|PT|324.9|ICD9CM|Intracranial and intraspinal abscess of unspecified site|Intracranial and intraspinal abscess of unspecified site
C0154662|T047|PT|325|ICD9CM|Phlebitis and thrombophlebitis of intracranial venous sinuses|Phlebitis and thrombophlebitis of intracranial venous sinuses
C0154662|T047|AB|325|ICD9CM|Phlebitis intrcran sinus|Phlebitis intrcran sinus
C0154663|T047|AB|326|ICD9CM|Late eff cns abscess|Late eff cns abscess
C0154663|T047|PT|326|ICD9CM|Late effects of intracranial abscess or pyogenic infection|Late effects of intracranial abscess or pyogenic infection
C1561892|T047|HT|327|ICD9CM|Organic sleep disorders|Organic sleep disorders
C1561892|T047|HT|327-327.99|ICD9CM|ORGANIC SLEEP DISORDERS|ORGANIC SLEEP DISORDERS
C1561852|T047|HT|327.0|ICD9CM|Organic disorders of initiating and maintaining sleep [Organic insomnia]|Organic disorders of initiating and maintaining sleep [Organic insomnia]
C0021607|T048|AB|327.00|ICD9CM|Organic insomnia NOS|Organic insomnia NOS
C0021607|T048|PT|327.00|ICD9CM|Organic insomnia, unspecified|Organic insomnia, unspecified
C1561849|T047|PT|327.01|ICD9CM|Insomnia due to medical condition classified elsewhere|Insomnia due to medical condition classified elsewhere
C1561849|T047|AB|327.01|ICD9CM|Insomnia in other dis|Insomnia in other dis
C1561850|T048|AB|327.02|ICD9CM|Insomnia dt mental disor|Insomnia dt mental disor
C1561850|T048|PT|327.02|ICD9CM|Insomnia due to mental disorder|Insomnia due to mental disorder
C1561851|T047|AB|327.09|ICD9CM|Organic insomnia NEC|Organic insomnia NEC
C1561851|T047|PT|327.09|ICD9CM|Other organic insomnia|Other organic insomnia
C1561860|T047|HT|327.1|ICD9CM|Organic disorder of excessive somnolence [Organic hypersomnia]|Organic disorder of excessive somnolence [Organic hypersomnia]
C0270543|T047|AB|327.10|ICD9CM|Organic hypersomnia NOS|Organic hypersomnia NOS
C0270543|T047|PT|327.10|ICD9CM|Organic hypersomnia, unspecified|Organic hypersomnia, unspecified
C2711059|T047|AB|327.11|ICD9CM|Idio hypersom-long sleep|Idio hypersom-long sleep
C2711059|T047|PT|327.11|ICD9CM|Idiopathic hypersomnia with long sleep time|Idiopathic hypersomnia with long sleep time
C1561855|T047|AB|327.12|ICD9CM|Idio hypersom-no lng slp|Idio hypersom-no lng slp
C1561855|T047|PT|327.12|ICD9CM|Idiopathic hypersomnia without long sleep time|Idiopathic hypersomnia without long sleep time
C0751226|T047|AB|327.13|ICD9CM|Recurrent hypersomnia|Recurrent hypersomnia
C0751226|T047|PT|327.13|ICD9CM|Recurrent hypersomnia|Recurrent hypersomnia
C1561857|T047|PT|327.14|ICD9CM|Hypersomnia due to medical condition classified elsewhere|Hypersomnia due to medical condition classified elsewhere
C1561857|T047|AB|327.14|ICD9CM|Hypersomnia in other dis|Hypersomnia in other dis
C1561858|T048|AB|327.15|ICD9CM|Hypersom dt mental disor|Hypersom dt mental disor
C1561858|T048|PT|327.15|ICD9CM|Hypersomnia due to mental disorder|Hypersomnia due to mental disorder
C1561859|T047|AB|327.19|ICD9CM|Organic hypersomnia NEC|Organic hypersomnia NEC
C1561859|T047|PT|327.19|ICD9CM|Other organic hypersomnia|Other organic hypersomnia
C1561861|T047|HT|327.2|ICD9CM|Organic sleep apnea|Organic sleep apnea
C1561861|T047|AB|327.20|ICD9CM|Organic sleep apnea NOS|Organic sleep apnea NOS
C1561861|T047|PT|327.20|ICD9CM|Organic sleep apnea, unspecified|Organic sleep apnea, unspecified
C0751762|T047|AB|327.21|ICD9CM|Prim central sleep apnea|Prim central sleep apnea
C0751762|T047|PT|327.21|ICD9CM|Primary central sleep apnea|Primary central sleep apnea
C1561862|T047|AB|327.22|ICD9CM|High altitude breathing|High altitude breathing
C1561862|T047|PT|327.22|ICD9CM|High altitude periodic breathing|High altitude periodic breathing
C0520679|T047|AB|327.23|ICD9CM|Obstructive sleep apnea|Obstructive sleep apnea
C0520679|T047|PT|327.23|ICD9CM|Obstructive sleep apnea (adult)(pediatric)|Obstructive sleep apnea (adult)(pediatric)
C2711232|T047|AB|327.24|ICD9CM|Idiopath sleep hypovent|Idiopath sleep hypovent
C2711232|T047|PT|327.24|ICD9CM|Idiopathic sleep related non-obstructive alveolar hypoventilation|Idiopathic sleep related non-obstructive alveolar hypoventilation
C1561866|T047|AB|327.25|ICD9CM|Cong cntrl hypovent synd|Cong cntrl hypovent synd
C1561866|T047|PT|327.25|ICD9CM|Congenital central alveolar hypoventilation syndrome|Congenital central alveolar hypoventilation syndrome
C1561867|T047|AB|327.26|ICD9CM|Sleep hypovent oth dis|Sleep hypovent oth dis
C1561867|T047|PT|327.26|ICD9CM|Sleep related hypoventilation/hypoxemia in conditions classifiable elsewhere|Sleep related hypoventilation/hypoxemia in conditions classifiable elsewhere
C1561868|T047|PT|327.27|ICD9CM|Central sleep apnea in conditions classified elsewhere|Central sleep apnea in conditions classified elsewhere
C1561868|T047|AB|327.27|ICD9CM|Cntrl sleep apnea ot dis|Cntrl sleep apnea ot dis
C1561869|T047|AB|327.29|ICD9CM|Organic sleep apnea NEC|Organic sleep apnea NEC
C1561869|T047|PT|327.29|ICD9CM|Other organic sleep apnea|Other organic sleep apnea
C0877792|T046|HT|327.3|ICD9CM|Circadian rhythm sleep disorder|Circadian rhythm sleep disorder
C1561871|T047|AB|327.30|ICD9CM|Circadian rhym sleep NOS|Circadian rhym sleep NOS
C1561871|T047|PT|327.30|ICD9CM|Circadian rhythm sleep disorder, unspecified|Circadian rhythm sleep disorder, unspecified
C0393770|T047|AB|327.31|ICD9CM|Circadian rhy-delay slp|Circadian rhy-delay slp
C0393770|T047|PT|327.31|ICD9CM|Circadian rhythm sleep disorder, delayed sleep phase type|Circadian rhythm sleep disorder, delayed sleep phase type
C0751758|T047|AB|327.32|ICD9CM|Circadian rhy-advc sleep|Circadian rhy-advc sleep
C0751758|T047|PT|327.32|ICD9CM|Circadian rhythm sleep disorder, advanced sleep phase type|Circadian rhythm sleep disorder, advanced sleep phase type
C1561874|T047|AB|327.33|ICD9CM|Circadian rhym-irreg slp|Circadian rhym-irreg slp
C1561874|T047|PT|327.33|ICD9CM|Circadian rhythm sleep disorder, irregular sleep-wake type|Circadian rhythm sleep disorder, irregular sleep-wake type
C0393772|T033|AB|327.34|ICD9CM|Circadian rhym-free run|Circadian rhym-free run
C0393772|T033|PT|327.34|ICD9CM|Circadian rhythm sleep disorder, free-running type|Circadian rhythm sleep disorder, free-running type
C0231311|T047|PT|327.35|ICD9CM|Circadian rhythm sleep disorder, jet lag type|Circadian rhythm sleep disorder, jet lag type
C0231311|T047|AB|327.35|ICD9CM|Circadian rhythm-jetlag|Circadian rhythm-jetlag
C0393773|T047|AB|327.36|ICD9CM|Circadian rhy-shift work|Circadian rhy-shift work
C0393773|T047|PT|327.36|ICD9CM|Circadian rhythm sleep disorder, shift work type|Circadian rhythm sleep disorder, shift work type
C1561878|T047|AB|327.37|ICD9CM|Circadian rhym oth dis|Circadian rhym oth dis
C1561878|T047|PT|327.37|ICD9CM|Circadian rhythm sleep disorder in conditions classified elsewhere|Circadian rhythm sleep disorder in conditions classified elsewhere
C1561879|T047|AB|327.39|ICD9CM|Circadian rhym sleep NEC|Circadian rhym sleep NEC
C1561879|T047|PT|327.39|ICD9CM|Other circadian rhythm sleep disorder|Other circadian rhythm sleep disorder
C1561882|T047|HT|327.4|ICD9CM|Organic parasomnia|Organic parasomnia
C1561882|T047|AB|327.40|ICD9CM|Organic parasomnia NOS|Organic parasomnia NOS
C1561882|T047|PT|327.40|ICD9CM|Organic parasomnia, unspecified|Organic parasomnia, unspecified
C0752295|T048|AB|327.41|ICD9CM|Confusional arousals|Confusional arousals
C0752295|T048|PT|327.41|ICD9CM|Confusional arousals|Confusional arousals
C0751772|T048|AB|327.42|ICD9CM|REM sleep behavior dis|REM sleep behavior dis
C0751772|T048|PT|327.42|ICD9CM|REM sleep behavior disorder|REM sleep behavior disorder
C1561883|T046|PT|327.43|ICD9CM|Recurrent isolated sleep paralysis|Recurrent isolated sleep paralysis
C1561883|T046|AB|327.43|ICD9CM|Recurrnt sleep paralysis|Recurrnt sleep paralysis
C3693456|T047|PT|327.44|ICD9CM|Parasomnia in conditions classified elsewhere|Parasomnia in conditions classified elsewhere
C3693456|T047|AB|327.44|ICD9CM|Parasomnia oth diseases|Parasomnia oth diseases
C1561885|T047|AB|327.49|ICD9CM|Organic parasomnia NEC|Organic parasomnia NEC
C1561885|T047|PT|327.49|ICD9CM|Other organic parasomnia|Other organic parasomnia
C1561890|T047|HT|327.5|ICD9CM|Organic sleep related movement disorders|Organic sleep related movement disorders
C0751774|T047|AB|327.51|ICD9CM|Periodic limb movement|Periodic limb movement
C0751774|T047|PT|327.51|ICD9CM|Periodic limb movement disorder|Periodic limb movement disorder
C1561888|T047|AB|327.52|ICD9CM|Sleep related leg cramps|Sleep related leg cramps
C1561888|T047|PT|327.52|ICD9CM|Sleep related leg cramps|Sleep related leg cramps
C0393774|T047|AB|327.53|ICD9CM|Sleep related bruxism|Sleep related bruxism
C0393774|T047|PT|327.53|ICD9CM|Sleep related bruxism|Sleep related bruxism
C1561889|T047|AB|327.59|ICD9CM|Organic sleep movemt NEC|Organic sleep movemt NEC
C1561889|T047|PT|327.59|ICD9CM|Other organic sleep related movement disorders|Other organic sleep related movement disorders
C1561891|T047|PT|327.8|ICD9CM|Other organic sleep disorders|Other organic sleep disorders
C1561891|T047|AB|327.8|ICD9CM|Sleep organic disord NEC|Sleep organic disord NEC
C0154664|T047|HT|330|ICD9CM|Cerebral degenerations usually manifest in childhood|Cerebral degenerations usually manifest in childhood
C1444208|T047|HT|330-337.99|ICD9CM|HEREDITARY AND DEGENERATIVE DISEASES OF THE CENTRAL NERVOUS SYSTEM|HEREDITARY AND DEGENERATIVE DISEASES OF THE CENTRAL NERVOUS SYSTEM
C0023520|T047|AB|330.0|ICD9CM|Leukodystrophy|Leukodystrophy
C0023520|T047|PT|330.0|ICD9CM|Leukodystrophy|Leukodystrophy
C0007788|T047|AB|330.1|ICD9CM|Cerebral lipidoses|Cerebral lipidoses
C0007788|T047|PT|330.1|ICD9CM|Cerebral lipidoses|Cerebral lipidoses
C1689951|T047|AB|330.2|ICD9CM|Cereb degen in lipidosis|Cereb degen in lipidosis
C1689951|T047|PT|330.2|ICD9CM|Cerebral degeneration in generalized lipidoses|Cerebral degeneration in generalized lipidoses
C0154666|T047|AB|330.3|ICD9CM|Cerb deg chld in oth dis|Cerb deg chld in oth dis
C0154666|T047|PT|330.3|ICD9CM|Cerebral degeneration of childhood in other diseases classified elsewhere|Cerebral degeneration of childhood in other diseases classified elsewhere
C0029753|T047|AB|330.8|ICD9CM|Cereb degen in child NEC|Cereb degen in child NEC
C0029753|T047|PT|330.8|ICD9CM|Other specified cerebral degenerations in childhood|Other specified cerebral degenerations in childhood
C0154667|T047|AB|330.9|ICD9CM|Cereb degen in child NOS|Cereb degen in child NOS
C0154667|T047|PT|330.9|ICD9CM|Unspecified cerebral degeneration in childhood|Unspecified cerebral degeneration in childhood
C0154668|T047|HT|331|ICD9CM|Other cerebral degenerations|Other cerebral degenerations
C0002395|T047|AB|331.0|ICD9CM|Alzheimer's disease|Alzheimer's disease
C0002395|T047|PT|331.0|ICD9CM|Alzheimer's disease|Alzheimer's disease
C0338451|T047|HT|331.1|ICD9CM|Frontotemporal dementia|Frontotemporal dementia
C0236642|T047|AB|331.11|ICD9CM|Pick's disease|Pick's disease
C0236642|T047|PT|331.11|ICD9CM|Pick's disease|Pick's disease
C1260406|T047|AB|331.19|ICD9CM|Frontotemp dementia NEC|Frontotemp dementia NEC
C1260406|T047|PT|331.19|ICD9CM|Other frontotemporal dementia|Other frontotemporal dementia
C0154669|T047|AB|331.2|ICD9CM|Senile degenerat brain|Senile degenerat brain
C0154669|T047|PT|331.2|ICD9CM|Senile degeneration of brain|Senile degeneration of brain
C0009451|T047|AB|331.3|ICD9CM|Communicat hydrocephalus|Communicat hydrocephalus
C0009451|T047|PT|331.3|ICD9CM|Communicating hydrocephalus|Communicating hydrocephalus
C0549423|T047|AB|331.4|ICD9CM|Obstructiv hydrocephalus|Obstructiv hydrocephalus
C0549423|T047|PT|331.4|ICD9CM|Obstructive hydrocephalus|Obstructive hydrocephalus
C1955760|T047|PT|331.5|ICD9CM|Idiopathic normal pressure hydrocephalus (INPH)|Idiopathic normal pressure hydrocephalus (INPH)
C1955760|T047|AB|331.5|ICD9CM|Norml pressure hydroceph|Norml pressure hydroceph
C0393570|T047|PT|331.6|ICD9CM|Corticobasal degeneration|Corticobasal degeneration
C0393570|T047|AB|331.6|ICD9CM|Corticobasal degneration|Corticobasal degneration
C0393647|T047|AB|331.7|ICD9CM|Cereb degen in oth dis|Cereb degen in oth dis
C0393647|T047|PT|331.7|ICD9CM|Cerebral degeneration in diseases classified elsewhere|Cerebral degeneration in diseases classified elsewhere
C0154668|T047|HT|331.8|ICD9CM|Other cerebral degeneration|Other cerebral degeneration
C0035400|T047|AB|331.81|ICD9CM|Reye's syndrome|Reye's syndrome
C0035400|T047|PT|331.81|ICD9CM|Reye's syndrome|Reye's syndrome
C0752347|T047|AB|331.82|ICD9CM|Dementia w Lewy bodies|Dementia w Lewy bodies
C0752347|T047|PT|331.82|ICD9CM|Dementia with lewy bodies|Dementia with lewy bodies
C1719378|T047|AB|331.83|ICD9CM|Mild cognitive impairemt|Mild cognitive impairemt
C1719378|T047|PT|331.83|ICD9CM|Mild cognitive impairment, so stated|Mild cognitive impairment, so stated
C0154668|T047|AB|331.89|ICD9CM|Cereb degeneration NEC|Cereb degeneration NEC
C0154668|T047|PT|331.89|ICD9CM|Other cerebral degeneration|Other cerebral degeneration
C0154671|T047|AB|331.9|ICD9CM|Cereb degeneration NOS|Cereb degeneration NOS
C0154671|T047|PT|331.9|ICD9CM|Cerebral degeneration, unspecified|Cerebral degeneration, unspecified
C0030567|T047|HT|332|ICD9CM|Parkinson's disease|Parkinson's disease
C0030567|T047|AB|332.0|ICD9CM|Paralysis agitans|Paralysis agitans
C0030567|T047|PT|332.0|ICD9CM|Paralysis agitans|Paralysis agitans
C0030569|T047|AB|332.1|ICD9CM|Secondary parkinsonism|Secondary parkinsonism
C0030569|T047|PT|332.1|ICD9CM|Secondary parkinsonism|Secondary parkinsonism
C0154678|T047|HT|333|ICD9CM|Other extrapyramidal disease and abnormal movement disorders|Other extrapyramidal disease and abnormal movement disorders
C0029571|T047|AB|333.0|ICD9CM|Degen basal ganglia NEC|Degen basal ganglia NEC
C0029571|T047|PT|333.0|ICD9CM|Other degenerative diseases of the basal ganglia|Other degenerative diseases of the basal ganglia
C1961111|T184|PT|333.1|ICD9CM|Essential and other specified forms of tremor|Essential and other specified forms of tremor
C1961111|T184|AB|333.1|ICD9CM|Tremor NEC|Tremor NEC
C0027066|T184|AB|333.2|ICD9CM|Myoclonus|Myoclonus
C0027066|T184|PT|333.2|ICD9CM|Myoclonus|Myoclonus
C0702141|T046|AB|333.3|ICD9CM|Tics of organic origin|Tics of organic origin
C0702141|T046|PT|333.3|ICD9CM|Tics of organic origin|Tics of organic origin
C0020179|T047|AB|333.4|ICD9CM|Huntington's chorea|Huntington's chorea
C0020179|T047|PT|333.4|ICD9CM|Huntington's chorea|Huntington's chorea
C0029542|T046|AB|333.5|ICD9CM|Chorea NEC|Chorea NEC
C0029542|T046|PT|333.5|ICD9CM|Other choreas|Other choreas
C0013423|T047|PT|333.6|ICD9CM|Genetic torsion dystonia|Genetic torsion dystonia
C0013423|T047|AB|333.6|ICD9CM|Genetic torsion dystonia|Genetic torsion dystonia
C1719382|T047|HT|333.7|ICD9CM|Acquired torsion dystonia|Acquired torsion dystonia
C0270742|T047|PT|333.71|ICD9CM|Athetoid cerebral palsy|Athetoid cerebral palsy
C0270742|T047|AB|333.71|ICD9CM|Athetoid cerebral palsy|Athetoid cerebral palsy
C0393596|T046|AB|333.72|ICD9CM|Acute dystonia d/t drugs|Acute dystonia d/t drugs
C0393596|T046|PT|333.72|ICD9CM|Acute dystonia due to drugs|Acute dystonia due to drugs
C1719381|T047|AB|333.79|ICD9CM|Acq torsion dystonia NEC|Acq torsion dystonia NEC
C1719381|T047|PT|333.79|ICD9CM|Other acquired torsion dystonia|Other acquired torsion dystonia
C0154675|T047|HT|333.8|ICD9CM|Fragments of torsion dystonia|Fragments of torsion dystonia
C0005747|T047|AB|333.81|ICD9CM|Blepharospasm|Blepharospasm
C0005747|T047|PT|333.81|ICD9CM|Blepharospasm|Blepharospasm
C0152115|T047|AB|333.82|ICD9CM|Orofacial dyskinesia|Orofacial dyskinesia
C0152115|T047|PT|333.82|ICD9CM|Orofacial dyskinesia|Orofacial dyskinesia
C0152116|T184|AB|333.83|ICD9CM|Spasmodic torticollis|Spasmodic torticollis
C0152116|T184|PT|333.83|ICD9CM|Spasmodic torticollis|Spasmodic torticollis
C0154676|T047|AB|333.84|ICD9CM|Organic writers' cramp|Organic writers' cramp
C0154676|T047|PT|333.84|ICD9CM|Organic writers' cramp|Organic writers' cramp
C3662039|T047|AB|333.85|ICD9CM|Subac dyskinesa d/t drug|Subac dyskinesa d/t drug
C3662039|T047|PT|333.85|ICD9CM|Subacute dyskinesia due to drugs|Subacute dyskinesia due to drugs
C0154677|T047|AB|333.89|ICD9CM|Fragm torsion dyston NEC|Fragm torsion dyston NEC
C0154677|T047|PT|333.89|ICD9CM|Other fragments of torsion dystonia|Other fragments of torsion dystonia
C0154678|T047|HT|333.9|ICD9CM|Other and unspecified extrapyramidal diseases and abnormal movement disorders|Other and unspecified extrapyramidal diseases and abnormal movement disorders
C0477355|T047|AB|333.90|ICD9CM|Extrapyramidal dis NOS|Extrapyramidal dis NOS
C0477355|T047|PT|333.90|ICD9CM|Unspecified extrapyramidal disease and abnormal movement disorder|Unspecified extrapyramidal disease and abnormal movement disorder
C0085292|T047|AB|333.91|ICD9CM|Stiff-man syndrome|Stiff-man syndrome
C0085292|T047|PT|333.91|ICD9CM|Stiff-man syndrome|Stiff-man syndrome
C0027849|T047|AB|333.92|ICD9CM|Neuroleptic malgnt synd|Neuroleptic malgnt synd
C0027849|T047|PT|333.92|ICD9CM|Neuroleptic malignant syndrome|Neuroleptic malignant syndrome
C0375200|T047|PT|333.93|ICD9CM|Benign shuddering attacks|Benign shuddering attacks
C0375200|T047|AB|333.93|ICD9CM|Bnign shuddering attacks|Bnign shuddering attacks
C0035258|T047|AB|333.94|ICD9CM|Restless legs syndrome|Restless legs syndrome
C0035258|T047|PT|333.94|ICD9CM|Restless legs syndrome (RLS)|Restless legs syndrome (RLS)
C0154678|T047|AB|333.99|ICD9CM|Extrapyramidal dis NEC|Extrapyramidal dis NEC
C0154678|T047|PT|333.99|ICD9CM|Other extrapyramidal diseases and abnormal movement disorders|Other extrapyramidal diseases and abnormal movement disorders
C0037952|T047|HT|334|ICD9CM|Spinocerebellar disease|Spinocerebellar disease
C0016719|T047|AB|334.0|ICD9CM|Friedreich's ataxia|Friedreich's ataxia
C0016719|T047|PT|334.0|ICD9CM|Friedreich's ataxia|Friedreich's ataxia
C0037773|T047|AB|334.1|ICD9CM|Hered spastic paraplegia|Hered spastic paraplegia
C0037773|T047|PT|334.1|ICD9CM|Hereditary spastic paraplegia|Hereditary spastic paraplegia
C0033132|T047|AB|334.2|ICD9CM|Primary cerebellar degen|Primary cerebellar degen
C0033132|T047|PT|334.2|ICD9CM|Primary cerebellar degeneration|Primary cerebellar degeneration
C0029534|T047|AB|334.3|ICD9CM|Cerebellar ataxia NEC|Cerebellar ataxia NEC
C0029534|T047|PT|334.3|ICD9CM|Other cerebellar ataxia|Other cerebellar ataxia
C0393517|T047|AB|334.4|ICD9CM|Cerebel atax in oth dis|Cerebel atax in oth dis
C0393517|T047|PT|334.4|ICD9CM|Cerebellar ataxia in diseases classified elsewhere|Cerebellar ataxia in diseases classified elsewhere
C0029849|T047|PT|334.8|ICD9CM|Other spinocerebellar diseases|Other spinocerebellar diseases
C0029849|T047|AB|334.8|ICD9CM|Spinocerebellar dis NEC|Spinocerebellar dis NEC
C0037952|T047|AB|334.9|ICD9CM|Spinocerebellar dis NOS|Spinocerebellar dis NOS
C0037952|T047|PT|334.9|ICD9CM|Spinocerebellar disease, unspecified|Spinocerebellar disease, unspecified
C0154681|T047|HT|335|ICD9CM|Anterior horn cell disease|Anterior horn cell disease
C0043116|T047|PT|335.0|ICD9CM|Werdnig-Hoffmann disease|Werdnig-Hoffmann disease
C0043116|T047|AB|335.0|ICD9CM|Werdnig-hoffmann disease|Werdnig-hoffmann disease
C0026847|T047|HT|335.1|ICD9CM|Spinal muscular atrophy|Spinal muscular atrophy
C0026847|T047|AB|335.10|ICD9CM|Spinal muscl atrophy NOS|Spinal muscl atrophy NOS
C0026847|T047|PT|335.10|ICD9CM|Spinal muscular atrophy, unspecified|Spinal muscular atrophy, unspecified
C0152109|T047|AB|335.11|ICD9CM|Kugelberg-welander dis|Kugelberg-welander dis
C0152109|T047|PT|335.11|ICD9CM|Kugelberg-Welander disease|Kugelberg-Welander disease
C0029848|T047|PT|335.19|ICD9CM|Other spinal muscular atrophy|Other spinal muscular atrophy
C0029848|T047|AB|335.19|ICD9CM|Spinal muscl atrophy NEC|Spinal muscl atrophy NEC
C0085084|T047|HT|335.2|ICD9CM|Motor neuron disease|Motor neuron disease
C0002736|T047|PT|335.20|ICD9CM|Amyotrophic lateral sclerosis|Amyotrophic lateral sclerosis
C0002736|T047|AB|335.20|ICD9CM|Amyotrophic sclerosis|Amyotrophic sclerosis
C0917981|T047|AB|335.21|ICD9CM|Prog muscular atrophy|Prog muscular atrophy
C0917981|T047|PT|335.21|ICD9CM|Progressive muscular atrophy|Progressive muscular atrophy
C0030442|T047|AB|335.22|ICD9CM|Progressive bulbar palsy|Progressive bulbar palsy
C0030442|T047|PT|335.22|ICD9CM|Progressive bulbar palsy|Progressive bulbar palsy
C0033790|T047|AB|335.23|ICD9CM|Pseudobulbar palsy|Pseudobulbar palsy
C0033790|T047|PT|335.23|ICD9CM|Pseudobulbar palsy|Pseudobulbar palsy
C0154682|T047|AB|335.24|ICD9CM|Prim lateral sclerosis|Prim lateral sclerosis
C0154682|T047|PT|335.24|ICD9CM|Primary lateral sclerosis|Primary lateral sclerosis
C0154683|T047|AB|335.29|ICD9CM|Motor neuron disease NEC|Motor neuron disease NEC
C0154683|T047|PT|335.29|ICD9CM|Other motor neuron disease|Other motor neuron disease
C0154684|T047|AB|335.8|ICD9CM|Ant horn cell dis NEC|Ant horn cell dis NEC
C0154684|T047|PT|335.8|ICD9CM|Other anterior horn cell diseases|Other anterior horn cell diseases
C0154681|T047|AB|335.9|ICD9CM|Ant horn cell dis NOS|Ant horn cell dis NOS
C0154681|T047|PT|335.9|ICD9CM|Anterior horn cell disease, unspecified|Anterior horn cell disease, unspecified
C0154688|T047|HT|336|ICD9CM|Other diseases of spinal cord|Other diseases of spinal cord
C0039145|T047|AB|336.0|ICD9CM|Syringomyelia|Syringomyelia
C0039145|T047|PT|336.0|ICD9CM|Syringomyelia and syringobulbia|Syringomyelia and syringobulbia
C0154685|T047|AB|336.1|ICD9CM|Vascular myelopathies|Vascular myelopathies
C0154685|T047|PT|336.1|ICD9CM|Vascular myelopathies|Vascular myelopathies
C0154686|T047|AB|336.2|ICD9CM|Comb deg cord in oth dis|Comb deg cord in oth dis
C0154686|T047|PT|336.2|ICD9CM|Subacute combined degeneration of spinal cord in diseases classified elsewhere|Subacute combined degeneration of spinal cord in diseases classified elsewhere
C0154687|T047|AB|336.3|ICD9CM|Myelopathy in oth dis|Myelopathy in oth dis
C0154687|T047|PT|336.3|ICD9CM|Myelopathy in other diseases classified elsewhere|Myelopathy in other diseases classified elsewhere
C1961841|T047|AB|336.8|ICD9CM|Myelopathy NEC|Myelopathy NEC
C1961841|T047|PT|336.8|ICD9CM|Other myelopathy|Other myelopathy
C0037928|T047|AB|336.9|ICD9CM|Spinal cord disease NOS|Spinal cord disease NOS
C0037928|T047|PT|336.9|ICD9CM|Unspecified disease of spinal cord|Unspecified disease of spinal cord
C1145628|T047|HT|337|ICD9CM|Disorders of the autonomic nervous system|Disorders of the autonomic nervous system
C0154690|T047|HT|337.0|ICD9CM|Idiopathic peripheral autonomic neuropathy|Idiopathic peripheral autonomic neuropathy
C2349410|T047|AB|337.00|ICD9CM|Idio perph auto neur NOS|Idio perph auto neur NOS
C2349410|T047|PT|337.00|ICD9CM|Idiopathic peripheral autonomic neuropathy, unspecified|Idiopathic peripheral autonomic neuropathy, unspecified
C0221046|T047|PT|337.01|ICD9CM|Carotid sinus syndrome|Carotid sinus syndrome
C0221046|T047|AB|337.01|ICD9CM|Carotid sinus syndrome|Carotid sinus syndrome
C2349411|T047|AB|337.09|ICD9CM|Idio perph auto neur NEC|Idio perph auto neur NEC
C2349411|T047|PT|337.09|ICD9CM|Other idiopathic peripheral autonomic neuropathy|Other idiopathic peripheral autonomic neuropathy
C0154691|T047|AB|337.1|ICD9CM|Aut neuropthy in oth dis|Aut neuropthy in oth dis
C0154691|T047|PT|337.1|ICD9CM|Peripheral autonomic neuropathy in disorders classified elsewhere|Peripheral autonomic neuropathy in disorders classified elsewhere
C0034931|T047|HT|337.2|ICD9CM|Reflex sympathetic dystrophy|Reflex sympathetic dystrophy
C0034931|T047|PT|337.20|ICD9CM|Reflex sympathetic dystrophy, unspecified|Reflex sympathetic dystrophy, unspecified
C0034931|T047|AB|337.20|ICD9CM|Unsp rflx sympth dystrph|Unsp rflx sympth dystrph
C4040007|T047|PT|337.21|ICD9CM|Reflex sympathetic dystrophy of the upper limb|Reflex sympathetic dystrophy of the upper limb
C4040007|T047|AB|337.21|ICD9CM|Rflx sym dystrph up limb|Rflx sym dystrph up limb
C0745890|T047|PT|337.22|ICD9CM|Reflex sympathetic dystrophy of the lower limb|Reflex sympathetic dystrophy of the lower limb
C0745890|T047|AB|337.22|ICD9CM|Rflx sym dystrph lwr lmb|Rflx sym dystrph lwr lmb
C0375204|T047|PT|337.29|ICD9CM|Reflex sympathetic dystrophy of other specified site|Reflex sympathetic dystrophy of other specified site
C0375204|T047|AB|337.29|ICD9CM|Rflx sym dystrph oth st|Rflx sym dystrph oth st
C0238015|T047|AB|337.3|ICD9CM|Autonomic dysreflexia|Autonomic dysreflexia
C0238015|T047|PT|337.3|ICD9CM|Autonomic dysreflexia|Autonomic dysreflexia
C1145628|T047|AB|337.9|ICD9CM|Autonomic nerve dis NEC|Autonomic nerve dis NEC
C1145628|T047|PT|337.9|ICD9CM|Unspecified disorder of autonomic nervous system|Unspecified disorder of autonomic nervous system
C0995154|T184|HT|338|ICD9CM|Pain, not elsewhere classified|Pain, not elsewhere classified
C0030193|T184|HT|338-338.99|ICD9CM|PAIN|PAIN
C1536114|T047|PT|338.0|ICD9CM|Central pain syndrome|Central pain syndrome
C1536114|T047|AB|338.0|ICD9CM|Central pain syndrome|Central pain syndrome
C0184567|T184|HT|338.1|ICD9CM|Acute pain|Acute pain
C1719389|T047|PT|338.11|ICD9CM|Acute pain due to trauma|Acute pain due to trauma
C1719389|T047|AB|338.11|ICD9CM|Acute pain due to trauma|Acute pain due to trauma
C1719390|T047|AB|338.12|ICD9CM|Acute post-thoracot pain|Acute post-thoracot pain
C1719390|T047|PT|338.12|ICD9CM|Acute post-thoracotomy pain|Acute post-thoracotomy pain
C1719392|T047|AB|338.18|ICD9CM|Acute postop pain NEC|Acute postop pain NEC
C1719392|T047|PT|338.18|ICD9CM|Other acute postoperative pain|Other acute postoperative pain
C1719723|T047|AB|338.19|ICD9CM|Acute pain NEC|Acute pain NEC
C1719723|T047|PT|338.19|ICD9CM|Other acute pain|Other acute pain
C0150055|T184|HT|338.2|ICD9CM|Chronic pain|Chronic pain
C1719393|T047|AB|338.21|ICD9CM|Chronc pain d/t trauma|Chronc pain d/t trauma
C1719393|T047|PT|338.21|ICD9CM|Chronic pain due to trauma|Chronic pain due to trauma
C1719710|T047|AB|338.22|ICD9CM|Chron post-thoracot pain|Chron post-thoracot pain
C1719710|T047|PT|338.22|ICD9CM|Chronic post-thoracotomy pain|Chronic post-thoracotomy pain
C1719394|T047|AB|338.28|ICD9CM|Chronic postop pain NEC|Chronic postop pain NEC
C1719394|T047|PT|338.28|ICD9CM|Other chronic postoperative pain|Other chronic postoperative pain
C0478148|T184|AB|338.29|ICD9CM|Chronic pain NEC|Chronic pain NEC
C0478148|T184|PT|338.29|ICD9CM|Other chronic pain|Other chronic pain
C1719395|T047|AB|338.3|ICD9CM|Neoplasm related pain|Neoplasm related pain
C1719395|T047|PT|338.3|ICD9CM|Neoplasm related pain (acute) (chronic)|Neoplasm related pain (acute) (chronic)
C1298685|T047|PT|338.4|ICD9CM|Chronic pain syndrome|Chronic pain syndrome
C1298685|T047|AB|338.4|ICD9CM|Chronic pain syndrome|Chronic pain syndrome
C0494479|T047|HT|339|ICD9CM|Other headache syndromes|Other headache syndromes
C0494479|T047|HT|339-339.99|ICD9CM|OTHER HEADACHE SYNDROMES|OTHER HEADACHE SYNDROMES
C2349419|T047|HT|339.0|ICD9CM|Cluster headaches and other trigeminal autonomic cephalgias|Cluster headaches and other trigeminal autonomic cephalgias
C0009088|T047|AB|339.00|ICD9CM|Cluster headache syn NOS|Cluster headache syn NOS
C0009088|T047|PT|339.00|ICD9CM|Cluster headache syndrome, unspecified|Cluster headache syndrome, unspecified
C0393739|T047|AB|339.01|ICD9CM|Episodc cluster headache|Episodc cluster headache
C0393739|T047|PT|339.01|ICD9CM|Episodic cluster headache|Episodic cluster headache
C0009088|T047|PT|339.02|ICD9CM|Chronic cluster headache|Chronic cluster headache
C0009088|T047|AB|339.02|ICD9CM|Chronic cluster headache|Chronic cluster headache
C1565171|T047|AB|339.03|ICD9CM|Episdc paroxyml hemicran|Episdc paroxyml hemicran
C1565171|T047|PT|339.03|ICD9CM|Episodic paroxysmal hemicrania|Episodic paroxysmal hemicrania
C0393743|T047|AB|339.04|ICD9CM|Chr paroxysml hemicrania|Chr paroxysml hemicrania
C0393743|T047|PT|339.04|ICD9CM|Chronic paroxysmal hemicrania|Chronic paroxysmal hemicrania
C2349417|T047|PT|339.05|ICD9CM|Short lasting unilateral neuralgiform headache with conjunctival injection and tearing|Short lasting unilateral neuralgiform headache with conjunctival injection and tearing
C2349417|T047|AB|339.05|ICD9CM|Shrt lst uni nral hdache|Shrt lst uni nral hdache
C2349418|T047|PT|339.09|ICD9CM|Other trigeminal autonomic cephalgias|Other trigeminal autonomic cephalgias
C2349418|T047|AB|339.09|ICD9CM|Trigem autonmc cephl NEC|Trigem autonmc cephl NEC
C0033893|T047|HT|339.1|ICD9CM|Tension type headache|Tension type headache
C0033893|T047|AB|339.10|ICD9CM|Tension headache NOS|Tension headache NOS
C0033893|T047|PT|339.10|ICD9CM|Tension type headache, unspecified|Tension type headache, unspecified
C0393737|T047|AB|339.11|ICD9CM|Episdic tension headache|Episdic tension headache
C0393737|T047|PT|339.11|ICD9CM|Episodic tension type headache|Episodic tension type headache
C0393738|T047|AB|339.12|ICD9CM|Chronic tension headache|Chronic tension headache
C0393738|T047|PT|339.12|ICD9CM|Chronic tension type headache|Chronic tension type headache
C0032816|T046|HT|339.2|ICD9CM|Post-traumatic headache|Post-traumatic headache
C0032816|T046|AB|339.20|ICD9CM|Post-trauma headache NOS|Post-trauma headache NOS
C0032816|T046|PT|339.20|ICD9CM|Post-traumatic headache, unspecified|Post-traumatic headache, unspecified
C2349421|T047|AB|339.21|ICD9CM|Ac post-trauma headache|Ac post-trauma headache
C2349421|T047|PT|339.21|ICD9CM|Acute post-traumatic headache|Acute post-traumatic headache
C0393745|T047|AB|339.22|ICD9CM|Chr post-trauma headache|Chr post-trauma headache
C0393745|T047|PT|339.22|ICD9CM|Chronic post-traumatic headache|Chronic post-traumatic headache
C2349422|T047|AB|339.3|ICD9CM|Drug induce headache NEC|Drug induce headache NEC
C2349422|T047|PT|339.3|ICD9CM|Drug induced headache, not elsewhere classified|Drug induced headache, not elsewhere classified
C2349428|T047|HT|339.4|ICD9CM|Complicated headache syndromes|Complicated headache syndromes
C2349425|T047|PT|339.41|ICD9CM|Hemicrania continua|Hemicrania continua
C2349425|T047|AB|339.41|ICD9CM|Hemicrania continua|Hemicrania continua
C2349426|T047|AB|339.42|ICD9CM|New daily pers headache|New daily pers headache
C2349426|T047|PT|339.42|ICD9CM|New daily persistent headache|New daily persistent headache
C0521668|T047|AB|339.43|ICD9CM|Prim thnderclap headache|Prim thnderclap headache
C0521668|T047|PT|339.43|ICD9CM|Primary thunderclap headache|Primary thunderclap headache
C2349427|T047|AB|339.44|ICD9CM|Comp headache synd NEC|Comp headache synd NEC
C2349427|T047|PT|339.44|ICD9CM|Other complicated headache syndrome|Other complicated headache syndrome
C0477374|T047|HT|339.8|ICD9CM|Other specified headache syndromes|Other specified headache syndromes
C0752150|T047|PT|339.81|ICD9CM|Hypnic headache|Hypnic headache
C0752150|T047|AB|339.81|ICD9CM|Hypnic headache|Hypnic headache
C0393754|T184|PT|339.82|ICD9CM|Headache associated with sexual activity|Headache associated with sexual activity
C0393754|T184|AB|339.82|ICD9CM|Headache w sex activity|Headache w sex activity
C0751185|T047|PT|339.83|ICD9CM|Primary cough headache|Primary cough headache
C0751185|T047|AB|339.83|ICD9CM|Primary cough headache|Primary cough headache
C0522253|T047|AB|339.84|ICD9CM|Prim exertion headache|Prim exertion headache
C0522253|T047|PT|339.84|ICD9CM|Primary exertional headache|Primary exertional headache
C0751191|T033|AB|339.85|ICD9CM|Prim stabbing headache|Prim stabbing headache
C0751191|T033|PT|339.85|ICD9CM|Primary stabbing headache|Primary stabbing headache
C0494479|T047|AB|339.89|ICD9CM|Headache syndrome NEC|Headache syndrome NEC
C0494479|T047|PT|339.89|ICD9CM|Other headache syndromes|Other headache syndromes
C0026769|T047|AB|340|ICD9CM|Multiple sclerosis|Multiple sclerosis
C0026769|T047|PT|340|ICD9CM|Multiple sclerosis|Multiple sclerosis
C0178266|T047|HT|340-349.99|ICD9CM|OTHER DISORDERS OF THE CENTRAL NERVOUS SYSTEM|OTHER DISORDERS OF THE CENTRAL NERVOUS SYSTEM
C0154692|T047|HT|341|ICD9CM|Other demyelinating diseases of central nervous system|Other demyelinating diseases of central nervous system
C0027873|T047|AB|341.0|ICD9CM|Neuromyelitis optica|Neuromyelitis optica
C0027873|T047|PT|341.0|ICD9CM|Neuromyelitis optica|Neuromyelitis optica
C0007795|T047|AB|341.1|ICD9CM|Schilder's disease|Schilder's disease
C0007795|T047|PT|341.1|ICD9CM|Schilder's disease|Schilder's disease
C0270627|T047|HT|341.2|ICD9CM|Acute (transverse) myelitis|Acute (transverse) myelitis
C0270627|T047|PT|341.20|ICD9CM|Acute (transverse) myelitis NOS|Acute (transverse) myelitis NOS
C0270627|T047|AB|341.20|ICD9CM|Acute myelitis NOS|Acute myelitis NOS
C1719403|T047|PT|341.21|ICD9CM|Acute (transverse) myelitis in conditions classified elsewhere|Acute (transverse) myelitis in conditions classified elsewhere
C1719403|T047|AB|341.21|ICD9CM|Acute myelitis oth cond|Acute myelitis oth cond
C1719404|T047|AB|341.22|ICD9CM|Idiopathc trans myelitis|Idiopathc trans myelitis
C1719404|T047|PT|341.22|ICD9CM|Idiopathic transverse myelitis|Idiopathic transverse myelitis
C0154692|T047|AB|341.8|ICD9CM|Cns demyelination NEC|Cns demyelination NEC
C0154692|T047|PT|341.8|ICD9CM|Other demyelinating diseases of central nervous system|Other demyelinating diseases of central nervous system
C0011302|T047|AB|341.9|ICD9CM|Cns demyelination NOS|Cns demyelination NOS
C0011302|T047|PT|341.9|ICD9CM|Demyelinating disease of central nervous system, unspecified|Demyelinating disease of central nervous system, unspecified
C0375206|T047|HT|342|ICD9CM|Hemiplegia and hemiparesis|Hemiplegia and hemiparesis
C0154693|T184|HT|342.0|ICD9CM|Flaccid hemiplegia|Flaccid hemiplegia
C0154693|T184|PT|342.00|ICD9CM|Flaccid hemiplegia and hemiparesis affecting unspecified side|Flaccid hemiplegia and hemiparesis affecting unspecified side
C0154693|T184|AB|342.00|ICD9CM|Flccd hmiplga unspf side|Flccd hmiplga unspf side
C0375208|T184|PT|342.01|ICD9CM|Flaccid hemiplegia and hemiparesis affecting dominant side|Flaccid hemiplegia and hemiparesis affecting dominant side
C0375208|T184|AB|342.01|ICD9CM|Flccd hmiplga domnt side|Flccd hmiplga domnt side
C0375209|T184|PT|342.02|ICD9CM|Flaccid hemiplegia and hemiparesis affecting nondominant side|Flaccid hemiplegia and hemiparesis affecting nondominant side
C0375209|T184|AB|342.02|ICD9CM|Flccd hmiplg nondmnt sde|Flccd hmiplg nondmnt sde
C0154694|T047|HT|342.1|ICD9CM|Spastic hemiplegia|Spastic hemiplegia
C0154694|T047|PT|342.10|ICD9CM|Spastic hemiplegia and hemiparesis affecting unspecified side|Spastic hemiplegia and hemiparesis affecting unspecified side
C0154694|T047|AB|342.10|ICD9CM|Spstc hmiplga unspf side|Spstc hmiplga unspf side
C0375211|T184|PT|342.11|ICD9CM|Spastic hemiplegia and hemiparesis affecting dominant side|Spastic hemiplegia and hemiparesis affecting dominant side
C0375211|T184|AB|342.11|ICD9CM|Spstc hmiplga domnt side|Spstc hmiplga domnt side
C0375212|T184|PT|342.12|ICD9CM|Spastic hemiplegia and hemiparesis affecting nondominant side|Spastic hemiplegia and hemiparesis affecting nondominant side
C0375212|T184|AB|342.12|ICD9CM|Spstc hmiplg nondmnt sde|Spstc hmiplg nondmnt sde
C0375213|T184|HT|342.8|ICD9CM|Other specified hemiplegia|Other specified hemiplegia
C0375214|T184|AB|342.80|ICD9CM|Ot sp hmiplga unspf side|Ot sp hmiplga unspf side
C0375214|T184|PT|342.80|ICD9CM|Other specified hemiplegia and hemiparesis affecting unspecified side|Other specified hemiplegia and hemiparesis affecting unspecified side
C0375215|T184|AB|342.81|ICD9CM|Ot sp hmiplga domnt side|Ot sp hmiplga domnt side
C0375215|T184|PT|342.81|ICD9CM|Other specified hemiplegia and hemiparesis affecting dominant side|Other specified hemiplegia and hemiparesis affecting dominant side
C0375216|T184|AB|342.82|ICD9CM|Ot sp hmiplg nondmnt sde|Ot sp hmiplg nondmnt sde
C0375216|T184|PT|342.82|ICD9CM|Other specified hemiplegia and hemiparesis affecting nondominant side|Other specified hemiplegia and hemiparesis affecting nondominant side
C0018991|T184|HT|342.9|ICD9CM|Hemiplegia, unspecified|Hemiplegia, unspecified
C0375218|T184|PT|342.90|ICD9CM|Hemiplegia, unspecified, affecting unspecified side|Hemiplegia, unspecified, affecting unspecified side
C0375218|T184|AB|342.90|ICD9CM|Unsp hemiplga unspf side|Unsp hemiplga unspf side
C0375219|T184|PT|342.91|ICD9CM|Hemiplegia, unspecified, affecting dominant side|Hemiplegia, unspecified, affecting dominant side
C0375219|T184|AB|342.91|ICD9CM|Unsp hemiplga domnt side|Unsp hemiplga domnt side
C0375220|T184|PT|342.92|ICD9CM|Hemiplegia, unspecified, affecting nondominant side|Hemiplegia, unspecified, affecting nondominant side
C0375220|T184|AB|342.92|ICD9CM|Unsp hmiplga nondmnt sde|Unsp hmiplga nondmnt sde
C0392549|T047|HT|343|ICD9CM|Infantile cerebral palsy|Infantile cerebral palsy
C0154695|T047|AB|343.0|ICD9CM|Congenital diplegia|Congenital diplegia
C0154695|T047|PT|343.0|ICD9CM|Congenital diplegia|Congenital diplegia
C0270805|T019|AB|343.1|ICD9CM|Congenital hemiplegia|Congenital hemiplegia
C0270805|T047|AB|343.1|ICD9CM|Congenital hemiplegia|Congenital hemiplegia
C0270805|T019|PT|343.1|ICD9CM|Congenital hemiplegia|Congenital hemiplegia
C0270805|T047|PT|343.1|ICD9CM|Congenital hemiplegia|Congenital hemiplegia
C0154697|T019|AB|343.2|ICD9CM|Congenital quadriplegia|Congenital quadriplegia
C0154697|T047|AB|343.2|ICD9CM|Congenital quadriplegia|Congenital quadriplegia
C0154697|T019|PT|343.2|ICD9CM|Congenital quadriplegia|Congenital quadriplegia
C0154697|T047|PT|343.2|ICD9CM|Congenital quadriplegia|Congenital quadriplegia
C0154698|T047|AB|343.3|ICD9CM|Congenital monoplegia|Congenital monoplegia
C0154698|T047|PT|343.3|ICD9CM|Congenital monoplegia|Congenital monoplegia
C0392550|T047|AB|343.4|ICD9CM|Infantile hemiplegia|Infantile hemiplegia
C0392550|T047|PT|343.4|ICD9CM|Infantile hemiplegia|Infantile hemiplegia
C0029806|T047|AB|343.8|ICD9CM|Cerebral palsy NEC|Cerebral palsy NEC
C0029806|T047|PT|343.8|ICD9CM|Other specified infantile cerebral palsy|Other specified infantile cerebral palsy
C0392549|T047|AB|343.9|ICD9CM|Cerebral palsy NOS|Cerebral palsy NOS
C0392549|T047|PT|343.9|ICD9CM|Infantile cerebral palsy, unspecified|Infantile cerebral palsy, unspecified
C0154700|T047|HT|344|ICD9CM|Other paralytic syndromes|Other paralytic syndromes
C0375221|T047|HT|344.0|ICD9CM|Quadriplegia and quadriparesis|Quadriplegia and quadriparesis
C0034372|T047|AB|344.00|ICD9CM|Quadriplegia, unspecifd|Quadriplegia, unspecifd
C0034372|T047|PT|344.00|ICD9CM|Quadriplegia, unspecified|Quadriplegia, unspecified
C0376129|T047|PT|344.01|ICD9CM|Quadriplegia, C1-C4, complete|Quadriplegia, C1-C4, complete
C0376129|T047|AB|344.01|ICD9CM|Quadrplg c1-c4, complete|Quadrplg c1-c4, complete
C0376130|T047|PT|344.02|ICD9CM|Quadriplegia, C1-C4, incomplete|Quadriplegia, C1-C4, incomplete
C0376130|T047|AB|344.02|ICD9CM|Quadrplg c1-c4, incomplt|Quadrplg c1-c4, incomplt
C0376131|T047|PT|344.03|ICD9CM|Quadriplegia, C5-C7, complete|Quadriplegia, C5-C7, complete
C0376131|T047|AB|344.03|ICD9CM|Quadrplg c5-c7, complete|Quadrplg c5-c7, complete
C0376132|T047|PT|344.04|ICD9CM|Quadriplegia, C5-C7, incomplete|Quadriplegia, C5-C7, incomplete
C0376132|T047|AB|344.04|ICD9CM|Quadrplg c5-c7, incomplt|Quadrplg c5-c7, incomplt
C0375223|T184|AB|344.09|ICD9CM|Other quadriplegia|Other quadriplegia
C0375223|T184|PT|344.09|ICD9CM|Other quadriplegia|Other quadriplegia
C0030486|T047|PT|344.1|ICD9CM|Paraplegia|Paraplegia
C0030486|T047|AB|344.1|ICD9CM|Paraplegia NOS|Paraplegia NOS
C0154701|T047|AB|344.2|ICD9CM|Diplegia of upper limbs|Diplegia of upper limbs
C0154701|T047|PT|344.2|ICD9CM|Diplegia of upper limbs|Diplegia of upper limbs
C0154702|T047|HT|344.3|ICD9CM|Monoplegia of lower limb|Monoplegia of lower limb
C0375224|T184|PT|344.30|ICD9CM|Monoplegia of lower limb affecting unspecified side|Monoplegia of lower limb affecting unspecified side
C0375224|T184|AB|344.30|ICD9CM|Monplga lwr lmb unsp sde|Monplga lwr lmb unsp sde
C0375225|T047|PT|344.31|ICD9CM|Monoplegia of lower limb affecting dominant side|Monoplegia of lower limb affecting dominant side
C0375225|T047|AB|344.31|ICD9CM|Monplga lwr lmb dmnt sde|Monplga lwr lmb dmnt sde
C0859832|T184|AB|344.32|ICD9CM|Mnplg lwr lmb nondmnt sd|Mnplg lwr lmb nondmnt sd
C0859832|T184|PT|344.32|ICD9CM|Monoplegia of lower limb affecting nondominant side|Monoplegia of lower limb affecting nondominant side
C0154703|T047|HT|344.4|ICD9CM|Monoplegia of upper limb|Monoplegia of upper limb
C0154703|T047|PT|344.40|ICD9CM|Monoplegia of upper limb affecting unspecified side|Monoplegia of upper limb affecting unspecified side
C0154703|T047|AB|344.40|ICD9CM|Monplga upr lmb unsp sde|Monplga upr lmb unsp sde
C0375228|T047|PT|344.41|ICD9CM|Monoplegia of upper limb affecting dominant side|Monoplegia of upper limb affecting dominant side
C0375228|T047|AB|344.41|ICD9CM|Monplga upr lmb dmnt sde|Monplga upr lmb dmnt sde
C0375229|T184|AB|344.42|ICD9CM|Mnplg upr lmb nondmnt sd|Mnplg upr lmb nondmnt sd
C0375229|T184|PT|344.42|ICD9CM|Monoplegia of upper limb affecting nondominant sde|Monoplegia of upper limb affecting nondominant sde
C0085622|T047|AB|344.5|ICD9CM|Monoplegia NOS|Monoplegia NOS
C0085622|T047|PT|344.5|ICD9CM|Unspecified monoplegia|Unspecified monoplegia
C0392548|T047|HT|344.6|ICD9CM|Cauda equina syndrome|Cauda equina syndrome
C0270799|T047|AB|344.60|ICD9CM|Cauda equina synd NOS|Cauda equina synd NOS
C0270799|T047|PT|344.60|ICD9CM|Cauda equina syndrome without mention of neurogenic bladder|Cauda equina syndrome without mention of neurogenic bladder
C0007459|T047|PT|344.61|ICD9CM|Cauda equina syndrome with neurogenic bladder|Cauda equina syndrome with neurogenic bladder
C0007459|T047|AB|344.61|ICD9CM|Neurogenic bladder|Neurogenic bladder
C0154706|T047|HT|344.8|ICD9CM|Other specified paralytic syndromes|Other specified paralytic syndromes
C0023944|T047|AB|344.81|ICD9CM|Locked-in state|Locked-in state
C0023944|T047|PT|344.81|ICD9CM|Locked-in state|Locked-in state
C0154706|T047|AB|344.89|ICD9CM|Oth spcf paralytic synd|Oth spcf paralytic synd
C0154706|T047|PT|344.89|ICD9CM|Other specified paralytic syndrome|Other specified paralytic syndrome
C0522224|T033|AB|344.9|ICD9CM|Paralysis NOS|Paralysis NOS
C0522224|T033|PT|344.9|ICD9CM|Paralysis, unspecified|Paralysis, unspecified
C1719410|T047|HT|345|ICD9CM|Epilepsy and recurrent seizures|Epilepsy and recurrent seizures
C0017332|T047|HT|345.0|ICD9CM|Generalized nonconvulsive epilepsy|Generalized nonconvulsive epilepsy
C0154707|T047|AB|345.00|ICD9CM|Gen noncv ep w/o intr ep|Gen noncv ep w/o intr ep
C0154707|T047|PT|345.00|ICD9CM|Generalized nonconvulsive epilepsy, without mention of intractable epilepsy|Generalized nonconvulsive epilepsy, without mention of intractable epilepsy
C1112693|T047|AB|345.01|ICD9CM|Gen nonconv ep w intr ep|Gen nonconv ep w intr ep
C1112693|T047|PT|345.01|ICD9CM|Generalized nonconvulsive epilepsy, with intractable epilepsy|Generalized nonconvulsive epilepsy, with intractable epilepsy
C0311334|T047|HT|345.1|ICD9CM|Generalized convulsive epilepsy|Generalized convulsive epilepsy
C0154709|T047|AB|345.10|ICD9CM|Gen cnv epil w/o intr ep|Gen cnv epil w/o intr ep
C0154709|T047|PT|345.10|ICD9CM|Generalized convulsive epilepsy, without mention of intractable epilepsy|Generalized convulsive epilepsy, without mention of intractable epilepsy
C0154710|T047|AB|345.11|ICD9CM|Gen cnv epil w intr epil|Gen cnv epil w intr epil
C0154710|T047|PT|345.11|ICD9CM|Generalized convulsive epilepsy, with intractable epilepsy|Generalized convulsive epilepsy, with intractable epilepsy
C0270823|T047|AB|345.2|ICD9CM|Petit mal status|Petit mal status
C0270823|T047|PT|345.2|ICD9CM|Petit mal status|Petit mal status
C0311335|T047|AB|345.3|ICD9CM|Grand mal status|Grand mal status
C0311335|T047|PT|345.3|ICD9CM|Grand mal status|Grand mal status
C1306246|T047|AB|345.40|ICD9CM|Psymotr epil w/o int epi|Psymotr epil w/o int epi
C0154713|T047|AB|345.41|ICD9CM|Psymotr epil w intr epil|Psymotr epil w intr epil
C1719407|T047|HT|345.5|ICD9CM|Localization-related (focal) (partial) epilepsy and epileptic syndromes with simple partial seizures|Localization-related (focal) (partial) epilepsy and epileptic syndromes with simple partial seizures
C0154714|T047|AB|345.50|ICD9CM|Part epil w/o intr epil|Part epil w/o intr epil
C0154712|T047|AB|345.51|ICD9CM|Part epil w intr epil|Part epil w intr epil
C0037769|T047|HT|345.6|ICD9CM|Infantile spasms|Infantile spasms
C0154715|T046|AB|345.60|ICD9CM|Inf spasm w/o intr epil|Inf spasm w/o intr epil
C0154715|T046|PT|345.60|ICD9CM|Infantile spasms, without mention of intractable epilepsy|Infantile spasms, without mention of intractable epilepsy
C0154716|T046|AB|345.61|ICD9CM|Inf spasm w intract epil|Inf spasm w intract epil
C0154716|T046|PT|345.61|ICD9CM|Infantile spasms, with intractable epilepsy|Infantile spasms, with intractable epilepsy
C0085543|T047|HT|345.7|ICD9CM|Epilepsia partialis continua|Epilepsia partialis continua
C0154717|T047|AB|345.70|ICD9CM|Epil par cont w/o int ep|Epil par cont w/o int ep
C0154717|T047|PT|345.70|ICD9CM|Epilepsia partialis continua, without mention of intractable epilepsy|Epilepsia partialis continua, without mention of intractable epilepsy
C0154718|T047|AB|345.71|ICD9CM|Epil par cont w intr epi|Epil par cont w intr epi
C0154718|T047|PT|345.71|ICD9CM|Epilepsia partialis continua, with intractable epilepsy|Epilepsia partialis continua, with intractable epilepsy
C1719409|T047|HT|345.8|ICD9CM|Other forms of epilepsy and recurrent seizures|Other forms of epilepsy and recurrent seizures
C0154719|T047|AB|345.80|ICD9CM|Epilep NEC w/o intr epil|Epilep NEC w/o intr epil
C0154719|T047|PT|345.80|ICD9CM|Other forms of epilepsy and recurrent seizures, without mention of intractable epilepsy|Other forms of epilepsy and recurrent seizures, without mention of intractable epilepsy
C0154720|T047|AB|345.81|ICD9CM|Epilepsy NEC w intr epil|Epilepsy NEC w intr epil
C0154720|T047|PT|345.81|ICD9CM|Other forms of epilepsy and recurrent seizures, with intractable epilepsy|Other forms of epilepsy and recurrent seizures, with intractable epilepsy
C0014544|T047|HT|345.9|ICD9CM|Epilepsy, unspecified|Epilepsy, unspecified
C0154721|T047|AB|345.90|ICD9CM|Epilep NOS w/o intr epil|Epilep NOS w/o intr epil
C0154721|T047|PT|345.90|ICD9CM|Epilepsy, unspecified, without mention of intractable epilepsy|Epilepsy, unspecified, without mention of intractable epilepsy
C0154722|T047|AB|345.91|ICD9CM|Epilepsy NOS w intr epil|Epilepsy NOS w intr epil
C0154722|T047|PT|345.91|ICD9CM|Epilepsy, unspecified, with intractable epilepsy|Epilepsy, unspecified, with intractable epilepsy
C0149931|T047|HT|346|ICD9CM|Migraine|Migraine
C0154723|T047|HT|346.0|ICD9CM|Migraine with aura|Migraine with aura
C2349432|T047|AB|346.00|ICD9CM|Mgrn w aura wo ntrc mgrn|Mgrn w aura wo ntrc mgrn
C2349432|T047|PT|346.00|ICD9CM|Migraine with aura, without mention of intractable migraine without mention of status migrainosus|Migraine with aura, without mention of intractable migraine without mention of status migrainosus
C2349433|T047|AB|346.01|ICD9CM|Mgrn w aura w ntrc mgrn|Mgrn w aura w ntrc mgrn
C2349433|T047|PT|346.01|ICD9CM|Migraine with aura, with intractable migraine, so stated, without mention of status migrainosus|Migraine with aura, with intractable migraine, so stated, without mention of status migrainosus
C2349434|T047|AB|346.02|ICD9CM|Mgrn w aur wo ntrc mgrn|Mgrn w aur wo ntrc mgrn
C2349434|T047|PT|346.02|ICD9CM|Migraine with aura, without mention of intractable migraine with status migrainosus|Migraine with aura, without mention of intractable migraine with status migrainosus
C2349435|T047|AB|346.03|ICD9CM|Mgrn w aura w ntrc mgrn|Mgrn w aura w ntrc mgrn
C2349435|T047|PT|346.03|ICD9CM|Migraine with aura, with intractable migraine, so stated, with status migrainosus|Migraine with aura, with intractable migraine, so stated, with status migrainosus
C0338480|T047|HT|346.1|ICD9CM|Migraine without aura|Migraine without aura
C2349438|T047|AB|346.10|ICD9CM|Mgrn wo aura wo ntrc mgr|Mgrn wo aura wo ntrc mgr
C2349438|T047|PT|346.10|ICD9CM|Migraine without aura, without mention of intractable migraine without mention of status migrainosus|Migraine without aura, without mention of intractable migraine without mention of status migrainosus
C2349439|T047|AB|346.11|ICD9CM|Mgrn wo aura w ntrc mgrn|Mgrn wo aura w ntrc mgrn
C2349439|T047|PT|346.11|ICD9CM|Migraine without aura, with intractable migraine, so stated, without mention of status migrainosus|Migraine without aura, with intractable migraine, so stated, without mention of status migrainosus
C2349440|T047|AB|346.12|ICD9CM|Mgrn wo aura wo ntrc mgr|Mgrn wo aura wo ntrc mgr
C2349440|T047|PT|346.12|ICD9CM|Migraine without aura, without mention of intractable migraine with status migrainosus|Migraine without aura, without mention of intractable migraine with status migrainosus
C2349441|T047|AB|346.13|ICD9CM|Mgrn wo aura w ntrc mgrn|Mgrn wo aura w ntrc mgrn
C2349441|T047|PT|346.13|ICD9CM|Migraine without aura, with intractable migraine, so stated, with status migrainosus|Migraine without aura, with intractable migraine, so stated, with status migrainosus
C2349446|T047|HT|346.2|ICD9CM|Variants of migraine, not elsewhere classified|Variants of migraine, not elsewhere classified
C2349442|T047|AB|346.20|ICD9CM|Vrnt mgrn wo ntr mgr NEC|Vrnt mgrn wo ntr mgr NEC
C2349443|T047|AB|346.21|ICD9CM|Vrnt mgrn w ntrc mgr NEC|Vrnt mgrn w ntrc mgr NEC
C2349444|T047|AB|346.22|ICD9CM|Var mgr NEC wo ntc mgr|Var mgr NEC wo ntc mgr
C2349445|T047|AB|346.23|ICD9CM|Var mgrn NEC w ntrc mgr|Var mgrn NEC w ntrc mgr
C0270862|T047|HT|346.3|ICD9CM|Hemiplegic migraine|Hemiplegic migraine
C2349449|T047|PT|346.30|ICD9CM|Hemiplegic migraine, without mention of intractable migraine without mention of status migrainosus|Hemiplegic migraine, without mention of intractable migraine without mention of status migrainosus
C2349449|T047|AB|346.30|ICD9CM|Hmplg mgr wo ntrc wo st|Hmplg mgr wo ntrc wo st
C2349450|T047|PT|346.31|ICD9CM|Hemiplegic migraine, with intractable migraine, so stated, without mention of status migrainosus|Hemiplegic migraine, with intractable migraine, so stated, without mention of status migrainosus
C2349450|T047|AB|346.31|ICD9CM|Hmplg mgrn w ntrc wo st|Hmplg mgrn w ntrc wo st
C2349451|T047|PT|346.32|ICD9CM|Hemiplegic migraine, without mention of intractable migraine with status migrainosus|Hemiplegic migraine, without mention of intractable migraine with status migrainosus
C2349451|T047|AB|346.32|ICD9CM|Hemplg mgr wo ntrc w st|Hemplg mgr wo ntrc w st
C2349452|T047|PT|346.33|ICD9CM|Hemiplegic migraine, with intractable migraine, so stated, with status migrainosus|Hemiplegic migraine, with intractable migraine, so stated, with status migrainosus
C2349452|T047|AB|346.33|ICD9CM|Hmplg mgrn w ntrc w st|Hmplg mgrn w ntrc w st
C0269226|T046|HT|346.4|ICD9CM|Menstrual migraine|Menstrual migraine
C2349455|T047|AB|346.40|ICD9CM|Menst mgr wo ntrc wo st|Menst mgr wo ntrc wo st
C2349455|T047|PT|346.40|ICD9CM|Menstrual migraine, without mention of intractable migraine without mention of status migrainosus|Menstrual migraine, without mention of intractable migraine without mention of status migrainosus
C2349456|T047|AB|346.41|ICD9CM|Menstl mgrn w ntrc wo st|Menstl mgrn w ntrc wo st
C2349456|T047|PT|346.41|ICD9CM|Menstrual migraine, with intractable migraine, so stated, without mention of status migrainosus|Menstrual migraine, with intractable migraine, so stated, without mention of status migrainosus
C2349457|T047|AB|346.42|ICD9CM|Menstl mgr wo ntrc w st|Menstl mgr wo ntrc w st
C2349457|T047|PT|346.42|ICD9CM|Menstrual migraine, without mention of intractable migraine with status migrainosus|Menstrual migraine, without mention of intractable migraine with status migrainosus
C2349458|T047|AB|346.43|ICD9CM|Menstl mgrn w ntrc w st|Menstl mgrn w ntrc w st
C2349458|T047|PT|346.43|ICD9CM|Menstrual migraine, with intractable migraine, so stated, with status migrainosus|Menstrual migraine, with intractable migraine, so stated, with status migrainosus
C2349465|T046|HT|346.5|ICD9CM|Persistent migraine aura without cerebral infarction|Persistent migraine aura without cerebral infarction
C2349461|T047|AB|346.50|ICD9CM|Prst aura wo inf/ntr/st|Prst aura wo inf/ntr/st
C2349462|T047|AB|346.51|ICD9CM|Prs ara w ntr wo inf/st|Prs ara w ntr wo inf/st
C2349463|T047|AB|346.52|ICD9CM|Prs ara wo inf/ntr w st|Prs ara wo inf/ntr w st
C2349464|T047|AB|346.53|ICD9CM|Prs ara wo inf w ntr/st|Prs ara wo inf w ntr/st
C2349471|T047|HT|346.6|ICD9CM|Persistent migraine aura with cerebral infarction|Persistent migraine aura with cerebral infarction
C2349467|T047|AB|346.60|ICD9CM|Prs ara w inf wo ntr/st|Prs ara w inf wo ntr/st
C2349468|T047|AB|346.61|ICD9CM|Prs ara w/inf/ntr wo st|Prs ara w/inf/ntr wo st
C2349469|T047|AB|346.62|ICD9CM|Prs ara wo ntr w inf/st|Prs ara wo ntr w inf/st
C2349470|T047|AB|346.63|ICD9CM|Prst ara w inf w ntr/st|Prst ara w inf w ntr/st
C2349476|T047|HT|346.7|ICD9CM|Chronic migraine without aura|Chronic migraine without aura
C2349472|T047|AB|346.70|ICD9CM|Ch mgr wo ar wo nt wo st|Ch mgr wo ar wo nt wo st
C2349473|T047|AB|346.71|ICD9CM|Ch mgr wo ara w nt wo st|Ch mgr wo ara w nt wo st
C2349474|T047|AB|346.72|ICD9CM|Ch mgr wo ara wo nt w st|Ch mgr wo ara wo nt w st
C2349474|T047|PT|346.72|ICD9CM|Chronic migraine without aura, without mention of intractable migraine with status migrainosus|Chronic migraine without aura, without mention of intractable migraine with status migrainosus
C2349475|T047|AB|346.73|ICD9CM|Ch mgr wo ara w ntr w st|Ch mgr wo ara w ntr w st
C2349475|T047|PT|346.73|ICD9CM|Chronic migraine without aura, with intractable migraine, so stated, with status migrainosus|Chronic migraine without aura, with intractable migraine, so stated, with status migrainosus
C0477373|T047|HT|346.8|ICD9CM|Other forms of migraine|Other forms of migraine
C2362836|T047|AB|346.80|ICD9CM|Othr migrne wo ntrc mgrn|Othr migrne wo ntrc mgrn
C2349478|T047|PT|346.81|ICD9CM|Other forms of migraine, with intractable migraine, so stated, without mention of status migrainosus|Other forms of migraine, with intractable migraine, so stated, without mention of status migrainosus
C2349478|T047|AB|346.81|ICD9CM|Othr migrne w ntrc mgrne|Othr migrne w ntrc mgrne
C2349479|T047|AB|346.82|ICD9CM|Oth mgr wo ntrc w st mgr|Oth mgr wo ntrc w st mgr
C2349479|T047|PT|346.82|ICD9CM|Other forms of migraine, without mention of intractable migraine with status migrainosus|Other forms of migraine, without mention of intractable migraine with status migrainosus
C2349480|T047|AB|346.83|ICD9CM|Oth mgr w ntrc w st mgr|Oth mgr w ntrc w st mgr
C2349480|T047|PT|346.83|ICD9CM|Other forms of migraine, with intractable migraine, so stated, with status migrainosus|Other forms of migraine, with intractable migraine, so stated, with status migrainosus
C0149931|T047|HT|346.9|ICD9CM|Migraine, unspecified|Migraine, unspecified
C0375239|T047|PT|346.90|ICD9CM|Migraine, unspecified, without mention of intractable migraine without mention of status migrainosus|Migraine, unspecified, without mention of intractable migraine without mention of status migrainosus
C0375239|T047|AB|346.90|ICD9CM|Migrne unsp wo ntrc mgrn|Migrne unsp wo ntrc mgrn
C0375240|T047|AB|346.91|ICD9CM|Mgrn unsp w ntrc mgr std|Mgrn unsp w ntrc mgr std
C0375240|T047|PT|346.91|ICD9CM|Migraine, unspecified, with intractable migraine, so stated, without mention of status migrainosus|Migraine, unspecified, with intractable migraine, so stated, without mention of status migrainosus
C2349481|T047|AB|346.92|ICD9CM|Mgr NOS wo ntrc w st mgr|Mgr NOS wo ntrc w st mgr
C2349481|T047|PT|346.92|ICD9CM|Migraine, unspecified, without mention of intractable migraine with status migrainosus|Migraine, unspecified, without mention of intractable migraine with status migrainosus
C2349482|T047|AB|346.93|ICD9CM|Mgrn NOS w ntrc w st mgr|Mgrn NOS w ntrc w st mgr
C2349482|T047|PT|346.93|ICD9CM|Migraine, unspecified, with intractable migraine, so stated, with status migrainosus|Migraine, unspecified, with intractable migraine, so stated, with status migrainosus
C0751362|T047|HT|347|ICD9CM|Cataplexy and narcolepsy|Cataplexy and narcolepsy
C0027404|T047|HT|347.0|ICD9CM|Narcolepsy|Narcolepsy
C1456240|T047|AB|347.00|ICD9CM|Narcolepsy w/o cataplexy|Narcolepsy w/o cataplexy
C1456240|T047|PT|347.00|ICD9CM|Narcolepsy, without cataplexy|Narcolepsy, without cataplexy
C0751362|T047|AB|347.01|ICD9CM|Narcolepsy w cataplexy|Narcolepsy w cataplexy
C0751362|T047|PT|347.01|ICD9CM|Narcolepsy, with cataplexy|Narcolepsy, with cataplexy
C1456243|T047|HT|347.1|ICD9CM|Narcolepsy in conditions classified elsewhere|Narcolepsy in conditions classified elsewhere
C1456241|T047|AB|347.10|ICD9CM|Narclpsy w/o cat oth dis|Narclpsy w/o cat oth dis
C1456241|T047|PT|347.10|ICD9CM|Narcolepsy in conditions classified elsewhere, without cataplexy|Narcolepsy in conditions classified elsewhere, without cataplexy
C1456242|T047|PT|347.11|ICD9CM|Narcolepsy in conditions classified elsewhere, with cataplexy|Narcolepsy in conditions classified elsewhere, with cataplexy
C1456242|T047|AB|347.11|ICD9CM|Narcolepsy w cat oth dis|Narcolepsy w cat oth dis
C0029551|T047|HT|348|ICD9CM|Other conditions of brain|Other conditions of brain
C0154724|T047|AB|348.0|ICD9CM|Cerebral cysts|Cerebral cysts
C0154724|T047|PT|348.0|ICD9CM|Cerebral cysts|Cerebral cysts
C0003132|T046|AB|348.1|ICD9CM|Anoxic brain damage|Anoxic brain damage
C0003132|T046|PT|348.1|ICD9CM|Anoxic brain damage|Anoxic brain damage
C0033845|T047|PT|348.2|ICD9CM|Benign intracranial hypertension|Benign intracranial hypertension
C0033845|T047|AB|348.2|ICD9CM|Pseudotumor cerebri|Pseudotumor cerebri
C0085584|T047|HT|348.3|ICD9CM|Encephalopathy, not elsewhere classified|Encephalopathy, not elsewhere classified
C0085584|T047|AB|348.30|ICD9CM|Encephalopathy NOS|Encephalopathy NOS
C0085584|T047|PT|348.30|ICD9CM|Encephalopathy, unspecified|Encephalopathy, unspecified
C0006112|T047|AB|348.31|ICD9CM|Metabolic encephalopathy|Metabolic encephalopathy
C0006112|T047|PT|348.31|ICD9CM|Metabolic encephalopathy|Metabolic encephalopathy
C1260408|T047|AB|348.39|ICD9CM|Encephalopathy NEC|Encephalopathy NEC
C1260408|T047|PT|348.39|ICD9CM|Other encephalopathy|Other encephalopathy
C0009592|T047|AB|348.4|ICD9CM|Compression of brain|Compression of brain
C0009592|T047|PT|348.4|ICD9CM|Compression of brain|Compression of brain
C0006114|T046|AB|348.5|ICD9CM|Cerebral edema|Cerebral edema
C0006114|T046|PT|348.5|ICD9CM|Cerebral edema|Cerebral edema
C0029551|T047|HT|348.8|ICD9CM|Other conditions of brain|Other conditions of brain
C2712987|T047|AB|348.81|ICD9CM|Temporal sclerosis|Temporal sclerosis
C2712987|T047|PT|348.81|ICD9CM|Temporal sclerosis|Temporal sclerosis
C0006110|T046|AB|348.82|ICD9CM|Brain death|Brain death
C0006110|T046|PT|348.82|ICD9CM|Brain death|Brain death
C2712887|T047|AB|348.89|ICD9CM|Brain conditions NEC|Brain conditions NEC
C2712887|T047|PT|348.89|ICD9CM|Other conditions of brain|Other conditions of brain
C0006111|T047|AB|348.9|ICD9CM|Brain condition NOS|Brain condition NOS
C0006111|T047|PT|348.9|ICD9CM|Unspecified condition of brain|Unspecified condition of brain
C0154725|T047|HT|349|ICD9CM|Other and unspecified disorders of the nervous system|Other and unspecified disorders of the nervous system
C0701795|T033|AB|349.0|ICD9CM|Lumbar puncture reaction|Lumbar puncture reaction
C0701795|T033|PT|349.0|ICD9CM|Reaction to spinal or lumbar puncture|Reaction to spinal or lumbar puncture
C0154727|T047|AB|349.1|ICD9CM|Complication cns device|Complication cns device
C0154727|T047|PT|349.1|ICD9CM|Nervous system complications from surgically implanted device|Nervous system complications from surgically implanted device
C0795685|T047|AB|349.2|ICD9CM|Disorder of meninges NEC|Disorder of meninges NEC
C0795685|T047|PT|349.2|ICD9CM|Disorders of meninges, not elsewhere classified|Disorders of meninges, not elsewhere classified
C1504340|T037|HT|349.3|ICD9CM|Dural tear|Dural tear
C2349483|T037|AB|349.31|ICD9CM|Accid punc/op lac dura|Accid punc/op lac dura
C2349483|T037|PT|349.31|ICD9CM|Accidental puncture or laceration of dura during a procedure|Accidental puncture or laceration of dura during a procedure
C2349485|T047|AB|349.39|ICD9CM|Dural tear NEC|Dural tear NEC
C2349485|T047|PT|349.39|ICD9CM|Other dural tear|Other dural tear
C0029784|T047|HT|349.8|ICD9CM|Other specified disorders of nervous system|Other specified disorders of nervous system
C0007815|T047|PT|349.81|ICD9CM|Cerebrospinal fluid rhinorrhea|Cerebrospinal fluid rhinorrhea
C0007815|T047|AB|349.81|ICD9CM|Cerebrospinal rhinorrhea|Cerebrospinal rhinorrhea
C0149504|T037|AB|349.82|ICD9CM|Toxic encephalopathy|Toxic encephalopathy
C0149504|T037|PT|349.82|ICD9CM|Toxic encephalopathy|Toxic encephalopathy
C0029784|T047|AB|349.89|ICD9CM|Cns disorder NEC|Cns disorder NEC
C0029784|T047|PT|349.89|ICD9CM|Other specified disorders of nervous system|Other specified disorders of nervous system
C0027765|T047|AB|349.9|ICD9CM|Cns disorder NOS|Cns disorder NOS
C0027765|T047|PT|349.9|ICD9CM|Unspecified disorders of nervous system|Unspecified disorders of nervous system
C0152177|T047|HT|350|ICD9CM|Trigeminal nerve disorders|Trigeminal nerve disorders
C4721453|T047|HT|350-359.99|ICD9CM|DISORDERS OF THE PERIPHERAL NERVOUS SYSTEM|DISORDERS OF THE PERIPHERAL NERVOUS SYSTEM
C0040997|T047|AB|350.1|ICD9CM|Trigeminal neuralgia|Trigeminal neuralgia
C0040997|T047|PT|350.1|ICD9CM|Trigeminal neuralgia|Trigeminal neuralgia
C0154729|T184|AB|350.2|ICD9CM|Atypical face pain|Atypical face pain
C0154729|T184|PT|350.2|ICD9CM|Atypical face pain|Atypical face pain
C0029834|T047|PT|350.8|ICD9CM|Other specified trigeminal nerve disorders|Other specified trigeminal nerve disorders
C0029834|T047|AB|350.8|ICD9CM|Trigeminal nerve dis NEC|Trigeminal nerve dis NEC
C0152177|T047|AB|350.9|ICD9CM|Trigeminal nerve dis NOS|Trigeminal nerve dis NOS
C0152177|T047|PT|350.9|ICD9CM|Trigeminal nerve disorder, unspecified|Trigeminal nerve disorder, unspecified
C0015464|T047|HT|351|ICD9CM|Facial nerve disorders|Facial nerve disorders
C0376175|T047|AB|351.0|ICD9CM|Bell's palsy|Bell's palsy
C0376175|T047|PT|351.0|ICD9CM|Bell's palsy|Bell's palsy
C0017407|T047|AB|351.1|ICD9CM|Geniculate ganglionitis|Geniculate ganglionitis
C0017407|T047|PT|351.1|ICD9CM|Geniculate ganglionitis|Geniculate ganglionitis
C0029616|T047|AB|351.8|ICD9CM|Facial nerve dis NEC|Facial nerve dis NEC
C0029616|T047|PT|351.8|ICD9CM|Other facial nerve disorders|Other facial nerve disorders
C0015464|T047|AB|351.9|ICD9CM|Facial nerve dis NOS|Facial nerve dis NOS
C0015464|T047|PT|351.9|ICD9CM|Facial nerve disorder, unspecified|Facial nerve disorder, unspecified
C0154730|T047|HT|352|ICD9CM|Disorders of other cranial nerves|Disorders of other cranial nerves
C0751937|T047|PT|352.0|ICD9CM|Disorders of olfactory (1st) nerve|Disorders of olfactory (1st) nerve
C0751937|T047|AB|352.0|ICD9CM|Olfactory nerve disorder|Olfactory nerve disorder
C0154731|T047|AB|352.1|ICD9CM|Glossopharyng neuralgia|Glossopharyng neuralgia
C0154731|T047|PT|352.1|ICD9CM|Glossopharyngeal neuralgia|Glossopharyngeal neuralgia
C0393797|T047|AB|352.2|ICD9CM|Glossophar nerve dis NEC|Glossophar nerve dis NEC
C0393797|T047|PT|352.2|ICD9CM|Other disorders of glossopharyngeal [9th] nerve|Other disorders of glossopharyngeal [9th] nerve
C0152179|T047|PT|352.3|ICD9CM|Disorders of pneumogastric [10th] nerve|Disorders of pneumogastric [10th] nerve
C0152179|T047|AB|352.3|ICD9CM|Pneumogastric nerve dis|Pneumogastric nerve dis
C0152180|T047|AB|352.4|ICD9CM|Accessory nerve disorder|Accessory nerve disorder
C0152180|T047|PT|352.4|ICD9CM|Disorders of accessory [11th] nerve|Disorders of accessory [11th] nerve
C0152181|T047|PT|352.5|ICD9CM|Disorders of hypoglossal [12th] nerve|Disorders of hypoglossal [12th] nerve
C0152181|T047|AB|352.5|ICD9CM|Hypoglossal nerve dis|Hypoglossal nerve dis
C0154733|T047|AB|352.6|ICD9CM|Mult cranial nerve palsy|Mult cranial nerve palsy
C0154733|T047|PT|352.6|ICD9CM|Multiple cranial nerve palsies|Multiple cranial nerve palsies
C0010266|T047|AB|352.9|ICD9CM|Cranial nerve dis NOS|Cranial nerve dis NOS
C0010266|T047|PT|352.9|ICD9CM|Unspecified disorder of cranial nerves|Unspecified disorder of cranial nerves
C0270890|T047|HT|353|ICD9CM|Nerve root and plexus disorders|Nerve root and plexus disorders
C0006091|T047|AB|353.0|ICD9CM|Brachial plexus lesions|Brachial plexus lesions
C0006091|T047|PT|353.0|ICD9CM|Brachial plexus lesions|Brachial plexus lesions
C0154735|T047|AB|353.1|ICD9CM|Lumbosacral plex lesion|Lumbosacral plex lesion
C0154735|T047|PT|353.1|ICD9CM|Lumbosacral plexus lesions|Lumbosacral plexus lesions
C0869208|T047|AB|353.2|ICD9CM|Cervical root lesion NEC|Cervical root lesion NEC
C0869208|T047|PT|353.2|ICD9CM|Cervical root lesions, not elsewhere classified|Cervical root lesions, not elsewhere classified
C0868842|T047|AB|353.3|ICD9CM|Thoracic root lesion NEC|Thoracic root lesion NEC
C0868842|T047|PT|353.3|ICD9CM|Thoracic root lesions, not elsewhere classified|Thoracic root lesions, not elsewhere classified
C0869447|T047|PT|353.4|ICD9CM|Lumbosacral root lesions, not elsewhere classified|Lumbosacral root lesions, not elsewhere classified
C0869447|T047|AB|353.4|ICD9CM|Lumbsacral root les NEC|Lumbsacral root les NEC
C1510479|T047|AB|353.5|ICD9CM|Neuralgic amyotrophy|Neuralgic amyotrophy
C1510479|T047|PT|353.5|ICD9CM|Neuralgic amyotrophy|Neuralgic amyotrophy
C0031315|T047|AB|353.6|ICD9CM|Phantom limb (syndrome)|Phantom limb (syndrome)
C0031315|T047|PT|353.6|ICD9CM|Phantom limb (syndrome)|Phantom limb (syndrome)
C0154739|T047|AB|353.8|ICD9CM|Nerv root/plexus dis NEC|Nerv root/plexus dis NEC
C0154739|T047|PT|353.8|ICD9CM|Other nerve root and plexus disorders|Other nerve root and plexus disorders
C0270890|T047|AB|353.9|ICD9CM|Nerv root/plexus dis NOS|Nerv root/plexus dis NOS
C0270890|T047|PT|353.9|ICD9CM|Unspecified nerve root and plexus disorder|Unspecified nerve root and plexus disorder
C0154741|T047|HT|354|ICD9CM|Mononeuritis of upper limb and mononeuritis multiplex|Mononeuritis of upper limb and mononeuritis multiplex
C0007286|T047|AB|354.0|ICD9CM|Carpal tunnel syndrome|Carpal tunnel syndrome
C0007286|T047|PT|354.0|ICD9CM|Carpal tunnel syndrome|Carpal tunnel syndrome
C0154742|T046|AB|354.1|ICD9CM|Median nerve lesion NEC|Median nerve lesion NEC
C0154742|T046|PT|354.1|ICD9CM|Other lesion of median nerve|Other lesion of median nerve
C1288279|T047|PT|354.2|ICD9CM|Lesion of ulnar nerve|Lesion of ulnar nerve
C1288279|T047|AB|354.2|ICD9CM|Ulnar nerve lesion|Ulnar nerve lesion
C0154744|T047|PT|354.3|ICD9CM|Lesion of radial nerve|Lesion of radial nerve
C0154744|T047|AB|354.3|ICD9CM|Radial nerve lesion|Radial nerve lesion
C1443291|T047|PT|354.4|ICD9CM|Causalgia of upper limb|Causalgia of upper limb
C1443291|T047|AB|354.4|ICD9CM|Causalgia upper limb|Causalgia upper limb
C0151295|T047|AB|354.5|ICD9CM|Mononeuritis multiplex|Mononeuritis multiplex
C0151295|T047|PT|354.5|ICD9CM|Mononeuritis multiplex|Mononeuritis multiplex
C0154745|T047|AB|354.8|ICD9CM|Mononeuritis arm NEC|Mononeuritis arm NEC
C0154745|T047|PT|354.8|ICD9CM|Other mononeuritis of upper limb|Other mononeuritis of upper limb
C0154746|T047|AB|354.9|ICD9CM|Mononeuritis arm NOS|Mononeuritis arm NOS
C0154746|T047|PT|354.9|ICD9CM|Mononeuritis of upper limb, unspecified|Mononeuritis of upper limb, unspecified
C0154747|T047|HT|355|ICD9CM|Mononeuritis of lower limb|Mononeuritis of lower limb
C0154748|T047|PT|355.0|ICD9CM|Lesion of sciatic nerve|Lesion of sciatic nerve
C0154748|T047|AB|355.0|ICD9CM|Sciatic nerve lesion|Sciatic nerve lesion
C0152110|T047|AB|355.1|ICD9CM|Meralgia paresthetica|Meralgia paresthetica
C0152110|T047|PT|355.1|ICD9CM|Meralgia paresthetica|Meralgia paresthetica
C0154749|T047|AB|355.2|ICD9CM|Femoral nerve lesion NEC|Femoral nerve lesion NEC
C0154749|T047|PT|355.2|ICD9CM|Other lesion of femoral nerve|Other lesion of femoral nerve
C0270909|T047|AB|355.3|ICD9CM|Lat popliteal nerve les|Lat popliteal nerve les
C0270909|T047|PT|355.3|ICD9CM|Lesion of lateral popliteal nerve|Lesion of lateral popliteal nerve
C1302325|T047|PT|355.4|ICD9CM|Lesion of medial popliteal nerve|Lesion of medial popliteal nerve
C1302325|T047|AB|355.4|ICD9CM|Med popliteal nerve les|Med popliteal nerve les
C0039319|T047|AB|355.5|ICD9CM|Tarsal tunnel syndrome|Tarsal tunnel syndrome
C0039319|T047|PT|355.5|ICD9CM|Tarsal tunnel syndrome|Tarsal tunnel syndrome
C0154752|T047|PT|355.6|ICD9CM|Lesion of plantar nerve|Lesion of plantar nerve
C0154752|T047|AB|355.6|ICD9CM|Plantar nerve lesion|Plantar nerve lesion
C0154753|T047|HT|355.7|ICD9CM|Other mononeuritis of lower limb|Other mononeuritis of lower limb
C0375242|T047|AB|355.71|ICD9CM|Causalgia lower limb|Causalgia lower limb
C0375242|T047|PT|355.71|ICD9CM|Causalgia of lower limb|Causalgia of lower limb
C0154753|T047|AB|355.79|ICD9CM|Oth mononeur lower limb|Oth mononeur lower limb
C0154753|T047|PT|355.79|ICD9CM|Other mononeuritis of lower limb|Other mononeuritis of lower limb
C0154747|T047|AB|355.8|ICD9CM|Mononeuritis leg NOS|Mononeuritis leg NOS
C0154747|T047|PT|355.8|ICD9CM|Mononeuritis of lower limb, unspecified|Mononeuritis of lower limb, unspecified
C0235880|T047|AB|355.9|ICD9CM|Mononeuritis NOS|Mononeuritis NOS
C0235880|T047|PT|355.9|ICD9CM|Mononeuritis of unspecified site|Mononeuritis of unspecified site
C0154754|T047|HT|356|ICD9CM|Hereditary and idiopathic peripheral neuropathy|Hereditary and idiopathic peripheral neuropathy
C0392553|T047|AB|356.0|ICD9CM|Hered periph neuropathy|Hered periph neuropathy
C0392553|T047|PT|356.0|ICD9CM|Hereditary peripheral neuropathy|Hereditary peripheral neuropathy
C0007959|T047|AB|356.1|ICD9CM|Peroneal muscle atrophy|Peroneal muscle atrophy
C0007959|T047|PT|356.1|ICD9CM|Peroneal muscular atrophy|Peroneal muscular atrophy
C0699739|T047|AB|356.2|ICD9CM|Hered sensory neuropathy|Hered sensory neuropathy
C0699739|T047|PT|356.2|ICD9CM|Hereditary sensory neuropathy|Hereditary sensory neuropathy
C0034960|T047|AB|356.3|ICD9CM|Refsum's disease|Refsum's disease
C0034960|T047|PT|356.3|ICD9CM|Refsum's disease|Refsum's disease
C0154756|T047|AB|356.4|ICD9CM|Idio prog polyneuropathy|Idio prog polyneuropathy
C0154756|T047|PT|356.4|ICD9CM|Idiopathic progressive polyneuropathy|Idiopathic progressive polyneuropathy
C0154757|T047|AB|356.8|ICD9CM|Idio periph neurpthy NEC|Idio periph neurpthy NEC
C0154757|T047|PT|356.8|ICD9CM|Other specified idiopathic peripheral neuropathy|Other specified idiopathic peripheral neuropathy
C0859673|T047|AB|356.9|ICD9CM|Idio periph neurpthy NOS|Idio periph neurpthy NOS
C0859673|T047|PT|356.9|ICD9CM|Unspecified hereditary and idiopathic peripheral neuropathy|Unspecified hereditary and idiopathic peripheral neuropathy
C0154758|T046|HT|357|ICD9CM|Inflammatory and toxic neuropathy|Inflammatory and toxic neuropathy
C3542501|T047|AB|357.0|ICD9CM|Ac infect polyneuritis|Ac infect polyneuritis
C3542501|T047|PT|357.0|ICD9CM|Acute infective polyneuritis|Acute infective polyneuritis
C0154759|T047|AB|357.1|ICD9CM|Neurpthy in col vasc dis|Neurpthy in col vasc dis
C0154759|T047|PT|357.1|ICD9CM|Polyneuropathy in collagen vascular disease|Polyneuropathy in collagen vascular disease
C0271680|T047|AB|357.2|ICD9CM|Neuropathy in diabetes|Neuropathy in diabetes
C0271680|T047|PT|357.2|ICD9CM|Polyneuropathy in diabetes|Polyneuropathy in diabetes
C0270932|T047|AB|357.3|ICD9CM|Neuropathy in malig dis|Neuropathy in malig dis
C0270932|T047|PT|357.3|ICD9CM|Polyneuropathy in malignant disease|Polyneuropathy in malignant disease
C0154761|T047|AB|357.4|ICD9CM|Neuropathy in other dis|Neuropathy in other dis
C0154761|T047|PT|357.4|ICD9CM|Polyneuropathy in other diseases classified elsewhere|Polyneuropathy in other diseases classified elsewhere
C0085677|T047|AB|357.5|ICD9CM|Alcoholic polyneuropathy|Alcoholic polyneuropathy
C0085677|T047|PT|357.5|ICD9CM|Alcoholic polyneuropathy|Alcoholic polyneuropathy
C0154762|T047|AB|357.6|ICD9CM|Neuropathy due to drugs|Neuropathy due to drugs
C0154762|T047|PT|357.6|ICD9CM|Polyneuropathy due to drugs|Polyneuropathy due to drugs
C0154763|T047|AB|357.7|ICD9CM|Neurpthy toxic agent NEC|Neurpthy toxic agent NEC
C0154763|T047|PT|357.7|ICD9CM|Polyneuropathy due to other toxic agents|Polyneuropathy due to other toxic agents
C0154764|T047|HT|357.8|ICD9CM|Other inflammatory and toxic neuropathies|Other inflammatory and toxic neuropathies
C0393819|T047|AB|357.81|ICD9CM|Chr inflam polyneuritis|Chr inflam polyneuritis
C0393819|T047|PT|357.81|ICD9CM|Chronic inflammatory demyelinating polyneuritis|Chronic inflammatory demyelinating polyneuritis
C0393851|T047|AB|357.82|ICD9CM|Crit illness neuropathy|Crit illness neuropathy
C0393851|T047|PT|357.82|ICD9CM|Critical illness polyneuropathy|Critical illness polyneuropathy
C0154764|T047|AB|357.89|ICD9CM|Inflam/tox neuropthy NEC|Inflam/tox neuropthy NEC
C0154764|T047|PT|357.89|ICD9CM|Other inflammatory and toxic neuropathy|Other inflammatory and toxic neuropathy
C0154758|T046|AB|357.9|ICD9CM|Inflam/tox neuropthy NOS|Inflam/tox neuropthy NOS
C0154758|T046|PT|357.9|ICD9CM|Unspecified inflammatory and toxic neuropathy|Unspecified inflammatory and toxic neuropathy
C0027868|T047|HT|358|ICD9CM|Myoneural disorders|Myoneural disorders
C0026896|T047|HT|358.0|ICD9CM|Myasthenia gravis|Myasthenia gravis
C1260409|T047|PT|358.00|ICD9CM|Myasthenia gravis without (acute) exacerbation|Myasthenia gravis without (acute) exacerbation
C1260409|T047|AB|358.00|ICD9CM|Mysthna grvs w/o ac exac|Mysthna grvs w/o ac exac
C0270942|T047|PT|358.01|ICD9CM|Myasthenia gravis with (acute) exacerbation|Myasthenia gravis with (acute) exacerbation
C0270942|T047|AB|358.01|ICD9CM|Myasthna gravs w ac exac|Myasthna gravs w ac exac
C0026897|T047|AB|358.1|ICD9CM|Myasthenia in oth dis|Myasthenia in oth dis
C0026897|T047|PT|358.1|ICD9CM|Myasthenic syndromes in diseases classified elsewhere|Myasthenic syndromes in diseases classified elsewhere
C0393939|T047|AB|358.2|ICD9CM|Toxic myoneural disorder|Toxic myoneural disorder
C0393939|T047|PT|358.2|ICD9CM|Toxic myoneural disorders|Toxic myoneural disorders
C0022972|T047|HT|358.3|ICD9CM|Lambert-Eaton syndrome|Lambert-Eaton syndrome
C3161080|T047|AB|358.30|ICD9CM|Lambert-Eaton synd NOS|Lambert-Eaton synd NOS
C3161080|T047|PT|358.30|ICD9CM|Lambert-Eaton syndrome, unspecified|Lambert-Eaton syndrome, unspecified
C3161081|T047|AB|358.31|ICD9CM|Lambert-Eaton synd neopl|Lambert-Eaton synd neopl
C3161081|T047|PT|358.31|ICD9CM|Lambert-Eaton syndrome in neoplastic disease|Lambert-Eaton syndrome in neoplastic disease
C3161082|T047|AB|358.39|ICD9CM|Lambert-Eaton syn ot dis|Lambert-Eaton syn ot dis
C3161082|T047|PT|358.39|ICD9CM|Lambert-Eaton syndrome in other diseases classified elsewhere|Lambert-Eaton syndrome in other diseases classified elsewhere
C0029816|T047|AB|358.8|ICD9CM|Myoneural disorders NEC|Myoneural disorders NEC
C0029816|T047|PT|358.8|ICD9CM|Other specified myoneural disorders|Other specified myoneural disorders
C0027868|T047|AB|358.9|ICD9CM|Myoneural disorders NOS|Myoneural disorders NOS
C0027868|T047|PT|358.9|ICD9CM|Myoneural disorders, unspecified|Myoneural disorders, unspecified
C0026849|T047|HT|359|ICD9CM|Muscular dystrophies and other myopathies|Muscular dystrophies and other myopathies
C2937300|T019|AB|359.0|ICD9CM|Cong hered musc dystrphy|Cong hered musc dystrphy
C2937300|T047|AB|359.0|ICD9CM|Cong hered musc dystrphy|Cong hered musc dystrphy
C2937300|T019|PT|359.0|ICD9CM|Congenital hereditary muscular dystrophy|Congenital hereditary muscular dystrophy
C2937300|T047|PT|359.0|ICD9CM|Congenital hereditary muscular dystrophy|Congenital hereditary muscular dystrophy
C4551827|T047|AB|359.1|ICD9CM|Hered prog musc dystrphy|Hered prog musc dystrphy
C4551827|T047|PT|359.1|ICD9CM|Hereditary progressive muscular dystrophy|Hereditary progressive muscular dystrophy
C0553604|T047|HT|359.2|ICD9CM|Myotonic disorders|Myotonic disorders
C0027126|T047|AB|359.21|ICD9CM|Myotonic musclr dystrphy|Myotonic musclr dystrphy
C0027126|T047|PT|359.21|ICD9CM|Myotonic muscular dystrophy|Myotonic muscular dystrophy
C0027127|T047|PT|359.22|ICD9CM|Myotonia congenita|Myotonia congenita
C0027127|T047|AB|359.22|ICD9CM|Myotonia congenita|Myotonia congenita
C0036391|T047|PT|359.23|ICD9CM|Myotonic chondrodystrophy|Myotonic chondrodystrophy
C0036391|T047|AB|359.23|ICD9CM|Myotonic chondrodystrphy|Myotonic chondrodystrphy
C1404542|T046|AB|359.24|ICD9CM|Drug induced myotonia|Drug induced myotonia
C1404542|T046|PT|359.24|ICD9CM|Drug- induced myotonia|Drug- induced myotonia
C0410224|T047|AB|359.29|ICD9CM|Myotonic disorder NEC|Myotonic disorder NEC
C0410224|T047|PT|359.29|ICD9CM|Other specified myotonic disorder|Other specified myotonic disorder
C1279412|T047|PT|359.3|ICD9CM|Periodic paralysis|Periodic paralysis
C1279412|T047|AB|359.3|ICD9CM|Periodic paralysis|Periodic paralysis
C0154769|T047|AB|359.4|ICD9CM|Toxic myopathy|Toxic myopathy
C0154769|T047|PT|359.4|ICD9CM|Toxic myopathy|Toxic myopathy
C0154770|T047|AB|359.5|ICD9CM|Myopathy in endocrin dis|Myopathy in endocrin dis
C0154770|T047|PT|359.5|ICD9CM|Myopathy in endocrine diseases classified elsewhere|Myopathy in endocrine diseases classified elsewhere
C0154771|T047|AB|359.6|ICD9CM|Infl myopathy in oth dis|Infl myopathy in oth dis
C0154771|T047|PT|359.6|ICD9CM|Symptomatic inflammatory myopathy in diseases classified elsewhere|Symptomatic inflammatory myopathy in diseases classified elsewhere
C2712761|T047|HT|359.7|ICD9CM|Inflammatory and immune myopathies, NEC|Inflammatory and immune myopathies, NEC
C0238190|T047|AB|359.71|ICD9CM|Inclusion body myositis|Inclusion body myositis
C0238190|T047|PT|359.71|ICD9CM|Inclusion body myositis|Inclusion body myositis
C2712808|T047|AB|359.79|ICD9CM|Inflm/immune myopath NEC|Inflm/immune myopath NEC
C2712808|T047|PT|359.79|ICD9CM|Other inflammatory and immune myopathies, NEC|Other inflammatory and immune myopathies, NEC
C0546839|T047|HT|359.8|ICD9CM|Other myopathies|Other myopathies
C1135188|T047|PT|359.81|ICD9CM|Critical illness myopathy|Critical illness myopathy
C1135188|T047|AB|359.81|ICD9CM|Critical illness myopthy|Critical illness myopthy
C0546839|T047|AB|359.89|ICD9CM|Myopathies NEC|Myopathies NEC
C0546839|T047|PT|359.89|ICD9CM|Other myopathies|Other myopathies
C0026848|T047|AB|359.9|ICD9CM|Myopathy NOS|Myopathy NOS
C0026848|T047|PT|359.9|ICD9CM|Myopathy, unspecified|Myopathy, unspecified
C0015397|T047|HT|360|ICD9CM|Disorders of the globe|Disorders of the globe
C1314803|T047|HT|360-379.99|ICD9CM|DISORDERS OF THE EYE AND ADNEXA|DISORDERS OF THE EYE AND ADNEXA
C0259800|T047|HT|360.0|ICD9CM|Purulent endophthalmitis|Purulent endophthalmitis
C0259800|T047|AB|360.00|ICD9CM|Purulent endophthalm NOS|Purulent endophthalm NOS
C0259800|T047|PT|360.00|ICD9CM|Purulent endophthalmitis, unspecified|Purulent endophthalmitis, unspecified
C0154773|T047|AB|360.01|ICD9CM|Acute endophthalmitis|Acute endophthalmitis
C0154773|T047|PT|360.01|ICD9CM|Acute endophthalmitis|Acute endophthalmitis
C0030332|T047|AB|360.02|ICD9CM|Panophthalmitis|Panophthalmitis
C0030332|T047|PT|360.02|ICD9CM|Panophthalmitis|Panophthalmitis
C0154774|T047|AB|360.03|ICD9CM|Chronic endophthalmitis|Chronic endophthalmitis
C0154774|T047|PT|360.03|ICD9CM|Chronic endophthalmitis|Chronic endophthalmitis
C0042904|T047|AB|360.04|ICD9CM|Vitreous abscess|Vitreous abscess
C0042904|T047|PT|360.04|ICD9CM|Vitreous abscess|Vitreous abscess
C0029610|T047|HT|360.1|ICD9CM|Other endophthalmitis|Other endophthalmitis
C0029077|T047|AB|360.11|ICD9CM|Sympathetic uveitis|Sympathetic uveitis
C0029077|T047|PT|360.11|ICD9CM|Sympathetic uveitis|Sympathetic uveitis
C0030343|T047|AB|360.12|ICD9CM|Panuveitis|Panuveitis
C0030343|T047|PT|360.12|ICD9CM|Panuveitis|Panuveitis
C0014238|T047|AB|360.13|ICD9CM|Parasitic endophthal NOS|Parasitic endophthal NOS
C0014238|T047|PT|360.13|ICD9CM|Parasitic endophthalmitis NOS|Parasitic endophthalmitis NOS
C0154775|T047|AB|360.14|ICD9CM|Ophthalmia nodosa|Ophthalmia nodosa
C0154775|T047|PT|360.14|ICD9CM|Ophthalmia nodosa|Ophthalmia nodosa
C0029610|T047|AB|360.19|ICD9CM|Endophthalmitis NEC|Endophthalmitis NEC
C0029610|T047|PT|360.19|ICD9CM|Other endophthalmitis|Other endophthalmitis
C0154777|T047|HT|360.2|ICD9CM|Degenerative disorders of globe|Degenerative disorders of globe
C0154777|T047|AB|360.20|ICD9CM|Degenerat globe dis NOS|Degenerat globe dis NOS
C0154777|T047|PT|360.20|ICD9CM|Degenerative disorder of globe, unspecified|Degenerative disorder of globe, unspecified
C0154778|T047|PT|360.21|ICD9CM|Progressive high (degenerative) myopia|Progressive high (degenerative) myopia
C0154778|T047|AB|360.21|ICD9CM|Progressive high myopia|Progressive high myopia
C0271001|T047|AB|360.23|ICD9CM|Siderosis|Siderosis
C0271001|T047|PT|360.23|ICD9CM|Siderosis of globe|Siderosis of globe
C0339034|T047|PT|360.24|ICD9CM|Other metallosis of globe|Other metallosis of globe
C0339034|T047|AB|360.24|ICD9CM|Other metallosis, eye|Other metallosis, eye
C0154780|T047|AB|360.29|ICD9CM|Degenerative globe NEC|Degenerative globe NEC
C0154780|T047|PT|360.29|ICD9CM|Other degenerative disorders of globe|Other degenerative disorders of globe
C0028841|T047|HT|360.3|ICD9CM|Hypotony of eye|Hypotony of eye
C0028841|T047|AB|360.30|ICD9CM|Hypotony NOS, eye|Hypotony NOS, eye
C0028841|T047|PT|360.30|ICD9CM|Hypotony of eye, unspecified|Hypotony of eye, unspecified
C0154782|T047|AB|360.31|ICD9CM|Primary hypotony|Primary hypotony
C0154782|T047|PT|360.31|ICD9CM|Primary hypotony of eye|Primary hypotony of eye
C0154783|T190|AB|360.32|ICD9CM|Hypotony due to fistula|Hypotony due to fistula
C0154783|T190|PT|360.32|ICD9CM|Ocular fistula causing hypotony|Ocular fistula causing hypotony
C0154784|T047|PT|360.33|ICD9CM|Hypotony associated with other ocular disorders|Hypotony associated with other ocular disorders
C0154784|T047|AB|360.33|ICD9CM|Hypotony w eye dis NEC|Hypotony w eye dis NEC
C0271004|T190|AB|360.34|ICD9CM|Flat anterior chamber|Flat anterior chamber
C0271004|T190|PT|360.34|ICD9CM|Flat anterior chamber of eye|Flat anterior chamber of eye
C0154777|T047|HT|360.4|ICD9CM|Degenerated conditions of globe|Degenerated conditions of globe
C0154777|T047|PT|360.40|ICD9CM|Degenerated globe or eye, unspecified|Degenerated globe or eye, unspecified
C0154777|T047|AB|360.40|ICD9CM|Degeneration of eye NOS|Degeneration of eye NOS
C0154788|T047|AB|360.41|ICD9CM|Blind hypotensive eye|Blind hypotensive eye
C0154788|T047|PT|360.41|ICD9CM|Blind hypotensive eye|Blind hypotensive eye
C0154789|T047|AB|360.42|ICD9CM|Blind hypertensive eye|Blind hypertensive eye
C0154789|T047|PT|360.42|ICD9CM|Blind hypertensive eye|Blind hypertensive eye
C1576412|T046|AB|360.43|ICD9CM|Hemophthalmos|Hemophthalmos
C1576412|T046|PT|360.43|ICD9CM|Hemophthalmos, except current injury|Hemophthalmos, except current injury
C0152458|T047|AB|360.44|ICD9CM|Leucocoria|Leucocoria
C0152458|T047|PT|360.44|ICD9CM|Leucocoria|Leucocoria
C0271008|T046|HT|360.5|ICD9CM|Retained (old) intraocular foreign body, magnetic|Retained (old) intraocular foreign body, magnetic
C0271008|T046|PT|360.50|ICD9CM|Foreign body, magnetic, intraocular, unspecified|Foreign body, magnetic, intraocular, unspecified
C0271008|T046|AB|360.50|ICD9CM|Old magnet fb, eye NOS|Old magnet fb, eye NOS
C0154792|T047|PT|360.51|ICD9CM|Foreign body, magnetic, in anterior chamber of eye|Foreign body, magnetic, in anterior chamber of eye
C0154792|T047|AB|360.51|ICD9CM|Old magnet fb, ant chamb|Old magnet fb, ant chamb
C0154793|T047|PT|360.52|ICD9CM|Foreign body, magnetic, in iris or ciliary body|Foreign body, magnetic, in iris or ciliary body
C0154793|T047|AB|360.52|ICD9CM|Old magnet fb, iris|Old magnet fb, iris
C0154794|T037|PT|360.53|ICD9CM|Foreign body, magnetic, in lens|Foreign body, magnetic, in lens
C0154794|T037|AB|360.53|ICD9CM|Old magnet fb, lens|Old magnet fb, lens
C0154795|T037|PT|360.54|ICD9CM|Foreign body, magnetic, in vitreous|Foreign body, magnetic, in vitreous
C0154795|T037|AB|360.54|ICD9CM|Old magnet fb, vitreous|Old magnet fb, vitreous
C0154796|T047|PT|360.55|ICD9CM|Foreign body, magnetic, in posterior wall|Foreign body, magnetic, in posterior wall
C0154796|T047|AB|360.55|ICD9CM|Old magnet fb, post wall|Old magnet fb, post wall
C0154797|T047|PT|360.59|ICD9CM|Intraocular foreign body, magnetic, in other or multiple sites|Intraocular foreign body, magnetic, in other or multiple sites
C0154797|T047|AB|360.59|ICD9CM|Old magnet fb, eye NEC|Old magnet fb, eye NEC
C0271015|T046|HT|360.6|ICD9CM|Retained (old) intraocular foreign body, nonmagnetic|Retained (old) intraocular foreign body, nonmagnetic
C0015401|T037|PT|360.60|ICD9CM|Foreign body, intraocular, unspecified|Foreign body, intraocular, unspecified
C0015401|T037|AB|360.60|ICD9CM|Intraocular FB NOS|Intraocular FB NOS
C0154799|T037|AB|360.61|ICD9CM|FB in anterior chamber|FB in anterior chamber
C0154799|T037|PT|360.61|ICD9CM|Foreign body in anterior chamber|Foreign body in anterior chamber
C0154800|T047|AB|360.62|ICD9CM|FB in iris or ciliary|FB in iris or ciliary
C0154800|T047|PT|360.62|ICD9CM|Foreign body in iris or ciliary body|Foreign body in iris or ciliary body
C0154801|T037|AB|360.63|ICD9CM|Foreign body in lens|Foreign body in lens
C0154801|T037|PT|360.63|ICD9CM|Foreign body in lens|Foreign body in lens
C0154802|T037|AB|360.64|ICD9CM|Foreign body in vitreous|Foreign body in vitreous
C0154802|T037|PT|360.64|ICD9CM|Foreign body in vitreous|Foreign body in vitreous
C0154803|T037|AB|360.65|ICD9CM|FB in posterior wall|FB in posterior wall
C0154803|T037|PT|360.65|ICD9CM|Foreign body in posterior wall of eye|Foreign body in posterior wall of eye
C0154804|T047|AB|360.69|ICD9CM|Intraocular FB NEC|Intraocular FB NEC
C0154804|T047|PT|360.69|ICD9CM|Intraocular foreign body in other or multiple sites|Intraocular foreign body in other or multiple sites
C0154805|T047|HT|360.8|ICD9CM|Other disorders of globe|Other disorders of globe
C0154806|T047|AB|360.81|ICD9CM|Luxation of globe|Luxation of globe
C0154806|T047|PT|360.81|ICD9CM|Luxation of globe|Luxation of globe
C0154805|T047|AB|360.89|ICD9CM|Disorder of globe NEC|Disorder of globe NEC
C0154805|T047|PT|360.89|ICD9CM|Other disorders of globe|Other disorders of globe
C0015397|T047|AB|360.9|ICD9CM|Disorder of globe NOS|Disorder of globe NOS
C0015397|T047|PT|360.9|ICD9CM|Unspecified disorder of globe|Unspecified disorder of globe
C1533659|T047|HT|361|ICD9CM|Retinal detachments and defects|Retinal detachments and defects
C0154808|T047|HT|361.0|ICD9CM|Retinal detachment with retinal defect|Retinal detachment with retinal defect
C0154808|T047|AB|361.00|ICD9CM|Detachmnt w defect NOS|Detachmnt w defect NOS
C0154808|T047|PT|361.00|ICD9CM|Retinal detachment with retinal defect, unspecified|Retinal detachment with retinal defect, unspecified
C0154809|T047|AB|361.01|ICD9CM|Part detach-singl defec|Part detach-singl defec
C0154809|T047|PT|361.01|ICD9CM|Recent retinal detachment, partial, with single defect|Recent retinal detachment, partial, with single defect
C0154810|T047|AB|361.02|ICD9CM|Part detach-mult defect|Part detach-mult defect
C0154810|T047|PT|361.02|ICD9CM|Recent retinal detachment, partial, with multiple defects|Recent retinal detachment, partial, with multiple defects
C0154811|T047|AB|361.03|ICD9CM|Part detach-giant tear|Part detach-giant tear
C0154811|T047|PT|361.03|ICD9CM|Recent retinal detachment, partial, with giant tear|Recent retinal detachment, partial, with giant tear
C0154812|T047|AB|361.04|ICD9CM|Part detach-dialysis|Part detach-dialysis
C0154812|T047|PT|361.04|ICD9CM|Recent retinal detachment, partial, with retinal dialysis|Recent retinal detachment, partial, with retinal dialysis
C0154813|T047|AB|361.05|ICD9CM|Recent detachment, total|Recent detachment, total
C0154813|T047|PT|361.05|ICD9CM|Recent retinal detachment, total or subtotal|Recent retinal detachment, total or subtotal
C0154814|T047|AB|361.06|ICD9CM|Old detachment, partial|Old detachment, partial
C0154814|T047|PT|361.06|ICD9CM|Old retinal detachment, partial|Old retinal detachment, partial
C0154815|T047|AB|361.07|ICD9CM|Old detachment, total|Old detachment, total
C0154815|T047|PT|361.07|ICD9CM|Old retinal detachment, total or subtotal|Old retinal detachment, total or subtotal
C0154816|T020|HT|361.1|ICD9CM|Retinoschisis and retinal cysts|Retinoschisis and retinal cysts
C0152439|T047|AB|361.10|ICD9CM|Retinoschisis NOS|Retinoschisis NOS
C0152439|T047|PT|361.10|ICD9CM|Retinoschisis, unspecified|Retinoschisis, unspecified
C0154817|T047|AB|361.11|ICD9CM|Flat retinoschisis|Flat retinoschisis
C0154817|T047|PT|361.11|ICD9CM|Flat retinoschisis|Flat retinoschisis
C0344289|T047|AB|361.12|ICD9CM|Bullous retinoschisis|Bullous retinoschisis
C0344289|T047|PT|361.12|ICD9CM|Bullous retinoschisis|Bullous retinoschisis
C0154819|T047|AB|361.13|ICD9CM|Primary retinal cysts|Primary retinal cysts
C0154819|T047|PT|361.13|ICD9CM|Primary retinal cysts|Primary retinal cysts
C0154820|T047|AB|361.14|ICD9CM|Secondary retinal cysts|Secondary retinal cysts
C0154820|T047|PT|361.14|ICD9CM|Secondary retinal cysts|Secondary retinal cysts
C0154821|T047|PT|361.19|ICD9CM|Other retinoschisis and retinal cysts|Other retinoschisis and retinal cysts
C0154821|T047|AB|361.19|ICD9CM|Retinoshisis or cyst NEC|Retinoshisis or cyst NEC
C0154822|T047|AB|361.2|ICD9CM|Serous retina detachment|Serous retina detachment
C0154822|T047|PT|361.2|ICD9CM|Serous retinal detachment|Serous retinal detachment
C0700508|T047|HT|361.3|ICD9CM|Retinal defects without detachment|Retinal defects without detachment
C0154823|T190|AB|361.30|ICD9CM|Retinal defect NOS|Retinal defect NOS
C0154823|T190|PT|361.30|ICD9CM|Retinal defect, unspecified|Retinal defect, unspecified
C0154825|T047|AB|361.31|ICD9CM|Round hole of retina|Round hole of retina
C0154825|T047|PT|361.31|ICD9CM|Round hole of retina without detachment|Round hole of retina without detachment
C0154826|T047|AB|361.32|ICD9CM|Horseshoe tear of retina|Horseshoe tear of retina
C0154826|T047|PT|361.32|ICD9CM|Horseshoe tear of retina without detachment|Horseshoe tear of retina without detachment
C0154827|T047|AB|361.33|ICD9CM|Mult defects of retina|Mult defects of retina
C0154827|T047|PT|361.33|ICD9CM|Multiple defects of retina without detachment|Multiple defects of retina without detachment
C0339440|T020|HT|361.8|ICD9CM|Other forms of retinal detachment|Other forms of retinal detachment
C0154828|T046|AB|361.81|ICD9CM|Retinal traction detach|Retinal traction detach
C0154828|T046|PT|361.81|ICD9CM|Traction detachment of retina|Traction detachment of retina
C0339440|T020|PT|361.89|ICD9CM|Other forms of retinal detachment|Other forms of retinal detachment
C0339440|T020|AB|361.89|ICD9CM|Retinal detachment NEC|Retinal detachment NEC
C0035305|T047|AB|361.9|ICD9CM|Retinal detachment NOS|Retinal detachment NOS
C0035305|T047|PT|361.9|ICD9CM|Unspecified retinal detachment|Unspecified retinal detachment
C0339438|T047|HT|362|ICD9CM|Other retinal disorders|Other retinal disorders
C0011884|T047|HT|362.0|ICD9CM|Diabetic retinopathy|Diabetic retinopathy
C0004606|T047|PT|362.01|ICD9CM|Background diabetic retinopathy|Background diabetic retinopathy
C0004606|T047|AB|362.01|ICD9CM|Diabetic retinopathy NOS|Diabetic retinopathy NOS
C0154830|T047|AB|362.02|ICD9CM|Prolif diab retinopathy|Prolif diab retinopathy
C0154830|T047|PT|362.02|ICD9CM|Proliferative diabetic retinopathy|Proliferative diabetic retinopathy
C0004606|T047|AB|362.03|ICD9CM|Nonprolf db retnoph NOS|Nonprolf db retnoph NOS
C0004606|T047|PT|362.03|ICD9CM|Nonproliferative diabetic retinopathy NOS|Nonproliferative diabetic retinopathy NOS
C0730276|T047|AB|362.04|ICD9CM|Mild nonprolf db retnoph|Mild nonprolf db retnoph
C0730276|T047|PT|362.04|ICD9CM|Mild nonproliferative diabetic retinopathy|Mild nonproliferative diabetic retinopathy
C0730277|T047|AB|362.05|ICD9CM|Mod nonprolf db retinoph|Mod nonprolf db retinoph
C0730277|T047|PT|362.05|ICD9CM|Moderate nonproliferative diabetic retinopathy|Moderate nonproliferative diabetic retinopathy
C0730278|T047|AB|362.06|ICD9CM|Sev nonprolf db retinoph|Sev nonprolf db retinoph
C0730278|T047|PT|362.06|ICD9CM|Severe nonproliferative diabetic retinopathy|Severe nonproliferative diabetic retinopathy
C0730285|T047|AB|362.07|ICD9CM|Diabetic macular edema|Diabetic macular edema
C0730285|T047|PT|362.07|ICD9CM|Diabetic macular edema|Diabetic macular edema
C0154831|T047|HT|362.1|ICD9CM|Other background retinopathy and retinal vascular changes|Other background retinopathy and retinal vascular changes
C0004608|T047|AB|362.10|ICD9CM|Backgrnd retinopathy NOS|Backgrnd retinopathy NOS
C0004608|T047|PT|362.10|ICD9CM|Background retinopathy, unspecified|Background retinopathy, unspecified
C0152132|T047|AB|362.11|ICD9CM|Hypertensive retinopathy|Hypertensive retinopathy
C0152132|T047|PT|362.11|ICD9CM|Hypertensive retinopathy|Hypertensive retinopathy
C0154832|T047|AB|362.12|ICD9CM|Exudative retinopathy|Exudative retinopathy
C0154832|T047|PT|362.12|ICD9CM|Exudative retinopathy|Exudative retinopathy
C1363843|T047|PT|362.13|ICD9CM|Changes in vascular appearance of retina|Changes in vascular appearance of retina
C1363843|T047|AB|362.13|ICD9CM|Retinal vascular changes|Retinal vascular changes
C0154834|T047|AB|362.14|ICD9CM|Retina microaneurysm NOS|Retina microaneurysm NOS
C0154834|T047|PT|362.14|ICD9CM|Retinal microaneurysms NOS|Retinal microaneurysms NOS
C0154835|T047|AB|362.15|ICD9CM|Retinal telangiectasia|Retinal telangiectasia
C0154835|T047|PT|362.15|ICD9CM|Retinal telangiectasia|Retinal telangiectasia
C0035320|T046|AB|362.16|ICD9CM|Retinal neovascular NOS|Retinal neovascular NOS
C0035320|T046|PT|362.16|ICD9CM|Retinal neovascularization NOS|Retinal neovascularization NOS
C0154836|T047|PT|362.17|ICD9CM|Other intraretinal microvascular abnormalities|Other intraretinal microvascular abnormalities
C0154836|T047|AB|362.17|ICD9CM|Retinal varices|Retinal varices
C0152026|T047|AB|362.18|ICD9CM|Retinal vasculitis|Retinal vasculitis
C0152026|T047|PT|362.18|ICD9CM|Retinal vasculitis|Retinal vasculitis
C0154837|T047|HT|362.2|ICD9CM|Other proliferative retinopathy|Other proliferative retinopathy
C0035344|T047|PT|362.20|ICD9CM|Retinopathy of prematurity, unspecified|Retinopathy of prematurity, unspecified
C0035344|T047|AB|362.20|ICD9CM|Retinoph prematurity NOS|Retinoph prematurity NOS
C0035344|T047|AB|362.21|ICD9CM|Retrolental fibroplasia|Retrolental fibroplasia
C0035344|T047|PT|362.21|ICD9CM|Retrolental fibroplasia|Retrolental fibroplasia
C3812410|T047|PT|362.22|ICD9CM|Retinopathy of prematurity, stage 0|Retinopathy of prematurity, stage 0
C3812410|T047|AB|362.22|ICD9CM|Retinoph prematr,stage 0|Retinoph prematr,stage 0
C1443381|T047|PT|362.23|ICD9CM|Retinopathy of prematurity, stage 1|Retinopathy of prematurity, stage 1
C1443381|T047|AB|362.23|ICD9CM|Retinoph prematr,stage 1|Retinoph prematr,stage 1
C1443382|T047|PT|362.24|ICD9CM|Retinopathy of prematurity, stage 2|Retinopathy of prematurity, stage 2
C1443382|T047|AB|362.24|ICD9CM|Retinoph prematr,stage 2|Retinoph prematr,stage 2
C1443383|T047|PT|362.25|ICD9CM|Retinopathy of prematurity, stage 3|Retinopathy of prematurity, stage 3
C1443383|T047|AB|362.25|ICD9CM|Retinoph prematr,stage 3|Retinoph prematr,stage 3
C1443384|T047|PT|362.26|ICD9CM|Retinopathy of prematurity, stage 4|Retinopathy of prematurity, stage 4
C1443384|T047|AB|362.26|ICD9CM|Retinoph prematr.stage 4|Retinoph prematr.stage 4
C1443385|T047|PT|362.27|ICD9CM|Retinopathy of prematurity, stage 5|Retinopathy of prematurity, stage 5
C1443385|T047|AB|362.27|ICD9CM|Retinoph prematr,stage 5|Retinoph prematr,stage 5
C0154838|T047|PT|362.29|ICD9CM|Other nondiabetic proliferative retinopathy|Other nondiabetic proliferative retinopathy
C0154838|T047|AB|362.29|ICD9CM|Prolif retinopathy NEC|Prolif retinopathy NEC
C0035326|T047|HT|362.3|ICD9CM|Retinal vascular occlusion|Retinal vascular occlusion
C0035326|T047|AB|362.30|ICD9CM|Retinal vasc occlus NOS|Retinal vasc occlus NOS
C0035326|T047|PT|362.30|ICD9CM|Retinal vascular occlusion, unspecified|Retinal vascular occlusion, unspecified
C0007688|T047|AB|362.31|ICD9CM|Cent retina artery occlu|Cent retina artery occlu
C0007688|T047|PT|362.31|ICD9CM|Central retinal artery occlusion|Central retinal artery occlusion
C0006123|T047|AB|362.32|ICD9CM|Arterial branch occlus|Arterial branch occlus
C0006123|T047|PT|362.32|ICD9CM|Retinal arterial branch occlusion|Retinal arterial branch occlusion
C0154839|T047|AB|362.33|ICD9CM|Part arterial occlusion|Part arterial occlusion
C0154839|T047|PT|362.33|ICD9CM|Partial retinal arterial occlusion|Partial retinal arterial occlusion
C0154840|T047|AB|362.34|ICD9CM|Transient arterial occlu|Transient arterial occlu
C0154840|T047|PT|362.34|ICD9CM|Transient retinal arterial occlusion|Transient retinal arterial occlusion
C0154841|T047|AB|362.35|ICD9CM|Cent retinal vein occlus|Cent retinal vein occlus
C0154841|T047|PT|362.35|ICD9CM|Central retinal vein occlusion|Central retinal vein occlusion
C0154842|T047|PT|362.36|ICD9CM|Venous tributary (branch) occlusion|Venous tributary (branch) occlusion
C0154842|T047|AB|362.36|ICD9CM|Venous tributary occlus|Venous tributary occlus
C0154843|T046|AB|362.37|ICD9CM|Retina venous engorgemnt|Retina venous engorgemnt
C0154843|T046|PT|362.37|ICD9CM|Venous engorgement|Venous engorgement
C0154844|T020|HT|362.4|ICD9CM|Separation of retinal layers|Separation of retinal layers
C0154844|T020|AB|362.40|ICD9CM|Retina layer separat NOS|Retina layer separat NOS
C0154844|T020|PT|362.40|ICD9CM|Retinal layer separation, unspecified|Retinal layer separation, unspecified
C0730328|T047|AB|362.41|ICD9CM|Cent serous retinopathy|Cent serous retinopathy
C0730328|T047|PT|362.41|ICD9CM|Central serous retinopathy|Central serous retinopathy
C0154845|T047|AB|362.42|ICD9CM|Serous detach pigm epith|Serous detach pigm epith
C0154845|T047|PT|362.42|ICD9CM|Serous detachment of retinal pigment epithelium|Serous detachment of retinal pigment epithelium
C0154846|T046|AB|362.43|ICD9CM|Hem detach pigmnt epith|Hem detach pigmnt epith
C0154846|T046|PT|362.43|ICD9CM|Hemorrhagic detachment of retinal pigment epithelium|Hemorrhagic detachment of retinal pigment epithelium
C0339436|T047|HT|362.5|ICD9CM|Degeneration of macula and posterior pole of retina|Degeneration of macula and posterior pole of retina
C0242383|T047|PT|362.50|ICD9CM|Macular degeneration (senile), unspecified|Macular degeneration (senile), unspecified
C0242383|T047|AB|362.50|ICD9CM|Macular degeneration NOS|Macular degeneration NOS
C0271083|T020|AB|362.51|ICD9CM|Nonexudat macular degen|Nonexudat macular degen
C0271083|T020|PT|362.51|ICD9CM|Nonexudative senile macular degeneration|Nonexudative senile macular degeneration
C0271084|T047|AB|362.52|ICD9CM|Exudative macular degen|Exudative macular degen
C0271084|T047|PT|362.52|ICD9CM|Exudative senile macular degeneration|Exudative senile macular degeneration
C0154850|T047|AB|362.53|ICD9CM|Cystoid macular degen|Cystoid macular degen
C0154850|T047|PT|362.53|ICD9CM|Cystoid macular degeneration|Cystoid macular degeneration
C1261331|T047|AB|362.54|ICD9CM|Macular cyst or hole|Macular cyst or hole
C1261331|T047|PT|362.54|ICD9CM|Macular cyst, hole, or pseudohole|Macular cyst, hole, or pseudohole
C0271086|T047|AB|362.55|ICD9CM|Toxic maculopathy|Toxic maculopathy
C0271086|T047|PT|362.55|ICD9CM|Toxic maculopathy|Toxic maculopathy
C0339543|T020|AB|362.56|ICD9CM|Macular puckering|Macular puckering
C0339543|T020|PT|362.56|ICD9CM|Macular puckering|Macular puckering
C0035312|T047|AB|362.57|ICD9CM|Drusen (degenerative)|Drusen (degenerative)
C0035312|T047|PT|362.57|ICD9CM|Drusen (degenerative)|Drusen (degenerative)
C1320640|T047|HT|362.6|ICD9CM|Peripheral retinal degenerations|Peripheral retinal degenerations
C1320640|T047|AB|362.60|ICD9CM|Periph retina degen NOS|Periph retina degen NOS
C1320640|T047|PT|362.60|ICD9CM|Peripheral retinal degeneration, unspecified|Peripheral retinal degeneration, unspecified
C0154854|T047|AB|362.61|ICD9CM|Paving stone degenerat|Paving stone degenerat
C0154854|T047|PT|362.61|ICD9CM|Paving stone degeneration|Paving stone degeneration
C0154855|T047|AB|362.62|ICD9CM|Microcystoid degenerat|Microcystoid degenerat
C0154855|T047|PT|362.62|ICD9CM|Microcystoid degeneration|Microcystoid degeneration
C0154856|T047|AB|362.63|ICD9CM|Lattice degeneration|Lattice degeneration
C0154856|T047|PT|362.63|ICD9CM|Lattice degeneration|Lattice degeneration
C0154857|T047|AB|362.64|ICD9CM|Senile reticular degen|Senile reticular degen
C0154857|T047|PT|362.64|ICD9CM|Senile reticular degeneration|Senile reticular degeneration
C0154858|T047|PT|362.65|ICD9CM|Secondary pigmentary degeneration|Secondary pigmentary degeneration
C0154858|T047|AB|362.65|ICD9CM|Secondry pigment degen|Secondry pigment degen
C0154859|T047|AB|362.66|ICD9CM|Sec vitreoretina degen|Sec vitreoretina degen
C0154859|T047|PT|362.66|ICD9CM|Secondary vitreoretinal degenerations|Secondary vitreoretinal degenerations
C0154860|T047|HT|362.7|ICD9CM|Hereditary retinal dystrophies|Hereditary retinal dystrophies
C0154860|T047|AB|362.70|ICD9CM|Hered retin dystrphy NOS|Hered retin dystrphy NOS
C0154860|T047|PT|362.70|ICD9CM|Hereditary retinal dystrophy, unspecified|Hereditary retinal dystrophy, unspecified
C0154861|T047|AB|362.71|ICD9CM|Ret dystrph in lipidoses|Ret dystrph in lipidoses
C0154861|T047|PT|362.71|ICD9CM|Retinal dystrophy in systemic or cerebroretinal lipidoses|Retinal dystrophy in systemic or cerebroretinal lipidoses
C0154862|T047|AB|362.72|ICD9CM|Ret dystrph in syst dis|Ret dystrph in syst dis
C0154862|T047|PT|362.72|ICD9CM|Retinal dystrophy in other systemic disorders and syndromes|Retinal dystrophy in other systemic disorders and syndromes
C0154863|T047|PT|362.73|ICD9CM|Vitreoretinal dystrophies|Vitreoretinal dystrophies
C0154863|T047|AB|362.73|ICD9CM|Vitreoretinal dystrophy|Vitreoretinal dystrophy
C4551633|T047|AB|362.74|ICD9CM|Pigment retina dystrophy|Pigment retina dystrophy
C4551633|T047|PT|362.74|ICD9CM|Pigmentary retinal dystrophy|Pigmentary retinal dystrophy
C0154864|T047|PT|362.75|ICD9CM|Other dystrophies primarily involving the sensory retina|Other dystrophies primarily involving the sensory retina
C0154864|T047|AB|362.75|ICD9CM|Sensory retina dystrophy|Sensory retina dystrophy
C0154865|T047|PT|362.76|ICD9CM|Dystrophies primarily involving the retinal pigment epithelium|Dystrophies primarily involving the retinal pigment epithelium
C0154865|T047|AB|362.76|ICD9CM|Vitelliform dystrophy|Vitelliform dystrophy
C0154866|T047|AB|362.77|ICD9CM|Bruch membrane dystrophy|Bruch membrane dystrophy
C0154866|T047|PT|362.77|ICD9CM|Dystrophies primarily involving Bruch's membrane|Dystrophies primarily involving Bruch's membrane
C0339438|T047|HT|362.8|ICD9CM|Other retinal disorders|Other retinal disorders
C0035317|T047|AB|362.81|ICD9CM|Retinal hemorrhage|Retinal hemorrhage
C0035317|T047|PT|362.81|ICD9CM|Retinal hemorrhage|Retinal hemorrhage
C0154867|T047|AB|362.82|ICD9CM|Retina exudates/deposits|Retina exudates/deposits
C0154867|T047|PT|362.82|ICD9CM|Retinal exudates and deposits|Retinal exudates and deposits
C0242420|T046|AB|362.83|ICD9CM|Retinal edema|Retinal edema
C0242420|T046|PT|362.83|ICD9CM|Retinal edema|Retinal edema
C0162291|T046|AB|362.84|ICD9CM|Retinal ischemia|Retinal ischemia
C0162291|T046|PT|362.84|ICD9CM|Retinal ischemia|Retinal ischemia
C0474334|T047|AB|362.85|ICD9CM|Retinal nerv fiber defec|Retinal nerv fiber defec
C0474334|T047|PT|362.85|ICD9CM|Retinal nerve fiber bundle defects|Retinal nerve fiber bundle defects
C0339438|T047|PT|362.89|ICD9CM|Other retinal disorders|Other retinal disorders
C0339438|T047|AB|362.89|ICD9CM|Retinal disorders NEC|Retinal disorders NEC
C0035309|T047|AB|362.9|ICD9CM|Retinal disorder NOS|Retinal disorder NOS
C0035309|T047|PT|362.9|ICD9CM|Unspecified retinal disorder|Unspecified retinal disorder
C0008511|T047|HT|363|ICD9CM|Chorioretinal inflammations, scars, and other disorders of choroid|Chorioretinal inflammations, scars, and other disorders of choroid
C0154870|T047|HT|363.0|ICD9CM|Focal chorioretinitis and focal retinochoroiditis|Focal chorioretinitis and focal retinochoroiditis
C0154870|T047|AB|363.00|ICD9CM|Focal chorioretinit NOS|Focal chorioretinit NOS
C0154870|T047|PT|363.00|ICD9CM|Focal chorioretinitis, unspecified|Focal chorioretinitis, unspecified
C0154871|T047|PT|363.01|ICD9CM|Focal choroiditis and chorioretinitis, juxtapapillary|Focal choroiditis and chorioretinitis, juxtapapillary
C0154871|T047|AB|363.01|ICD9CM|Juxtapap foc choroiditis|Juxtapap foc choroiditis
C0154872|T047|AB|363.03|ICD9CM|Foc choroiditis post NEC|Foc choroiditis post NEC
C0154872|T047|PT|363.03|ICD9CM|Focal choroiditis and chorioretinitis of other posterior pole|Focal choroiditis and chorioretinitis of other posterior pole
C0339394|T047|PT|363.04|ICD9CM|Focal choroiditis and chorioretinitis, peripheral|Focal choroiditis and chorioretinitis, peripheral
C0339394|T047|AB|363.04|ICD9CM|Periph focal choroiditis|Periph focal choroiditis
C3665438|T047|PT|363.05|ICD9CM|Focal retinitis and retinochoroiditis, juxtapapillary|Focal retinitis and retinochoroiditis, juxtapapillary
C3665438|T047|AB|363.05|ICD9CM|Juxtapap focal retinitis|Juxtapap focal retinitis
C0154875|T047|PT|363.06|ICD9CM|Focal retinitis and retinochoroiditis, macular or paramacular|Focal retinitis and retinochoroiditis, macular or paramacular
C0154875|T047|AB|363.06|ICD9CM|Macular focal retinitis|Macular focal retinitis
C0154876|T047|AB|363.07|ICD9CM|Foc retinitis post NEC|Foc retinitis post NEC
C0154876|T047|PT|363.07|ICD9CM|Focal retinitis and retinochoroiditis of other posterior pole|Focal retinitis and retinochoroiditis of other posterior pole
C0154877|T047|PT|363.08|ICD9CM|Focal retinitis and retinochoroiditis, peripheral|Focal retinitis and retinochoroiditis, peripheral
C0154877|T047|AB|363.08|ICD9CM|Periph focal retinitis|Periph focal retinitis
C0154879|T047|HT|363.1|ICD9CM|Disseminated chorioretinitis and disseminated retinochoroiditis|Disseminated chorioretinitis and disseminated retinochoroiditis
C0154879|T047|AB|363.10|ICD9CM|Dissem chorioretinit NOS|Dissem chorioretinit NOS
C0154879|T047|PT|363.10|ICD9CM|Disseminated chorioretinitis, unspecified|Disseminated chorioretinitis, unspecified
C0154880|T047|AB|363.11|ICD9CM|Dissem choroiditis, post|Dissem choroiditis, post
C0154880|T047|PT|363.11|ICD9CM|Disseminated choroiditis and chorioretinitis, posterior pole|Disseminated choroiditis and chorioretinitis, posterior pole
C0154881|T047|PT|363.12|ICD9CM|Disseminated choroiditis and chorioretinitis, peripheral|Disseminated choroiditis and chorioretinitis, peripheral
C0154881|T047|AB|363.12|ICD9CM|Periph disem choroiditis|Periph disem choroiditis
C0154882|T047|PT|363.13|ICD9CM|Disseminated choroiditis and chorioretinitis, generalized|Disseminated choroiditis and chorioretinitis, generalized
C0154882|T047|AB|363.13|ICD9CM|Gen dissem choroiditis|Gen dissem choroiditis
C0154883|T047|PT|363.14|ICD9CM|Disseminated retinitis and retinochoroiditis, metastatic|Disseminated retinitis and retinochoroiditis, metastatic
C0154883|T047|AB|363.14|ICD9CM|Metastat dissem retinit|Metastat dissem retinit
C0154884|T047|PT|363.15|ICD9CM|Disseminated retinitis and retinochoroiditis, pigment epitheliopathy|Disseminated retinitis and retinochoroiditis, pigment epitheliopathy
C0154884|T047|AB|363.15|ICD9CM|Pigment epitheliopathy|Pigment epitheliopathy
C2239106|T047|HT|363.2|ICD9CM|Other and unspecified forms of chorioretinitis and retinochoroiditis|Other and unspecified forms of chorioretinitis and retinochoroiditis
C0008513|T047|AB|363.20|ICD9CM|Chorioretinitis NOS|Chorioretinitis NOS
C0008513|T047|PT|363.20|ICD9CM|Chorioretinitis, unspecified|Chorioretinitis, unspecified
C0030593|T047|AB|363.21|ICD9CM|Pars planitis|Pars planitis
C0030593|T047|PT|363.21|ICD9CM|Pars planitis|Pars planitis
C0042170|T047|AB|363.22|ICD9CM|Harada's disease|Harada's disease
C0042170|T047|PT|363.22|ICD9CM|Harada's disease|Harada's disease
C0008512|T020|HT|363.3|ICD9CM|Chorioretinal scars|Chorioretinal scars
C0008512|T020|AB|363.30|ICD9CM|Chorioretinal scar NOS|Chorioretinal scar NOS
C0008512|T020|PT|363.30|ICD9CM|Chorioretinal scar, unspecified|Chorioretinal scar, unspecified
C0152131|T047|AB|363.31|ICD9CM|Solar retinopathy|Solar retinopathy
C0152131|T047|PT|363.31|ICD9CM|Solar retinopathy|Solar retinopathy
C0339418|T020|AB|363.32|ICD9CM|Macular scars NEC|Macular scars NEC
C0339418|T020|PT|363.32|ICD9CM|Other macular scars|Other macular scars
C0339419|T020|PT|363.33|ICD9CM|Other scars of posterior pole|Other scars of posterior pole
C0339419|T020|AB|363.33|ICD9CM|Posterior pole scar NEC|Posterior pole scar NEC
C0154888|T047|AB|363.34|ICD9CM|Peripheral retinal scars|Peripheral retinal scars
C0154888|T047|PT|363.34|ICD9CM|Peripheral scars|Peripheral scars
C0154889|T047|AB|363.35|ICD9CM|Disseminated retina scar|Disseminated retina scar
C0154889|T047|PT|363.35|ICD9CM|Disseminated scars|Disseminated scars
C0344297|T047|HT|363.4|ICD9CM|Choroidal degenerations|Choroidal degenerations
C0344297|T047|AB|363.40|ICD9CM|Choroidal degen NOS|Choroidal degen NOS
C0344297|T047|PT|363.40|ICD9CM|Choroidal degeneration, unspecified|Choroidal degeneration, unspecified
C0154891|T047|PT|363.41|ICD9CM|Senile atrophy of choroid|Senile atrophy of choroid
C0154891|T047|AB|363.41|ICD9CM|Senile atrophy, choroid|Senile atrophy, choroid
C0154892|T047|PT|363.42|ICD9CM|Diffuse secondary atrophy of choroid|Diffuse secondary atrophy of choroid
C0154892|T047|AB|363.42|ICD9CM|Difus sec atroph choroid|Difus sec atroph choroid
C0002983|T047|PT|363.43|ICD9CM|Angioid streaks of choroid|Angioid streaks of choroid
C0002983|T047|AB|363.43|ICD9CM|Angioid streaks, choroid|Angioid streaks, choroid
C0154893|T047|HT|363.5|ICD9CM|Hereditary choroidal dystrophies|Hereditary choroidal dystrophies
C0154893|T047|AB|363.50|ICD9CM|Hered choroid atroph NOS|Hered choroid atroph NOS
C0154893|T047|PT|363.50|ICD9CM|Hereditary choroidal dystrophy or atrophy, unspecified|Hereditary choroidal dystrophy or atrophy, unspecified
C0154895|T047|PT|363.51|ICD9CM|Circumpapillary dystrophy of choroid, partial|Circumpapillary dystrophy of choroid, partial
C0154895|T047|AB|363.51|ICD9CM|Prt circmpap choroid dys|Prt circmpap choroid dys
C0154896|T047|PT|363.52|ICD9CM|Circumpapillary dystrophy of choroid, total|Circumpapillary dystrophy of choroid, total
C0154896|T047|AB|363.52|ICD9CM|Tot circmpap choroid dys|Tot circmpap choroid dys
C0339427|T047|PT|363.53|ICD9CM|Central dystrophy of choroid, partial|Central dystrophy of choroid, partial
C0339427|T047|AB|363.53|ICD9CM|Part cent choroid dystr|Part cent choroid dystr
C0154898|T047|PT|363.54|ICD9CM|Central choroidal atrophy, total|Central choroidal atrophy, total
C0154898|T047|AB|363.54|ICD9CM|Tot cent choroid atrophy|Tot cent choroid atrophy
C0008525|T047|AB|363.55|ICD9CM|Choroideremia|Choroideremia
C0008525|T047|PT|363.55|ICD9CM|Choroideremia|Choroideremia
C0154899|T047|PT|363.56|ICD9CM|Other diffuse or generalized dystrophy of choroid, partial|Other diffuse or generalized dystrophy of choroid, partial
C0154899|T047|AB|363.56|ICD9CM|Prt gen choroid dyst NEC|Prt gen choroid dyst NEC
C0154900|T047|PT|363.57|ICD9CM|Other diffuse or generalized dystrophy of choroid, total|Other diffuse or generalized dystrophy of choroid, total
C0154900|T047|AB|363.57|ICD9CM|Tot gen choroid dyst NEC|Tot gen choroid dyst NEC
C0154901|T046|HT|363.6|ICD9CM|Choroidal hemorrhage and rupture|Choroidal hemorrhage and rupture
C0008522|T046|AB|363.61|ICD9CM|Choroidal hemorrhage NOS|Choroidal hemorrhage NOS
C0008522|T046|PT|363.61|ICD9CM|Choroidal hemorrhage, unspecified|Choroidal hemorrhage, unspecified
C0154902|T047|AB|363.62|ICD9CM|Expulsive choroid hemorr|Expulsive choroid hemorr
C0154902|T047|PT|363.62|ICD9CM|Expulsive choroidal hemorrhage|Expulsive choroidal hemorrhage
C0154903|T047|AB|363.63|ICD9CM|Choroidal rupture|Choroidal rupture
C0154903|T047|PT|363.63|ICD9CM|Choroidal rupture|Choroidal rupture
C0162279|T020|HT|363.7|ICD9CM|Choroidal detachment|Choroidal detachment
C0162279|T020|AB|363.70|ICD9CM|Choroidal detachment NOS|Choroidal detachment NOS
C0162279|T020|PT|363.70|ICD9CM|Choroidal detachment, unspecified|Choroidal detachment, unspecified
C0154904|T047|AB|363.71|ICD9CM|Serous choroid detachmnt|Serous choroid detachmnt
C0154904|T047|PT|363.71|ICD9CM|Serous choroidal detachment|Serous choroidal detachment
C0154905|T047|AB|363.72|ICD9CM|Hemorr choroid detachmnt|Hemorr choroid detachmnt
C0154905|T047|PT|363.72|ICD9CM|Hemorrhagic choroidal detachment|Hemorrhagic choroidal detachment
C0154906|T047|AB|363.8|ICD9CM|Disorders of choroid NEC|Disorders of choroid NEC
C0154906|T047|PT|363.8|ICD9CM|Other disorders of choroid|Other disorders of choroid
C0008521|T047|AB|363.9|ICD9CM|Choroidal disorder NOS|Choroidal disorder NOS
C0008521|T047|PT|363.9|ICD9CM|Unspecified disorder of choroid|Unspecified disorder of choroid
C0154907|T047|HT|364|ICD9CM|Disorders of iris and ciliary body|Disorders of iris and ciliary body
C0154908|T047|HT|364.0|ICD9CM|Acute and subacute iridocyclitis|Acute and subacute iridocyclitis
C0154908|T047|PT|364.00|ICD9CM|Acute and subacute iridocyclitis, unspecified|Acute and subacute iridocyclitis, unspecified
C0154908|T047|AB|364.00|ICD9CM|Acute iridocyclitis NOS|Acute iridocyclitis NOS
C0154909|T047|AB|364.01|ICD9CM|Primary iridocyclitis|Primary iridocyclitis
C0154909|T047|PT|364.01|ICD9CM|Primary iridocyclitis|Primary iridocyclitis
C0154910|T047|AB|364.02|ICD9CM|Recurrent iridocyclitis|Recurrent iridocyclitis
C0154910|T047|PT|364.02|ICD9CM|Recurrent iridocyclitis|Recurrent iridocyclitis
C0154911|T047|PT|364.03|ICD9CM|Secondary iridocyclitis, infectious|Secondary iridocyclitis, infectious
C0154911|T047|AB|364.03|ICD9CM|Secondry iritis, infect|Secondry iritis, infect
C2937264|T047|AB|364.04|ICD9CM|Second iritis, noninfec|Second iritis, noninfec
C2937264|T047|PT|364.04|ICD9CM|Secondary iridocyclitis, noninfectious|Secondary iridocyclitis, noninfectious
C0020641|T047|AB|364.05|ICD9CM|Hypopyon|Hypopyon
C0020641|T047|PT|364.05|ICD9CM|Hypopyon|Hypopyon
C1510449|T047|HT|364.1|ICD9CM|Chronic iridocyclitis|Chronic iridocyclitis
C1510449|T047|AB|364.10|ICD9CM|Chr iridocyclitis NOS|Chr iridocyclitis NOS
C1510449|T047|PT|364.10|ICD9CM|Chronic iridocyclitis, unspecified|Chronic iridocyclitis, unspecified
C0339319|T047|AB|364.11|ICD9CM|Chr iridocyl in oth dis|Chr iridocyl in oth dis
C0339319|T047|PT|364.11|ICD9CM|Chronic iridocyclitis in diseases classified elsewhere|Chronic iridocyclitis in diseases classified elsewhere
C0007832|T047|HT|364.2|ICD9CM|Certain types of iridocyclitis|Certain types of iridocyclitis
C0016782|T047|AB|364.21|ICD9CM|Fuch hetrochrom cyclitis|Fuch hetrochrom cyclitis
C0016782|T047|PT|364.21|ICD9CM|Fuchs' heterochromic cyclitis|Fuchs' heterochromic cyclitis
C0152138|T047|AB|364.22|ICD9CM|Glaucomatocyclit crises|Glaucomatocyclit crises
C0152138|T047|PT|364.22|ICD9CM|Glaucomatocyclitic crises|Glaucomatocyclitic crises
C0339320|T047|AB|364.23|ICD9CM|Lens-induced iridocyclit|Lens-induced iridocyclit
C0339320|T047|PT|364.23|ICD9CM|Lens-induced iridocyclitis|Lens-induced iridocyclitis
C0042170|T047|AB|364.24|ICD9CM|Vogt-koyanagi syndrome|Vogt-koyanagi syndrome
C0042170|T047|PT|364.24|ICD9CM|Vogt-koyanagi syndrome|Vogt-koyanagi syndrome
C0022073|T047|AB|364.3|ICD9CM|Iridocyclitis NOS|Iridocyclitis NOS
C0022073|T047|PT|364.3|ICD9CM|Unspecified iridocyclitis|Unspecified iridocyclitis
C0154915|T047|HT|364.4|ICD9CM|Vascular disorders of iris and ciliary body|Vascular disorders of iris and ciliary body
C0020582|T047|AB|364.41|ICD9CM|Hyphema|Hyphema
C0020582|T047|PT|364.41|ICD9CM|Hyphema of iris and ciliary body|Hyphema of iris and ciliary body
C0154916|T047|AB|364.42|ICD9CM|Rubeosis iridis|Rubeosis iridis
C0154916|T047|PT|364.42|ICD9CM|Rubeosis iridis|Rubeosis iridis
C0154917|T020|HT|364.5|ICD9CM|Degenerations of iris and ciliary body|Degenerations of iris and ciliary body
C0271111|T047|PT|364.51|ICD9CM|Essential or progressive iris atrophy|Essential or progressive iris atrophy
C0271111|T047|AB|364.51|ICD9CM|Progressive iris atrophy|Progressive iris atrophy
C0154919|T047|AB|364.52|ICD9CM|Iridoschisis|Iridoschisis
C0154919|T047|PT|364.52|ICD9CM|Iridoschisis|Iridoschisis
C0154920|T033|AB|364.53|ICD9CM|Pigment iris degenerat|Pigment iris degenerat
C0154920|T033|PT|364.53|ICD9CM|Pigmentary iris degeneration|Pigmentary iris degeneration
C0154921|T047|PT|364.54|ICD9CM|Degeneration of pupillary margin|Degeneration of pupillary margin
C0154921|T047|AB|364.54|ICD9CM|Pupillary margin degen|Pupillary margin degen
C0154922|T047|AB|364.55|ICD9CM|Miotic cyst pupil margin|Miotic cyst pupil margin
C0154922|T047|PT|364.55|ICD9CM|Miotic cysts of pupillary margin|Miotic cysts of pupillary margin
C0154923|T020|AB|364.56|ICD9CM|Degen chamber angle|Degen chamber angle
C0154923|T020|PT|364.56|ICD9CM|Degenerative changes of chamber angle|Degenerative changes of chamber angle
C0154924|T047|AB|364.57|ICD9CM|Degen ciliary body|Degen ciliary body
C0154924|T047|PT|364.57|ICD9CM|Degenerative changes of ciliary body|Degenerative changes of ciliary body
C0154925|T047|AB|364.59|ICD9CM|Iris atrophy NEC|Iris atrophy NEC
C0154925|T047|PT|364.59|ICD9CM|Other iris atrophy|Other iris atrophy
C0154926|T047|HT|364.6|ICD9CM|Cysts of iris, ciliary body, and anterior chamber|Cysts of iris, ciliary body, and anterior chamber
C0154927|T047|AB|364.60|ICD9CM|Idiopathic cysts|Idiopathic cysts
C0154927|T047|PT|364.60|ICD9CM|Idiopathic cysts of iris, ciliary body, and anterior chamber|Idiopathic cysts of iris, ciliary body, and anterior chamber
C0271128|T047|AB|364.61|ICD9CM|Implantation cysts|Implantation cysts
C0271128|T047|PT|364.61|ICD9CM|Implantation cysts of iris, ciliary body, and anterior chamber|Implantation cysts of iris, ciliary body, and anterior chamber
C0154929|T047|AB|364.62|ICD9CM|Exud cyst iris/ant chamb|Exud cyst iris/ant chamb
C0154929|T047|PT|364.62|ICD9CM|Exudative cysts of iris or anterior chamber|Exudative cysts of iris or anterior chamber
C0154930|T047|PT|364.63|ICD9CM|Primary cyst of pars plana|Primary cyst of pars plana
C0154930|T047|AB|364.63|ICD9CM|Primary cyst pars plana|Primary cyst pars plana
C0154931|T047|AB|364.64|ICD9CM|Exudat cyst pars plana|Exudat cyst pars plana
C0154931|T047|PT|364.64|ICD9CM|Exudative cyst of pars plana|Exudative cyst of pars plana
C0154932|T047|HT|364.7|ICD9CM|Adhesions and disruptions of iris and ciliary body|Adhesions and disruptions of iris and ciliary body
C0154933|T047|AB|364.70|ICD9CM|Adhesions of iris NOS|Adhesions of iris NOS
C0154933|T047|PT|364.70|ICD9CM|Adhesions of iris, unspecified|Adhesions of iris, unspecified
C0152253|T047|AB|364.71|ICD9CM|Posterior synechiae|Posterior synechiae
C0152253|T047|PT|364.71|ICD9CM|Posterior synechiae of iris|Posterior synechiae of iris
C0152252|T047|AB|364.72|ICD9CM|Anterior synechiae|Anterior synechiae
C0152252|T047|PT|364.72|ICD9CM|Anterior synechiae of iris|Anterior synechiae of iris
C0154934|T047|AB|364.73|ICD9CM|Goniosynechiae|Goniosynechiae
C0154934|T047|PT|364.73|ICD9CM|Goniosynechiae|Goniosynechiae
C0154935|T047|PT|364.74|ICD9CM|Adhesions and disruptions of pupillary membranes|Adhesions and disruptions of pupillary membranes
C0154935|T047|AB|364.74|ICD9CM|Pupillary membranes|Pupillary membranes
C0154936|T033|AB|364.75|ICD9CM|Pupillary abnormalities|Pupillary abnormalities
C0154936|T033|PT|364.75|ICD9CM|Pupillary abnormalities|Pupillary abnormalities
C0152246|T047|AB|364.76|ICD9CM|Iridodialysis|Iridodialysis
C0152246|T047|PT|364.76|ICD9CM|Iridodialysis|Iridodialysis
C0154937|T046|PT|364.77|ICD9CM|Recession of chamber angle of eye|Recession of chamber angle of eye
C0154937|T046|AB|364.77|ICD9CM|Recession, chamber angle|Recession, chamber angle
C0339308|T047|HT|364.8|ICD9CM|Other disorders of iris and ciliary body|Other disorders of iris and ciliary body
C1735601|T046|PT|364.81|ICD9CM|Floppy iris syndrome|Floppy iris syndrome
C1735601|T046|AB|364.81|ICD9CM|Floppy iris syndrome|Floppy iris syndrome
C1321345|T047|PT|364.82|ICD9CM|Plateau iris syndrome|Plateau iris syndrome
C1321345|T047|AB|364.82|ICD9CM|Plateau iris syndrome|Plateau iris syndrome
C0348538|T047|AB|364.89|ICD9CM|Iris/ciliary disord NEC|Iris/ciliary disord NEC
C0348538|T047|PT|364.89|ICD9CM|Other disorders of iris and ciliary body|Other disorders of iris and ciliary body
C0154907|T047|AB|364.9|ICD9CM|Iris/ciliary dis NOS|Iris/ciliary dis NOS
C0154907|T047|PT|364.9|ICD9CM|Unspecified disorder of iris and ciliary body|Unspecified disorder of iris and ciliary body
C0017601|T047|HT|365|ICD9CM|Glaucoma|Glaucoma
C1533674|T047|HT|365.0|ICD9CM|Borderline glaucoma [glaucoma suspect]|Borderline glaucoma [glaucoma suspect]
C0549470|T047|AB|365.00|ICD9CM|Preglaucoma NOS|Preglaucoma NOS
C0549470|T047|PT|365.00|ICD9CM|Preglaucoma, unspecified|Preglaucoma, unspecified
C3264152|T047|PT|365.01|ICD9CM|Open angle with borderline findings, low risk|Open angle with borderline findings, low risk
C3264152|T047|AB|365.01|ICD9CM|Opn angl brderln lo risk|Opn angl brderln lo risk
C0154941|T047|AB|365.02|ICD9CM|Anatomical narrow angle|Anatomical narrow angle
C0154941|T047|PT|365.02|ICD9CM|Anatomical narrow angle borderline glaucoma|Anatomical narrow angle borderline glaucoma
C0339572|T047|AB|365.03|ICD9CM|Steroid responders|Steroid responders
C0339572|T047|PT|365.03|ICD9CM|Steroid responders borderline glaucoma|Steroid responders borderline glaucoma
C0028840|T047|AB|365.04|ICD9CM|Ocular hypertension|Ocular hypertension
C0028840|T047|PT|365.04|ICD9CM|Ocular hypertension|Ocular hypertension
C3161083|T047|PT|365.05|ICD9CM|Open angle with borderline findings, high risk|Open angle with borderline findings, high risk
C3161083|T047|AB|365.05|ICD9CM|Opn ang w brdrlne hi rsk|Opn ang w brdrlne hi rsk
C3161084|T047|AB|365.06|ICD9CM|Prim angle clos w/o dmg|Prim angle clos w/o dmg
C3161084|T047|PT|365.06|ICD9CM|Primary angle closure without glaucoma damage|Primary angle closure without glaucoma damage
C0017612|T047|HT|365.1|ICD9CM|Open-angle glaucoma|Open-angle glaucoma
C0017612|T047|AB|365.10|ICD9CM|Open-angle glaucoma NOS|Open-angle glaucoma NOS
C0017612|T047|PT|365.10|ICD9CM|Open-angle glaucoma, unspecified|Open-angle glaucoma, unspecified
C0339573|T047|AB|365.11|ICD9CM|Prim open angle glaucoma|Prim open angle glaucoma
C0339573|T047|PT|365.11|ICD9CM|Primary open angle glaucoma|Primary open angle glaucoma
C0152136|T047|AB|365.12|ICD9CM|Low tension glaucoma|Low tension glaucoma
C0152136|T047|PT|365.12|ICD9CM|Low tension open-angle glaucoma|Low tension open-angle glaucoma
C0017612|T047|AB|365.13|ICD9CM|Pigmentary glaucoma|Pigmentary glaucoma
C0017612|T047|PT|365.13|ICD9CM|Pigmentary open-angle glaucoma|Pigmentary open-angle glaucoma
C2981140|T047|AB|365.14|ICD9CM|Glaucoma of childhood|Glaucoma of childhood
C2981140|T047|PT|365.14|ICD9CM|Glaucoma of childhood|Glaucoma of childhood
C0154944|T047|AB|365.15|ICD9CM|Residual opn ang glaucma|Residual opn ang glaucma
C0154944|T047|PT|365.15|ICD9CM|Residual stage of open angle glaucoma|Residual stage of open angle glaucoma
C0017606|T047|HT|365.2|ICD9CM|Primary angle-closure glaucoma|Primary angle-closure glaucoma
C0017606|T047|AB|365.20|ICD9CM|Prim angl-clos glauc NOS|Prim angl-clos glauc NOS
C0017606|T047|PT|365.20|ICD9CM|Primary angle-closure glaucoma, unspecified|Primary angle-closure glaucoma, unspecified
C0154945|T047|AB|365.21|ICD9CM|Intermit angl-clos glauc|Intermit angl-clos glauc
C0154945|T047|PT|365.21|ICD9CM|Intermittent angle-closure glaucoma|Intermittent angle-closure glaucoma
C0154946|T047|AB|365.22|ICD9CM|Acute angl-clos glaucoma|Acute angl-clos glaucoma
C0154946|T047|PT|365.22|ICD9CM|Acute angle-closure glaucoma|Acute angle-closure glaucoma
C0154947|T047|AB|365.23|ICD9CM|Chr angle-clos glaucoma|Chr angle-clos glaucoma
C0154947|T047|PT|365.23|ICD9CM|Chronic angle-closure glaucoma|Chronic angle-closure glaucoma
C0154948|T047|AB|365.24|ICD9CM|Residual angl-clos glauc|Residual angl-clos glauc
C0154948|T047|PT|365.24|ICD9CM|Residual stage of angle-closure glaucoma|Residual stage of angle-closure glaucoma
C0339578|T047|HT|365.3|ICD9CM|Corticosteroid-induced glaucoma|Corticosteroid-induced glaucoma
C0339579|T047|PT|365.31|ICD9CM|Corticosteroid-induced glaucoma, glaucomatous stage|Corticosteroid-induced glaucoma, glaucomatous stage
C0339579|T047|AB|365.31|ICD9CM|Glauc stage-ster induced|Glauc stage-ster induced
C0339580|T047|PT|365.32|ICD9CM|Corticosteroid-induced glaucoma, residual stage|Corticosteroid-induced glaucoma, residual stage
C0339580|T047|AB|365.32|ICD9CM|Glauc resid-ster induced|Glauc resid-ster induced
C0154952|T047|HT|365.4|ICD9CM|Glaucoma associated with congenital anomalies, dystrophies, and systemic syndromes|Glaucoma associated with congenital anomalies, dystrophies, and systemic syndromes
C0154953|T047|AB|365.41|ICD9CM|Glauc w chamb angle anom|Glauc w chamb angle anom
C0154953|T047|PT|365.41|ICD9CM|Glaucoma associated with chamber angle anomalies|Glaucoma associated with chamber angle anomalies
C0154954|T047|PT|365.42|ICD9CM|Glaucoma associated with anomalies of iris|Glaucoma associated with anomalies of iris
C0154954|T047|AB|365.42|ICD9CM|Glaucoma w iris anomaly|Glaucoma w iris anomaly
C0154955|T047|AB|365.43|ICD9CM|Glauc w ant seg anom NEC|Glauc w ant seg anom NEC
C0154955|T047|PT|365.43|ICD9CM|Glaucoma associated with other anterior segment anomalies|Glaucoma associated with other anterior segment anomalies
C0154956|T047|PT|365.44|ICD9CM|Glaucoma associated with systemic syndromes|Glaucoma associated with systemic syndromes
C0154956|T047|AB|365.44|ICD9CM|Glaucoma w systemic synd|Glaucoma w systemic synd
C0271142|T047|HT|365.5|ICD9CM|Glaucoma associated with disorders of the lens|Glaucoma associated with disorders of the lens
C0152137|T047|AB|365.51|ICD9CM|Phacolytic glaucoma|Phacolytic glaucoma
C0152137|T047|PT|365.51|ICD9CM|Phacolytic glaucoma|Phacolytic glaucoma
C0206368|T047|AB|365.52|ICD9CM|Pseudoexfoliat glaucoma|Pseudoexfoliat glaucoma
C0206368|T047|PT|365.52|ICD9CM|Pseudoexfoliation glaucoma|Pseudoexfoliation glaucoma
C0154959|T047|PT|365.59|ICD9CM|Glaucoma associated with other lens disorders|Glaucoma associated with other lens disorders
C0154959|T047|AB|365.59|ICD9CM|Glaucoma w lens dis NEC|Glaucoma w lens dis NEC
C0154960|T047|HT|365.6|ICD9CM|Glaucoma associated with other ocular disorders|Glaucoma associated with other ocular disorders
C0154961|T047|AB|365.60|ICD9CM|Glauc w ocular dis NOS|Glauc w ocular dis NOS
C0154961|T047|PT|365.60|ICD9CM|Glaucoma associated with unspecified ocular disorder|Glaucoma associated with unspecified ocular disorder
C0339598|T047|AB|365.61|ICD9CM|Glauc w pupillary block|Glauc w pupillary block
C0339598|T047|PT|365.61|ICD9CM|Glaucoma associated with pupillary block|Glaucoma associated with pupillary block
C0339593|T047|PT|365.62|ICD9CM|Glaucoma associated with ocular inflammations|Glaucoma associated with ocular inflammations
C0339593|T047|AB|365.62|ICD9CM|Glaucoma w ocular inflam|Glaucoma w ocular inflam
C0154964|T047|PT|365.63|ICD9CM|Glaucoma associated with vascular disorders|Glaucoma associated with vascular disorders
C0154964|T047|AB|365.63|ICD9CM|Glaucoma w vascular dis|Glaucoma w vascular dis
C0154965|T047|PT|365.64|ICD9CM|Glaucoma associated with tumors or cysts|Glaucoma associated with tumors or cysts
C0154965|T047|AB|365.64|ICD9CM|Glaucoma w tumor or cyst|Glaucoma w tumor or cyst
C0339594|T047|PT|365.65|ICD9CM|Glaucoma associated with ocular trauma|Glaucoma associated with ocular trauma
C0339594|T047|AB|365.65|ICD9CM|Glaucoma w ocular trauma|Glaucoma w ocular trauma
C3161085|T033|HT|365.7|ICD9CM|Glaucoma stage|Glaucoma stage
C3161085|T033|AB|365.70|ICD9CM|Glaucoma stage NOS|Glaucoma stage NOS
C3161085|T033|PT|365.70|ICD9CM|Glaucoma stage, unspecified|Glaucoma stage, unspecified
C3161086|T033|AB|365.71|ICD9CM|Mild stage glaucoma|Mild stage glaucoma
C3161086|T033|PT|365.71|ICD9CM|Mild stage glaucoma|Mild stage glaucoma
C3161087|T033|AB|365.72|ICD9CM|Moderate stage glaucoma|Moderate stage glaucoma
C3161087|T033|PT|365.72|ICD9CM|Moderate stage glaucoma|Moderate stage glaucoma
C3161088|T033|AB|365.73|ICD9CM|Severe stage glaucoma|Severe stage glaucoma
C3161088|T033|PT|365.73|ICD9CM|Severe stage glaucoma|Severe stage glaucoma
C3161089|T047|AB|365.74|ICD9CM|Indeterm stage glaucoma|Indeterm stage glaucoma
C3161089|T047|PT|365.74|ICD9CM|Indeterminate stage glaucoma|Indeterminate stage glaucoma
C0029802|T047|HT|365.8|ICD9CM|Other specified forms of glaucoma|Other specified forms of glaucoma
C0154968|T047|AB|365.81|ICD9CM|Hypersecretion glaucoma|Hypersecretion glaucoma
C0154968|T047|PT|365.81|ICD9CM|Hypersecretion glaucoma|Hypersecretion glaucoma
C0339596|T047|AB|365.82|ICD9CM|Glauc w inc episcl press|Glauc w inc episcl press
C0339596|T047|PT|365.82|ICD9CM|Glaucoma with increased episcleral venous pressure|Glaucoma with increased episcleral venous pressure
C1135189|T047|AB|365.83|ICD9CM|Aqueous misdirection|Aqueous misdirection
C1135189|T047|PT|365.83|ICD9CM|Aqueous misdirection|Aqueous misdirection
C0029802|T047|AB|365.89|ICD9CM|Glaucoma NEC|Glaucoma NEC
C0029802|T047|PT|365.89|ICD9CM|Other specified glaucoma|Other specified glaucoma
C0017601|T047|AB|365.9|ICD9CM|Glaucoma NOS|Glaucoma NOS
C0017601|T047|PT|365.9|ICD9CM|Unspecified glaucoma|Unspecified glaucoma
C0086543|T020|HT|366|ICD9CM|Cataract|Cataract
C0154970|T047|HT|366.0|ICD9CM|Infantile, juvenile, and presenile cataract|Infantile, juvenile, and presenile cataract
C2607928|T020|AB|366.00|ICD9CM|Nonsenile cataract NOS|Nonsenile cataract NOS
C2607928|T020|PT|366.00|ICD9CM|Nonsenile cataract, unspecified|Nonsenile cataract, unspecified
C1112690|T020|AB|366.01|ICD9CM|Ant subcaps pol cataract|Ant subcaps pol cataract
C1112690|T020|PT|366.01|ICD9CM|Anterior subcapsular polar cataract|Anterior subcapsular polar cataract
C1112781|T020|AB|366.02|ICD9CM|Post subcaps pol catarct|Post subcaps pol catarct
C1112781|T020|PT|366.02|ICD9CM|Posterior subcapsular polar cataract|Posterior subcapsular polar cataract
C0154974|T047|AB|366.03|ICD9CM|Cortical cataract|Cortical cataract
C0154974|T047|PT|366.03|ICD9CM|Cortical, lamellar, or zonular cataract|Cortical, lamellar, or zonular cataract
C1112705|T047|AB|366.04|ICD9CM|Nuclear cataract|Nuclear cataract
C1112705|T047|PT|366.04|ICD9CM|Nuclear cataract|Nuclear cataract
C0154976|T020|AB|366.09|ICD9CM|Nonsenile cataract NEC|Nonsenile cataract NEC
C0154976|T020|PT|366.09|ICD9CM|Other and combined forms of nonsenile cataract|Other and combined forms of nonsenile cataract
C0036646|T020|HT|366.1|ICD9CM|Senile cataract|Senile cataract
C0036646|T020|AB|366.10|ICD9CM|Senile cataract NOS|Senile cataract NOS
C0036646|T020|PT|366.10|ICD9CM|Senile cataract, unspecified|Senile cataract, unspecified
C0311341|T047|AB|366.11|ICD9CM|Pseudoexfol lens capsule|Pseudoexfol lens capsule
C0311341|T047|PT|366.11|ICD9CM|Pseudoexfoliation of lens capsule|Pseudoexfoliation of lens capsule
C2939157|T047|AB|366.12|ICD9CM|Incipient cataract|Incipient cataract
C2939157|T047|PT|366.12|ICD9CM|Incipient senile cataract|Incipient senile cataract
C0154978|T047|AB|366.13|ICD9CM|Ant subcaps senile catar|Ant subcaps senile catar
C0154978|T047|PT|366.13|ICD9CM|Anterior subcapsular polar senile cataract|Anterior subcapsular polar senile cataract
C0154979|T047|AB|366.14|ICD9CM|Post subcap senile catar|Post subcap senile catar
C0154979|T047|PT|366.14|ICD9CM|Posterior subcapsular polar senile cataract|Posterior subcapsular polar senile cataract
C0154980|T047|AB|366.15|ICD9CM|Cortical senile cataract|Cortical senile cataract
C0154980|T047|PT|366.15|ICD9CM|Cortical senile cataract|Cortical senile cataract
C0271166|T020|AB|366.16|ICD9CM|Senile nuclear cataract|Senile nuclear cataract
C0271166|T020|PT|366.16|ICD9CM|Senile nuclear sclerosis|Senile nuclear sclerosis
C3665439|T020|AB|366.17|ICD9CM|Mature cataract|Mature cataract
C3665439|T020|PT|366.17|ICD9CM|Total or mature cataract|Total or mature cataract
C0152258|T047|AB|366.18|ICD9CM|Hypermature cataract|Hypermature cataract
C0152258|T047|PT|366.18|ICD9CM|Hypermature cataract|Hypermature cataract
C0154982|T020|PT|366.19|ICD9CM|Other and combined forms of senile cataract|Other and combined forms of senile cataract
C0154982|T020|AB|366.19|ICD9CM|Senile cataract NEC|Senile cataract NEC
C0154983|T037|HT|366.2|ICD9CM|Traumatic cataract|Traumatic cataract
C0154983|T037|AB|366.20|ICD9CM|Traumatic cataract NOS|Traumatic cataract NOS
C0154983|T037|PT|366.20|ICD9CM|Traumatic cataract, unspecified|Traumatic cataract, unspecified
C0154984|T037|AB|366.21|ICD9CM|Local traumatic opacity|Local traumatic opacity
C0154984|T037|PT|366.21|ICD9CM|Localized traumatic opacities|Localized traumatic opacities
C0154985|T037|AB|366.22|ICD9CM|Total traumatic cataract|Total traumatic cataract
C0154985|T037|PT|366.22|ICD9CM|Total traumatic cataract|Total traumatic cataract
C0154986|T037|AB|366.23|ICD9CM|Part resolv traum catar|Part resolv traum catar
C0154986|T037|PT|366.23|ICD9CM|Partially resolved traumatic cataract|Partially resolved traumatic cataract
C0152259|T047|HT|366.3|ICD9CM|Cataract secondary to ocular disorders|Cataract secondary to ocular disorders
C4721766|T047|AB|366.30|ICD9CM|Cataracta complicata NOS|Cataracta complicata NOS
C4721766|T047|PT|366.30|ICD9CM|Cataracta complicata, unspecified|Cataracta complicata, unspecified
C0154989|T047|AB|366.31|ICD9CM|Glaucomatous flecks|Glaucomatous flecks
C0154989|T047|PT|366.31|ICD9CM|Glaucomatous flecks (subcapsular)|Glaucomatous flecks (subcapsular)
C0154990|T047|AB|366.32|ICD9CM|Cataract in inflam dis|Cataract in inflam dis
C0154990|T047|PT|366.32|ICD9CM|Cataract in inflammatory ocular disorders|Cataract in inflammatory ocular disorders
C0271172|T020|AB|366.33|ICD9CM|Cataract w neovasculizat|Cataract w neovasculizat
C0271172|T020|PT|366.33|ICD9CM|Cataract with neovascularization|Cataract with neovascularization
C0154992|T047|AB|366.34|ICD9CM|Cataract in degen dis|Cataract in degen dis
C0154992|T047|PT|366.34|ICD9CM|Cataract in degenerative ocular disorders|Cataract in degenerative ocular disorders
C0154994|T047|HT|366.4|ICD9CM|Cataract associated with other disorders|Cataract associated with other disorders
C0011876|T047|AB|366.41|ICD9CM|Diabetic cataract|Diabetic cataract
C0011876|T047|PT|366.41|ICD9CM|Diabetic cataract|Diabetic cataract
C0039613|T047|AB|366.42|ICD9CM|Tetanic cataract|Tetanic cataract
C0039613|T047|PT|366.42|ICD9CM|Tetanic cataract|Tetanic cataract
C0027128|T047|AB|366.43|ICD9CM|Myotonic cataract|Myotonic cataract
C0027128|T047|PT|366.43|ICD9CM|Myotonic cataract|Myotonic cataract
C0154994|T047|PT|366.44|ICD9CM|Cataract associated with other syndromes|Cataract associated with other syndromes
C0154994|T047|AB|366.44|ICD9CM|Cataract w syndrome NEC|Cataract w syndrome NEC
C0154995|T037|AB|366.45|ICD9CM|Toxic cataract|Toxic cataract
C0154995|T037|PT|366.45|ICD9CM|Toxic cataract|Toxic cataract
C0154996|T020|PT|366.46|ICD9CM|Cataract associated with radiation and other physical influences|Cataract associated with radiation and other physical influences
C0154996|T020|AB|366.46|ICD9CM|Cataract w radiation|Cataract w radiation
C1306068|T047|HT|366.5|ICD9CM|After-cataract|After-cataract
C1306068|T047|AB|366.50|ICD9CM|After-cataract NOS|After-cataract NOS
C1306068|T047|PT|366.50|ICD9CM|After-cataract, unspecified|After-cataract, unspecified
C0152260|T033|AB|366.51|ICD9CM|Soemmering's ring|Soemmering's ring
C0152260|T033|PT|366.51|ICD9CM|Soemmering's ring|Soemmering's ring
C0154997|T020|AB|366.52|ICD9CM|After-cataract NEC|After-cataract NEC
C0154997|T020|PT|366.52|ICD9CM|Other after-cataract, not obscuring vision|Other after-cataract, not obscuring vision
C0154998|T020|PT|366.53|ICD9CM|After-cataract, obscuring vision|After-cataract, obscuring vision
C0154998|T020|AB|366.53|ICD9CM|Aftr-catar obscur vision|Aftr-catar obscur vision
C0029531|T047|AB|366.8|ICD9CM|Cataract NEC|Cataract NEC
C0029531|T047|PT|366.8|ICD9CM|Other cataract|Other cataract
C0086543|T020|AB|366.9|ICD9CM|Cataract NOS|Cataract NOS
C0086543|T020|PT|366.9|ICD9CM|Unspecified cataract|Unspecified cataract
C0339670|T047|HT|367|ICD9CM|Disorders of refraction and accommodation|Disorders of refraction and accommodation
C0020490|T047|AB|367.0|ICD9CM|Hypermetropia|Hypermetropia
C0020490|T047|PT|367.0|ICD9CM|Hypermetropia|Hypermetropia
C0027092|T047|AB|367.1|ICD9CM|Myopia|Myopia
C0027092|T047|PT|367.1|ICD9CM|Myopia|Myopia
C0004106|T047|HT|367.2|ICD9CM|Astigmatism|Astigmatism
C0004106|T047|AB|367.20|ICD9CM|Astigmatism NOS|Astigmatism NOS
C0004106|T047|PT|367.20|ICD9CM|Astigmatism, unspecified|Astigmatism, unspecified
C0152193|T047|AB|367.21|ICD9CM|Regular astigmatism|Regular astigmatism
C0152193|T047|PT|367.21|ICD9CM|Regular astigmatism|Regular astigmatism
C0152194|T047|AB|367.22|ICD9CM|Irregular astigmatism|Irregular astigmatism
C0152194|T047|PT|367.22|ICD9CM|Irregular astigmatism|Irregular astigmatism
C0154999|T047|HT|367.3|ICD9CM|Anisometropia and aniseikonia|Anisometropia and aniseikonia
C0003081|T047|AB|367.31|ICD9CM|Anisometropia|Anisometropia
C0003081|T047|PT|367.31|ICD9CM|Anisometropia|Anisometropia
C0003078|T184|AB|367.32|ICD9CM|Aniseikonia|Aniseikonia
C0003078|T184|PT|367.32|ICD9CM|Aniseikonia|Aniseikonia
C0033075|T047|AB|367.4|ICD9CM|Presbyopia|Presbyopia
C0033075|T047|PT|367.4|ICD9CM|Presbyopia|Presbyopia
C0152198|T047|HT|367.5|ICD9CM|Disorders of accommodation|Disorders of accommodation
C0235238|T047|AB|367.51|ICD9CM|Paresis of accommodation|Paresis of accommodation
C0235238|T047|PT|367.51|ICD9CM|Paresis of accommodation|Paresis of accommodation
C0152197|T047|AB|367.52|ICD9CM|Tot intern ophthalmopleg|Tot intern ophthalmopleg
C0152197|T047|PT|367.52|ICD9CM|Total or complete internal ophthalmoplegia|Total or complete internal ophthalmoplegia
C0152196|T047|AB|367.53|ICD9CM|Spasm of accommodation|Spasm of accommodation
C0152196|T047|PT|367.53|ICD9CM|Spasm of accommodation|Spasm of accommodation
C0029596|T047|HT|367.8|ICD9CM|Other disorders of refraction and accommodation|Other disorders of refraction and accommodation
C0155000|T047|AB|367.81|ICD9CM|Transient refract change|Transient refract change
C0155000|T047|PT|367.81|ICD9CM|Transient refractive change|Transient refractive change
C0029596|T047|PT|367.89|ICD9CM|Other disorders of refraction and accommodation|Other disorders of refraction and accommodation
C0029596|T047|AB|367.89|ICD9CM|Refraction disorder NEC|Refraction disorder NEC
C0339670|T047|AB|367.9|ICD9CM|Refraction disorder NOS|Refraction disorder NOS
C0339670|T047|PT|367.9|ICD9CM|Unspecified disorder of refraction and accommodation|Unspecified disorder of refraction and accommodation
C0547030|T033|HT|368|ICD9CM|Visual disturbances|Visual disturbances
C0152187|T020|HT|368.0|ICD9CM|Amblyopia ex anopsia|Amblyopia ex anopsia
C0002418|T047|AB|368.00|ICD9CM|Amblyopia NOS|Amblyopia NOS
C0002418|T047|PT|368.00|ICD9CM|Amblyopia, unspecified|Amblyopia, unspecified
C0750903|T047|AB|368.01|ICD9CM|Strabismic amblyopia|Strabismic amblyopia
C0750903|T047|PT|368.01|ICD9CM|Strabismic amblyopia|Strabismic amblyopia
C0152189|T047|AB|368.02|ICD9CM|Deprivation amblyopia|Deprivation amblyopia
C0152189|T047|PT|368.02|ICD9CM|Deprivation amblyopia|Deprivation amblyopia
C0152190|T047|AB|368.03|ICD9CM|Refractive amblyopia|Refractive amblyopia
C0152190|T047|PT|368.03|ICD9CM|Refractive amblyopia|Refractive amblyopia
C0155001|T184|HT|368.1|ICD9CM|Subjective visual disturbances|Subjective visual disturbances
C0155001|T184|AB|368.10|ICD9CM|Subj visual disturb NOS|Subj visual disturb NOS
C0155001|T184|PT|368.10|ICD9CM|Subjective visual disturbance, unspecified|Subjective visual disturbance, unspecified
C0155002|T184|AB|368.11|ICD9CM|Sudden visual loss|Sudden visual loss
C0155002|T184|PT|368.11|ICD9CM|Sudden visual loss|Sudden visual loss
C0155003|T046|AB|368.12|ICD9CM|Transient visual loss|Transient visual loss
C0155003|T046|PT|368.12|ICD9CM|Transient visual loss|Transient visual loss
C0042818|T184|AB|368.13|ICD9CM|Visual discomfort|Visual discomfort
C0042818|T184|PT|368.13|ICD9CM|Visual discomfort|Visual discomfort
C0155004|T184|AB|368.14|ICD9CM|Distortion of shape/size|Distortion of shape/size
C0155004|T184|PT|368.14|ICD9CM|Visual distortions of shape and size|Visual distortions of shape and size
C0155005|T047|PT|368.15|ICD9CM|Other visual distortions and entoptic phenomena|Other visual distortions and entoptic phenomena
C0155005|T047|AB|368.15|ICD9CM|Visual distortions NEC|Visual distortions NEC
C0155006|T047|AB|368.16|ICD9CM|Psychophysic visual dist|Psychophysic visual dist
C0155006|T047|PT|368.16|ICD9CM|Psychophysical visual disturbances|Psychophysical visual disturbances
C0012569|T033|AB|368.2|ICD9CM|Diplopia|Diplopia
C0012569|T033|PT|368.2|ICD9CM|Diplopia|Diplopia
C0155007|T047|HT|368.3|ICD9CM|Other disorders of binocular vision|Other disorders of binocular vision
C0005461|T047|AB|368.30|ICD9CM|Binocular vision dis NOS|Binocular vision dis NOS
C0005461|T047|PT|368.30|ICD9CM|Binocular vision disorder, unspecified|Binocular vision disorder, unspecified
C0221103|T046|AB|368.31|ICD9CM|Binocular vis suppress|Binocular vis suppress
C0221103|T046|PT|368.31|ICD9CM|Suppression of binocular vision|Suppression of binocular vision
C0155008|T047|PT|368.32|ICD9CM|Simultaneous visual perception without fusion|Simultaneous visual perception without fusion
C0155008|T047|AB|368.32|ICD9CM|Visual percept w/o fusn|Visual percept w/o fusn
C0155009|T047|AB|368.33|ICD9CM|Fusion w def stereopsis|Fusion w def stereopsis
C0155009|T047|PT|368.33|ICD9CM|Fusion with defective stereopsis|Fusion with defective stereopsis
C0155010|T047|AB|368.34|ICD9CM|Abn retina correspond|Abn retina correspond
C0155010|T047|PT|368.34|ICD9CM|Abnormal retinal correspondence|Abnormal retinal correspondence
C3887875|T033|HT|368.4|ICD9CM|Visual field defects|Visual field defects
C3887875|T033|AB|368.40|ICD9CM|Visual field defect NOS|Visual field defect NOS
C3887875|T033|PT|368.40|ICD9CM|Visual field defect, unspecified|Visual field defect, unspecified
C0152191|T033|AB|368.41|ICD9CM|Central scotoma|Central scotoma
C0152191|T033|PT|368.41|ICD9CM|Scotoma involving central area|Scotoma involving central area
C0152192|T033|AB|368.42|ICD9CM|Scotoma of blind spot|Scotoma of blind spot
C0152192|T033|PT|368.42|ICD9CM|Scotoma of blind spot area|Scotoma of blind spot area
C3839935|T033|AB|368.43|ICD9CM|Sector or arcuate defect|Sector or arcuate defect
C3839935|T033|PT|368.43|ICD9CM|Sector or arcuate visual field defects|Sector or arcuate visual field defects
C0029657|T047|PT|368.44|ICD9CM|Other localized visual field defect|Other localized visual field defect
C0029657|T047|AB|368.44|ICD9CM|Visual field defect NEC|Visual field defect NEC
C0155012|T047|AB|368.45|ICD9CM|Gen visual contraction|Gen visual contraction
C0155012|T047|PT|368.45|ICD9CM|Generalized visual field contraction or constriction|Generalized visual field contraction or constriction
C0271202|T047|PT|368.46|ICD9CM|Homonymous bilateral field defects|Homonymous bilateral field defects
C0271202|T047|AB|368.46|ICD9CM|Homonymous hemianopsia|Homonymous hemianopsia
C0271207|T033|PT|368.47|ICD9CM|Heteronymous bilateral field defects|Heteronymous bilateral field defects
C0271207|T033|AB|368.47|ICD9CM|Heteronymous hemianopsia|Heteronymous hemianopsia
C0242225|T047|HT|368.5|ICD9CM|Color vision deficiencies|Color vision deficiencies
C0155015|T047|AB|368.51|ICD9CM|Protan defect|Protan defect
C0155015|T047|PT|368.51|ICD9CM|Protan defect|Protan defect
C0155016|T047|AB|368.52|ICD9CM|Deutan defect|Deutan defect
C0155016|T047|PT|368.52|ICD9CM|Deutan defect|Deutan defect
C0155017|T047|AB|368.53|ICD9CM|Tritan defect|Tritan defect
C0155017|T047|PT|368.53|ICD9CM|Tritan defect|Tritan defect
C0152200|T047|AB|368.54|ICD9CM|Achromatopsia|Achromatopsia
C0152200|T047|PT|368.54|ICD9CM|Achromatopsia|Achromatopsia
C0155018|T047|AB|368.55|ICD9CM|Acq color deficiency|Acq color deficiency
C0155018|T047|PT|368.55|ICD9CM|Acquired color vision deficiencies|Acquired color vision deficiencies
C0029548|T047|AB|368.59|ICD9CM|Color deficiency NEC|Color deficiency NEC
C0029548|T047|PT|368.59|ICD9CM|Other color vision deficiencies|Other color vision deficiencies
C0028077|T047|HT|368.6|ICD9CM|Night blindness|Night blindness
C0028077|T047|AB|368.60|ICD9CM|Night blindness NOS|Night blindness NOS
C0028077|T047|PT|368.60|ICD9CM|Night blindness, unspecified|Night blindness, unspecified
C1306122|T047|AB|368.61|ICD9CM|Congen night blindness|Congen night blindness
C1306122|T047|PT|368.61|ICD9CM|Congenital night blindness|Congenital night blindness
C0152202|T020|AB|368.62|ICD9CM|Acquired night blindness|Acquired night blindness
C0152202|T020|PT|368.62|ICD9CM|Acquired night blindness|Acquired night blindness
C0155019|T047|AB|368.63|ICD9CM|Abn dark adaptat curve|Abn dark adaptat curve
C0155019|T047|PT|368.63|ICD9CM|Abnormal dark adaptation curve|Abnormal dark adaptation curve
C0029672|T047|AB|368.69|ICD9CM|Night blindness NEC|Night blindness NEC
C0029672|T047|PT|368.69|ICD9CM|Other night blindness|Other night blindness
C0029844|T184|PT|368.8|ICD9CM|Other specified visual disturbances|Other specified visual disturbances
C0029844|T184|AB|368.8|ICD9CM|Visual disturbances NEC|Visual disturbances NEC
C0547030|T033|PT|368.9|ICD9CM|Unspecified visual disturbance|Unspecified visual disturbance
C0547030|T033|AB|368.9|ICD9CM|Visual disturbance NOS|Visual disturbance NOS
C0155020|T047|HT|369|ICD9CM|Blindness and low vision|Blindness and low vision
C0155021|T047|HT|369.0|ICD9CM|Profound vision impairment, both eyes|Profound vision impairment, both eyes
C1879328|T047|AB|369.00|ICD9CM|Both eyes blind-who def|Both eyes blind-who def
C1879328|T047|PT|369.00|ICD9CM|Profound impairment, both eyes, impairment level not further specified|Profound impairment, both eyes, impairment level not further specified
C0155022|T047|PT|369.01|ICD9CM|Better eye: total vision impairment; lesser eye: total vision impairment|Better eye: total vision impairment; lesser eye: total vision impairment
C0155022|T047|AB|369.01|ICD9CM|Tot impairment-both eyes|Tot impairment-both eyes
C0521709|T047|PT|369.02|ICD9CM|Better eye: near-total vision impairment; lesser eye: not further specified|Better eye: near-total vision impairment; lesser eye: not further specified
C0521709|T047|AB|369.02|ICD9CM|One eye-near tot/oth-NOS|One eye-near tot/oth-NOS
C0392558|T047|PT|369.03|ICD9CM|Better eye: near-total vision impairment; lesser eye: total vision impairment|Better eye: near-total vision impairment; lesser eye: total vision impairment
C0392558|T047|AB|369.03|ICD9CM|One eye-near tot/oth-tot|One eye-near tot/oth-tot
C0271220|T033|PT|369.04|ICD9CM|Better eye: near-total vision impairment; lesser eye: near-total vision impairment|Better eye: near-total vision impairment; lesser eye: near-total vision impairment
C0271220|T033|AB|369.04|ICD9CM|Near-tot impair-both eye|Near-tot impair-both eye
C0392559|T047|PT|369.05|ICD9CM|Better eye: profound vision impairment; lesser eye: not further specified|Better eye: profound vision impairment; lesser eye: not further specified
C0392559|T047|AB|369.05|ICD9CM|One eye-profound/oth-NOS|One eye-profound/oth-NOS
C0392560|T033|PT|369.06|ICD9CM|Better eye: profound vision impairment; lesser eye: total vision impairment|Better eye: profound vision impairment; lesser eye: total vision impairment
C0392560|T033|AB|369.06|ICD9CM|One eye-profound/oth-tot|One eye-profound/oth-tot
C0392561|T047|PT|369.07|ICD9CM|Better eye: profound vision impairment; lesser eye: near-total vision impairment|Better eye: profound vision impairment; lesser eye: near-total vision impairment
C0392561|T047|AB|369.07|ICD9CM|One eye-prfnd/oth-nr tot|One eye-prfnd/oth-nr tot
C0271224|T047|PT|369.08|ICD9CM|Better eye: profound vision impairment; lesser eye: profound vision impairment|Better eye: profound vision impairment; lesser eye: profound vision impairment
C0271224|T047|AB|369.08|ICD9CM|Profound impair both eye|Profound impair both eye
C0339701|T047|HT|369.1|ICD9CM|Moderate or severe vision impairment, better eye; profound vision impairment of lesser eye|Moderate or severe vision impairment, better eye; profound vision impairment of lesser eye
C0271225|T047|AB|369.10|ICD9CM|Blindness/low vision|Blindness/low vision
C0271225|T047|PT|369.10|ICD9CM|Moderate or severe impairment, better eye, impairment level not further specified|Moderate or severe impairment, better eye, impairment level not further specified
C0392562|T047|AB|369.11|ICD9CM|1 eye-sev/oth-blind NOS|1 eye-sev/oth-blind NOS
C0392562|T047|PT|369.11|ICD9CM|Better eye: severe vision impairment; lesser eye: blind, not further specified|Better eye: severe vision impairment; lesser eye: blind, not further specified
C0392563|T033|PT|369.12|ICD9CM|Better eye: severe vision impairment; lesser eye: total vision impairment|Better eye: severe vision impairment; lesser eye: total vision impairment
C0392563|T033|AB|369.12|ICD9CM|One eye-severe/oth-total|One eye-severe/oth-total
C0392564|T033|PT|369.13|ICD9CM|Better eye: severe vision impairment; lesser eye: near-total vision impairment|Better eye: severe vision impairment; lesser eye: near-total vision impairment
C0392564|T033|AB|369.13|ICD9CM|One eye-sev/oth-near tot|One eye-sev/oth-near tot
C0392565|T033|PT|369.14|ICD9CM|Better eye: severe vision impairment; lesser eye: profound vision impairment|Better eye: severe vision impairment; lesser eye: profound vision impairment
C0392565|T033|AB|369.14|ICD9CM|One eye-sev/oth-prfnd|One eye-sev/oth-prfnd
C0392566|T033|PT|369.15|ICD9CM|Better eye: moderate vision impairment; lesser eye: blind, not further specified|Better eye: moderate vision impairment; lesser eye: blind, not further specified
C0392566|T033|AB|369.15|ICD9CM|One eye-mod/oth-blind|One eye-mod/oth-blind
C0392567|T033|PT|369.16|ICD9CM|Better eye: moderate vision impairment; lesser eye: total vision impairment|Better eye: moderate vision impairment; lesser eye: total vision impairment
C0392567|T033|AB|369.16|ICD9CM|One eye-moderate/oth-tot|One eye-moderate/oth-tot
C0392568|T033|PT|369.17|ICD9CM|Better eye: moderate vision impairment; lesser eye: near-total vision impairment|Better eye: moderate vision impairment; lesser eye: near-total vision impairment
C0392568|T033|AB|369.17|ICD9CM|One eye-mod/oth-near tot|One eye-mod/oth-near tot
C0392569|T033|PT|369.18|ICD9CM|Better eye: moderate vision impairment; lesser eye: profound vision impairment|Better eye: moderate vision impairment; lesser eye: profound vision impairment
C0392569|T033|AB|369.18|ICD9CM|One eye-mod/oth-profound|One eye-mod/oth-profound
C0155040|T047|HT|369.2|ICD9CM|Moderate or severe vision impairment, both eyes|Moderate or severe vision impairment, both eyes
C0271234|T047|AB|369.20|ICD9CM|Low vision, 2 eyes NOS|Low vision, 2 eyes NOS
C0271234|T047|PT|369.20|ICD9CM|Moderate or severe impairment, both eyes, impairment level not further specified|Moderate or severe impairment, both eyes, impairment level not further specified
C0392570|T033|PT|369.21|ICD9CM|Better eye: severe vision impairment; lesser eye; impairment not further specified|Better eye: severe vision impairment; lesser eye; impairment not further specified
C0392570|T033|AB|369.21|ICD9CM|One eye-severe/oth-NOS|One eye-severe/oth-NOS
C0271236|T033|PT|369.22|ICD9CM|Better eye: severe vision impairment; lesser eye: severe vision impairment|Better eye: severe vision impairment; lesser eye: severe vision impairment
C0271236|T033|AB|369.22|ICD9CM|Severe impair-both eyes|Severe impair-both eyes
C0392571|T047|PT|369.23|ICD9CM|Better eye: moderate vision impairment; lesser eye: impairment not further specified|Better eye: moderate vision impairment; lesser eye: impairment not further specified
C0392571|T047|AB|369.23|ICD9CM|One eye-moderate/oth-NOS|One eye-moderate/oth-NOS
C0392572|T033|PT|369.24|ICD9CM|Better eye: moderate vision impairment; lesser eye: severe vision impairment|Better eye: moderate vision impairment; lesser eye: severe vision impairment
C0392572|T033|AB|369.24|ICD9CM|One eye-moderate/oth-sev|One eye-moderate/oth-sev
C0271239|T033|PT|369.25|ICD9CM|Better eye: moderate vision impairment; lesser eye: moderate vision impairment|Better eye: moderate vision impairment; lesser eye: moderate vision impairment
C0271239|T033|AB|369.25|ICD9CM|Moderate impair-both eye|Moderate impair-both eye
C0155047|T184|AB|369.3|ICD9CM|Blindness NOS, both eyes|Blindness NOS, both eyes
C0155047|T184|PT|369.3|ICD9CM|Unqualified visual loss, both eyes|Unqualified visual loss, both eyes
C0339711|T033|AB|369.4|ICD9CM|Legal blindness-usa def|Legal blindness-usa def
C0339711|T033|PT|369.4|ICD9CM|Legal blindness, as defined in U.S.A.|Legal blindness, as defined in U.S.A.
C0155049|T047|HT|369.6|ICD9CM|Profound vision impairment, one eye|Profound vision impairment, one eye
C0392578|T033|AB|369.60|ICD9CM|Blindness, one eye|Blindness, one eye
C0392578|T033|PT|369.60|ICD9CM|Profound impairment, one eye, impairment level not further specified|Profound impairment, one eye, impairment level not further specified
C0521710|T033|AB|369.61|ICD9CM|One eye-total/oth-unknwn|One eye-total/oth-unknwn
C0521710|T033|PT|369.61|ICD9CM|One eye: total vision impairment; other eye: not specified|One eye: total vision impairment; other eye: not specified
C0392573|T033|AB|369.62|ICD9CM|One eye-tot/oth-near nor|One eye-tot/oth-near nor
C0392573|T033|PT|369.62|ICD9CM|One eye: total vision impairment; other eye: near-normal vision|One eye: total vision impairment; other eye: near-normal vision
C0392574|T033|AB|369.63|ICD9CM|One eye-total/oth-normal|One eye-total/oth-normal
C0392574|T033|PT|369.63|ICD9CM|One eye: total vision impairment; other eye: normal vision|One eye: total vision impairment; other eye: normal vision
C0392575|T033|AB|369.64|ICD9CM|One eye-near tot/oth-NOS|One eye-near tot/oth-NOS
C0392575|T033|PT|369.64|ICD9CM|One eye: near-total vision impairment; other eye: vision not specified|One eye: near-total vision impairment; other eye: vision not specified
C0392576|T033|AB|369.65|ICD9CM|Near-tot imp/near-normal|Near-tot imp/near-normal
C0392576|T033|PT|369.65|ICD9CM|One eye: near-total vision impairment; other eye: near-normal vision|One eye: near-total vision impairment; other eye: near-normal vision
C0392577|T033|AB|369.66|ICD9CM|Near-total impair/normal|Near-total impair/normal
C0392577|T033|PT|369.66|ICD9CM|One eye: near-total vision impairment; other eye: normal vision|One eye: near-total vision impairment; other eye: normal vision
C0392578|T033|AB|369.67|ICD9CM|One eye-prfound/oth-unkn|One eye-prfound/oth-unkn
C0392578|T033|PT|369.67|ICD9CM|One eye: profound vision impairment; other eye: vision not specified|One eye: profound vision impairment; other eye: vision not specified
C0392579|T033|PT|369.68|ICD9CM|One eye: profound vision impairment; other eye: near-normal vision|One eye: profound vision impairment; other eye: near-normal vision
C0392579|T033|AB|369.68|ICD9CM|Profnd impair/near norm|Profnd impair/near norm
C0392580|T033|PT|369.69|ICD9CM|One eye: profound vision impairment; other eye: normal vision|One eye: profound vision impairment; other eye: normal vision
C0392580|T033|AB|369.69|ICD9CM|Profound impair/normal|Profound impair/normal
C0155058|T047|HT|369.7|ICD9CM|Moderate or severe vision impairment, one eye|Moderate or severe vision impairment, one eye
C0520728|T047|AB|369.70|ICD9CM|Low vision, one eye|Low vision, one eye
C0520728|T047|PT|369.70|ICD9CM|Moderate or severe impairment, one eye, impairment level not further specified|Moderate or severe impairment, one eye, impairment level not further specified
C0392581|T033|AB|369.71|ICD9CM|One eye-severe/oth-unknw|One eye-severe/oth-unknw
C0392581|T033|PT|369.71|ICD9CM|One eye: severe vision impairment; other eye: vision not specified|One eye: severe vision impairment; other eye: vision not specified
C0392582|T033|AB|369.72|ICD9CM|One eye-sev/oth-nr norm|One eye-sev/oth-nr norm
C0392582|T033|PT|369.72|ICD9CM|One eye: severe vision impairment; other eye: near-normal vision|One eye: severe vision impairment; other eye: near-normal vision
C0392583|T033|AB|369.73|ICD9CM|One eye-severe/oth-norm|One eye-severe/oth-norm
C0392583|T033|PT|369.73|ICD9CM|One eye: severe vision impairment; other eye: normal vision|One eye: severe vision impairment; other eye: normal vision
C0392584|T033|AB|369.74|ICD9CM|One eye-mod/other-unknwn|One eye-mod/other-unknwn
C0392584|T033|PT|369.74|ICD9CM|One eye: moderate vision impairment; other eye: vision not specified|One eye: moderate vision impairment; other eye: vision not specified
C0392585|T033|AB|369.75|ICD9CM|One eye-mod/oth-nr norm|One eye-mod/oth-nr norm
C0392585|T033|PT|369.75|ICD9CM|One eye: moderate vision impairment; other eye: near-normal vision|One eye: moderate vision impairment; other eye: near-normal vision
C0392586|T033|AB|369.76|ICD9CM|One eye-mod/oth normal|One eye-mod/oth normal
C0392586|T033|PT|369.76|ICD9CM|One eye: moderate vision impairment; other eye: normal vision|One eye: moderate vision impairment; other eye: normal vision
C0155066|T184|PT|369.8|ICD9CM|Unqualified visual loss, one eye|Unqualified visual loss, one eye
C0155066|T184|AB|369.8|ICD9CM|Visual loss, one eye NOS|Visual loss, one eye NOS
C3665346|T184|PT|369.9|ICD9CM|Unspecified visual loss|Unspecified visual loss
C3665346|T184|AB|369.9|ICD9CM|Visual loss NOS|Visual loss NOS
C0022568|T047|HT|370|ICD9CM|Keratitis|Keratitis
C0010043|T047|HT|370.0|ICD9CM|Corneal ulcer|Corneal ulcer
C0010043|T047|AB|370.00|ICD9CM|Corneal ulcer NOS|Corneal ulcer NOS
C0010043|T047|PT|370.00|ICD9CM|Corneal ulcer, unspecified|Corneal ulcer, unspecified
C0155067|T047|AB|370.01|ICD9CM|Marginal corneal ulcer|Marginal corneal ulcer
C0155067|T047|PT|370.01|ICD9CM|Marginal corneal ulcer|Marginal corneal ulcer
C0155068|T047|AB|370.02|ICD9CM|Ring corneal ulcer|Ring corneal ulcer
C0155068|T047|PT|370.02|ICD9CM|Ring corneal ulcer|Ring corneal ulcer
C0155069|T047|AB|370.03|ICD9CM|Central corneal ulcer|Central corneal ulcer
C0155069|T047|PT|370.03|ICD9CM|Central corneal ulcer|Central corneal ulcer
C0155070|T047|AB|370.04|ICD9CM|Hypopyon ulcer|Hypopyon ulcer
C0155070|T047|PT|370.04|ICD9CM|Hypopyon ulcer|Hypopyon ulcer
C0155071|T047|AB|370.05|ICD9CM|Mycotic corneal ulcer|Mycotic corneal ulcer
C0155071|T047|PT|370.05|ICD9CM|Mycotic corneal ulcer|Mycotic corneal ulcer
C0151844|T047|AB|370.06|ICD9CM|Perforated corneal ulcer|Perforated corneal ulcer
C0151844|T047|PT|370.06|ICD9CM|Perforated corneal ulcer|Perforated corneal ulcer
C0155072|T047|AB|370.07|ICD9CM|Mooren's ulcer|Mooren's ulcer
C0155072|T047|PT|370.07|ICD9CM|Mooren's ulcer|Mooren's ulcer
C0155073|T047|HT|370.2|ICD9CM|Superficial keratitis without conjunctivitis|Superficial keratitis without conjunctivitis
C0155074|T047|AB|370.20|ICD9CM|Superfic keratitis NOS|Superfic keratitis NOS
C0155074|T047|PT|370.20|ICD9CM|Superficial keratitis, unspecified|Superficial keratitis, unspecified
C0259799|T047|AB|370.21|ICD9CM|Punctate keratitis|Punctate keratitis
C0259799|T047|PT|370.21|ICD9CM|Punctate keratitis|Punctate keratitis
C0155076|T047|AB|370.22|ICD9CM|Macular keratitis|Macular keratitis
C0155076|T047|PT|370.22|ICD9CM|Macular keratitis|Macular keratitis
C0155077|T047|AB|370.23|ICD9CM|Filamentary keratitis|Filamentary keratitis
C0155077|T047|PT|370.23|ICD9CM|Filamentary keratitis|Filamentary keratitis
C0155078|T047|AB|370.24|ICD9CM|Photokeratitis|Photokeratitis
C0155078|T047|PT|370.24|ICD9CM|Photokeratitis|Photokeratitis
C0155079|T047|HT|370.3|ICD9CM|Certain types of keratoconjunctivitis|Certain types of keratoconjunctivitis
C0155080|T047|AB|370.31|ICD9CM|Phlycten keratoconjunct|Phlycten keratoconjunct
C0155080|T047|PT|370.31|ICD9CM|Phlyctenular keratoconjunctivitis|Phlyctenular keratoconjunctivitis
C0155081|T047|PT|370.32|ICD9CM|Limbar and corneal involvement in vernal conjunctivitis|Limbar and corneal involvement in vernal conjunctivitis
C0155081|T047|AB|370.32|ICD9CM|Limbar keratoconjunctiv|Limbar keratoconjunctiv
C0155082|T047|AB|370.33|ICD9CM|Keratoconjunctivit sicca|Keratoconjunctivit sicca
C0155082|T047|PT|370.33|ICD9CM|Keratoconjunctivitis sicca, not specified as Sjogren's|Keratoconjunctivitis sicca, not specified as Sjogren's
C0339295|T047|PT|370.34|ICD9CM|Exposure keratoconjunctivitis|Exposure keratoconjunctivitis
C0339295|T047|AB|370.34|ICD9CM|Expsure keratoconjunctiv|Expsure keratoconjunctiv
C0155084|T047|AB|370.35|ICD9CM|Neurotroph keratoconjunc|Neurotroph keratoconjunc
C0155084|T047|PT|370.35|ICD9CM|Neurotrophic keratoconjunctivitis|Neurotrophic keratoconjunctivitis
C0155085|T047|HT|370.4|ICD9CM|Other and unspecified keratoconjunctivitis|Other and unspecified keratoconjunctivitis
C0022573|T047|AB|370.40|ICD9CM|Keratoconjunctivitis NOS|Keratoconjunctivitis NOS
C0022573|T047|PT|370.40|ICD9CM|Keratoconjunctivitis, unspecified|Keratoconjunctivitis, unspecified
C0155086|T047|AB|370.44|ICD9CM|Keratitis in exanthema|Keratitis in exanthema
C0155086|T047|PT|370.44|ICD9CM|Keratitis or keratoconjunctivitis in exanthema|Keratitis or keratoconjunctivitis in exanthema
C0029650|T047|AB|370.49|ICD9CM|Keratoconjunctivitis NEC|Keratoconjunctivitis NEC
C0029650|T047|PT|370.49|ICD9CM|Other keratoconjunctivitis|Other keratoconjunctivitis
C0155087|T047|HT|370.5|ICD9CM|Interstitial and deep keratitis|Interstitial and deep keratitis
C0155088|T047|AB|370.50|ICD9CM|Interstit keratitis NOS|Interstit keratitis NOS
C0155088|T047|PT|370.50|ICD9CM|Interstitial keratitis, unspecified|Interstitial keratitis, unspecified
C0155089|T047|AB|370.52|ICD9CM|Diffus interstit keratit|Diffus interstit keratit
C0155089|T047|PT|370.52|ICD9CM|Diffuse interstitial keratitis|Diffuse interstitial keratitis
C0155090|T047|AB|370.54|ICD9CM|Sclerosing keratitis|Sclerosing keratitis
C0155090|T047|PT|370.54|ICD9CM|Sclerosing keratitis|Sclerosing keratitis
C0155091|T047|AB|370.55|ICD9CM|Corneal abscess|Corneal abscess
C0155091|T047|PT|370.55|ICD9CM|Corneal abscess|Corneal abscess
C0155092|T047|AB|370.59|ICD9CM|Interstit keratitis NEC|Interstit keratitis NEC
C0155092|T047|PT|370.59|ICD9CM|Other interstitial and deep keratitis|Other interstitial and deep keratitis
C0085109|T047|HT|370.6|ICD9CM|Corneal neovascularization|Corneal neovascularization
C0085109|T047|AB|370.60|ICD9CM|Cornea neovasculariz NOS|Cornea neovasculariz NOS
C0085109|T047|PT|370.60|ICD9CM|Corneal neovascularization, unspecified|Corneal neovascularization, unspecified
C0155093|T047|AB|370.61|ICD9CM|Local vasculariza cornea|Local vasculariza cornea
C0155093|T047|PT|370.61|ICD9CM|Localized vascularization of cornea|Localized vascularization of cornea
C0155094|T047|AB|370.62|ICD9CM|Corneal pannus|Corneal pannus
C0155094|T047|PT|370.62|ICD9CM|Pannus (corneal)|Pannus (corneal)
C0155095|T047|AB|370.63|ICD9CM|Deep vasculariza cornea|Deep vasculariza cornea
C0155095|T047|PT|370.63|ICD9CM|Deep vascularization of cornea|Deep vascularization of cornea
C0155096|T190|AB|370.64|ICD9CM|Corneal ghost vessels|Corneal ghost vessels
C0155096|T190|PT|370.64|ICD9CM|Ghost vessels (corneal)|Ghost vessels (corneal)
C0348526|T047|AB|370.8|ICD9CM|Keratitis NEC|Keratitis NEC
C0348526|T047|PT|370.8|ICD9CM|Other forms of keratitis|Other forms of keratitis
C0022568|T047|AB|370.9|ICD9CM|Keratitis NOS|Keratitis NOS
C0022568|T047|PT|370.9|ICD9CM|Unspecified keratitis|Unspecified keratitis
C0155097|T047|HT|371|ICD9CM|Corneal opacity and other disorders of cornea|Corneal opacity and other disorders of cornea
C0155098|T020|HT|371.0|ICD9CM|Corneal scars and opacities|Corneal scars and opacities
C0010038|T033|AB|371.00|ICD9CM|Corneal opacity NOS|Corneal opacity NOS
C0010038|T033|PT|371.00|ICD9CM|Corneal opacity, unspecified|Corneal opacity, unspecified
C0155099|T033|AB|371.01|ICD9CM|Minor opacity of cornea|Minor opacity of cornea
C0155099|T033|PT|371.01|ICD9CM|Minor opacity of cornea|Minor opacity of cornea
C0155100|T033|AB|371.02|ICD9CM|Periph opacity of cornea|Periph opacity of cornea
C0155100|T033|PT|371.02|ICD9CM|Peripheral opacity of cornea|Peripheral opacity of cornea
C0007686|T033|PT|371.03|ICD9CM|Central opacity of cornea|Central opacity of cornea
C0007686|T033|AB|371.03|ICD9CM|Central opacity, cornea|Central opacity, cornea
C0271275|T033|AB|371.04|ICD9CM|Adherent leucoma|Adherent leucoma
C0271275|T033|PT|371.04|ICD9CM|Adherent leucoma|Adherent leucoma
C0155102|T047|AB|371.05|ICD9CM|Phthisical cornea|Phthisical cornea
C0155102|T047|PT|371.05|ICD9CM|Phthisical cornea|Phthisical cornea
C0339249|T033|HT|371.1|ICD9CM|Corneal pigmentations and deposits|Corneal pigmentations and deposits
C0162281|T047|AB|371.10|ICD9CM|Corneal deposit NOS|Corneal deposit NOS
C0162281|T047|PT|371.10|ICD9CM|Corneal deposit, unspecified|Corneal deposit, unspecified
C0155104|T047|AB|371.11|ICD9CM|Ant cornea pigmentation|Ant cornea pigmentation
C0155104|T047|PT|371.11|ICD9CM|Anterior corneal pigmentations|Anterior corneal pigmentations
C0155105|T047|AB|371.12|ICD9CM|Stromal cornea pigment|Stromal cornea pigment
C0155105|T047|PT|371.12|ICD9CM|Stromal corneal pigmentations|Stromal corneal pigmentations
C0155106|T047|AB|371.13|ICD9CM|Post cornea pigmentation|Post cornea pigmentation
C0155106|T047|PT|371.13|ICD9CM|Posterior corneal pigmentations|Posterior corneal pigmentations
C0152457|T047|PT|371.14|ICD9CM|Kayser-Fleischer ring|Kayser-Fleischer ring
C0152457|T047|AB|371.14|ICD9CM|Kayser-fleischer ring|Kayser-fleischer ring
C0155107|T047|AB|371.15|ICD9CM|Oth deposit w metab dis|Oth deposit w metab dis
C0155107|T047|PT|371.15|ICD9CM|Other corneal deposits associated with metabolic disorders|Other corneal deposits associated with metabolic disorders
C0155108|T047|AB|371.16|ICD9CM|Argentous cornea deposit|Argentous cornea deposit
C0155108|T047|PT|371.16|ICD9CM|Argentous corneal deposits|Argentous corneal deposits
C0010037|T046|HT|371.2|ICD9CM|Corneal edema|Corneal edema
C0010037|T046|AB|371.20|ICD9CM|Corneal edema NOS|Corneal edema NOS
C0010037|T046|PT|371.20|ICD9CM|Corneal edema, unspecified|Corneal edema, unspecified
C0155109|T047|AB|371.21|ICD9CM|Idiopathic corneal edema|Idiopathic corneal edema
C0155109|T047|PT|371.21|ICD9CM|Idiopathic corneal edema|Idiopathic corneal edema
C0155110|T047|AB|371.22|ICD9CM|Secondary corneal edema|Secondary corneal edema
C0155110|T047|PT|371.22|ICD9CM|Secondary corneal edema|Secondary corneal edema
C0155111|T047|AB|371.23|ICD9CM|Bullous keratopathy|Bullous keratopathy
C0155111|T047|PT|371.23|ICD9CM|Bullous keratopathy|Bullous keratopathy
C0474442|T047|PT|371.24|ICD9CM|Corneal edema due to wearing of contact lenses|Corneal edema due to wearing of contact lenses
C0474442|T047|AB|371.24|ICD9CM|Edema d/t contact lens|Edema d/t contact lens
C0155114|T020|HT|371.3|ICD9CM|Changes of corneal membranes|Changes of corneal membranes
C0155114|T020|AB|371.30|ICD9CM|Cornea memb change NOS|Cornea memb change NOS
C0155114|T020|PT|371.30|ICD9CM|Corneal membrane change, unspecified|Corneal membrane change, unspecified
C0155115|T047|AB|371.31|ICD9CM|Fold of bowman membrane|Fold of bowman membrane
C0155115|T047|PT|371.31|ICD9CM|Folds and rupture of bowman's membrane|Folds and rupture of bowman's membrane
C0155116|T190|AB|371.32|ICD9CM|Fold in descemet membran|Fold in descemet membran
C0155116|T190|PT|371.32|ICD9CM|Folds in descemet's membrane|Folds in descemet's membrane
C0155117|T020|AB|371.33|ICD9CM|Rupture descemet membran|Rupture descemet membran
C0155117|T020|PT|371.33|ICD9CM|Rupture in descemet's membrane|Rupture in descemet's membrane
C0155118|T047|HT|371.4|ICD9CM|Corneal degenerations|Corneal degenerations
C0155118|T047|AB|371.40|ICD9CM|Corneal degeneration NOS|Corneal degeneration NOS
C0155118|T047|PT|371.40|ICD9CM|Corneal degeneration, unspecified|Corneal degeneration, unspecified
C0036647|T020|AB|371.41|ICD9CM|Senile corneal changes|Senile corneal changes
C0036647|T020|PT|371.41|ICD9CM|Senile corneal changes|Senile corneal changes
C0155119|T047|AB|371.42|ICD9CM|Recurrent cornea erosion|Recurrent cornea erosion
C0155119|T047|PT|371.42|ICD9CM|Recurrent erosion of cornea|Recurrent erosion of cornea
C0155120|T047|AB|371.43|ICD9CM|Band-shaped keratopathy|Band-shaped keratopathy
C0155120|T047|PT|371.43|ICD9CM|Band-shaped keratopathy|Band-shaped keratopathy
C0155121|T047|AB|371.44|ICD9CM|Calcer cornea degen NEC|Calcer cornea degen NEC
C0155121|T047|PT|371.44|ICD9CM|Other calcerous degenerations of cornea|Other calcerous degenerations of cornea
C0152455|T047|AB|371.45|ICD9CM|Keratomalacia NOS|Keratomalacia NOS
C0152455|T047|PT|371.45|ICD9CM|Keratomalacia NOS|Keratomalacia NOS
C0155122|T047|AB|371.46|ICD9CM|Nodular cornea degen|Nodular cornea degen
C0155122|T047|PT|371.46|ICD9CM|Nodular degeneration of cornea|Nodular degeneration of cornea
C0155123|T047|AB|371.48|ICD9CM|Peripheral cornea degen|Peripheral cornea degen
C0155123|T047|PT|371.48|ICD9CM|Peripheral degenerations of cornea|Peripheral degenerations of cornea
C0155124|T047|AB|371.49|ICD9CM|Cornea degeneration NEC|Cornea degeneration NEC
C0155124|T047|PT|371.49|ICD9CM|Other corneal degenerations|Other corneal degenerations
C0010035|T047|HT|371.5|ICD9CM|Hereditary corneal dystrophies|Hereditary corneal dystrophies
C0010035|T047|AB|371.50|ICD9CM|Corneal dystrophy NOS|Corneal dystrophy NOS
C0010035|T047|PT|371.50|ICD9CM|Hereditary corneal dystrophy, unspecified|Hereditary corneal dystrophy, unspecified
C0339277|T019|AB|371.51|ICD9CM|Juv epith cornea dystrph|Juv epith cornea dystrph
C0339277|T019|PT|371.51|ICD9CM|Juvenile epithelial corneal dystrophy|Juvenile epithelial corneal dystrophy
C0155126|T047|AB|371.52|ICD9CM|Ant cornea dystrophy NEC|Ant cornea dystrophy NEC
C0155126|T047|PT|371.52|ICD9CM|Other anterior corneal dystrophies|Other anterior corneal dystrophies
C0018179|T047|AB|371.53|ICD9CM|Granular cornea dystrphy|Granular cornea dystrphy
C0018179|T047|PT|371.53|ICD9CM|Granular corneal dystrophy|Granular corneal dystrophy
C0155127|T047|AB|371.54|ICD9CM|Lattice cornea dystrophy|Lattice cornea dystrophy
C0155127|T047|PT|371.54|ICD9CM|Lattice corneal dystrophy|Lattice corneal dystrophy
C0024439|T047|AB|371.55|ICD9CM|Macular cornea dystrophy|Macular cornea dystrophy
C0024439|T047|PT|371.55|ICD9CM|Macular corneal dystrophy|Macular corneal dystrophy
C0155128|T047|PT|371.56|ICD9CM|Other stromal corneal dystrophies|Other stromal corneal dystrophies
C0155128|T047|AB|371.56|ICD9CM|Strom cornea dystrph NEC|Strom cornea dystrph NEC
C0544008|T047|AB|371.57|ICD9CM|Endothel cornea dystrphy|Endothel cornea dystrphy
C0544008|T047|PT|371.57|ICD9CM|Endothelial corneal dystrophy|Endothelial corneal dystrophy
C0155130|T047|PT|371.58|ICD9CM|Other posterior corneal dystrophies|Other posterior corneal dystrophies
C0155130|T047|AB|371.58|ICD9CM|Post cornea dystrphy NEC|Post cornea dystrphy NEC
C0022578|T047|HT|371.6|ICD9CM|Keratoconus|Keratoconus
C0022578|T047|AB|371.60|ICD9CM|Keratoconus NOS|Keratoconus NOS
C0022578|T047|PT|371.60|ICD9CM|Keratoconus, unspecified|Keratoconus, unspecified
C0155131|T047|AB|371.61|ICD9CM|Keratoconus, stable|Keratoconus, stable
C0155131|T047|PT|371.61|ICD9CM|Keratoconus, stable condition|Keratoconus, stable condition
C0339286|T047|AB|371.62|ICD9CM|Keratoconus, ac hydrops|Keratoconus, ac hydrops
C0339286|T047|PT|371.62|ICD9CM|Keratoconus, acute hydrops|Keratoconus, acute hydrops
C0155133|T190|HT|371.7|ICD9CM|Other corneal deformities|Other corneal deformities
C0339212|T190|AB|371.70|ICD9CM|Corneal deformity NOS|Corneal deformity NOS
C0339212|T190|PT|371.70|ICD9CM|Corneal deformity, unspecified|Corneal deformity, unspecified
C0155135|T047|AB|371.71|ICD9CM|Corneal ectasia|Corneal ectasia
C0155135|T047|PT|371.71|ICD9CM|Corneal ectasia|Corneal ectasia
C0155136|T190|AB|371.72|ICD9CM|Descemetocele|Descemetocele
C0155136|T190|PT|371.72|ICD9CM|Descemetocele|Descemetocele
C0152440|T047|AB|371.73|ICD9CM|Corneal staphyloma|Corneal staphyloma
C0152440|T047|PT|371.73|ICD9CM|Corneal staphyloma|Corneal staphyloma
C0155137|T047|HT|371.8|ICD9CM|Other corneal disorders|Other corneal disorders
C0155138|T047|AB|371.81|ICD9CM|Corneal anesthesia|Corneal anesthesia
C0155138|T047|PT|371.81|ICD9CM|Corneal anesthesia and hypoesthesia|Corneal anesthesia and hypoesthesia
C0375253|T020|PT|371.82|ICD9CM|Corneal disorder due to contact lens|Corneal disorder due to contact lens
C0375253|T020|AB|371.82|ICD9CM|Corneal dsdr contct lens|Corneal dsdr contct lens
C0155137|T047|AB|371.89|ICD9CM|Corneal disorder NEC|Corneal disorder NEC
C0155137|T047|PT|371.89|ICD9CM|Other corneal disorders|Other corneal disorders
C0010034|T047|AB|371.9|ICD9CM|Corneal disorder NOS|Corneal disorder NOS
C0010034|T047|PT|371.9|ICD9CM|Unspecified corneal disorder|Unspecified corneal disorder
C0009759|T047|HT|372|ICD9CM|Disorders of conjunctiva|Disorders of conjunctiva
C0155141|T047|HT|372.0|ICD9CM|Acute conjunctivitis|Acute conjunctivitis
C0155141|T047|AB|372.00|ICD9CM|Acute conjunctivitis NOS|Acute conjunctivitis NOS
C0155141|T047|PT|372.00|ICD9CM|Acute conjunctivitis, unspecified|Acute conjunctivitis, unspecified
C0155142|T047|AB|372.01|ICD9CM|Serous conjunctivitis|Serous conjunctivitis
C0155142|T047|PT|372.01|ICD9CM|Serous conjunctivitis, except viral|Serous conjunctivitis, except viral
C0155143|T047|AB|372.02|ICD9CM|Ac follic conjunctivitis|Ac follic conjunctivitis
C0155143|T047|PT|372.02|ICD9CM|Acute follicular conjunctivitis|Acute follicular conjunctivitis
C0029668|T047|AB|372.03|ICD9CM|Mucopur conjunctivit NEC|Mucopur conjunctivit NEC
C0029668|T047|PT|372.03|ICD9CM|Other mucopurulent conjunctivitis|Other mucopurulent conjunctivitis
C0155144|T047|AB|372.04|ICD9CM|Pseudomemb conjunctivit|Pseudomemb conjunctivit
C0155144|T047|PT|372.04|ICD9CM|Pseudomembranous conjunctivitis|Pseudomembranous conjunctivitis
C0001309|T047|AB|372.05|ICD9CM|Ac atopic conjunctivitis|Ac atopic conjunctivitis
C0001309|T047|PT|372.05|ICD9CM|Acute atopic conjunctivitis|Acute atopic conjunctivitis
C2712777|T047|AB|372.06|ICD9CM|Ac chem conjunctivitis|Ac chem conjunctivitis
C2712777|T047|PT|372.06|ICD9CM|Acute chemical conjunctivitis|Acute chemical conjunctivitis
C0155145|T047|HT|372.1|ICD9CM|Chronic conjunctivitis|Chronic conjunctivitis
C0155145|T047|AB|372.10|ICD9CM|Chr conjunctivitis NOS|Chr conjunctivitis NOS
C0155145|T047|PT|372.10|ICD9CM|Chronic conjunctivitis, unspecified|Chronic conjunctivitis, unspecified
C0155146|T047|AB|372.11|ICD9CM|Simpl chr conjunctivitis|Simpl chr conjunctivitis
C0155146|T047|PT|372.11|ICD9CM|Simple chronic conjunctivitis|Simple chronic conjunctivitis
C0155147|T047|AB|372.12|ICD9CM|Chr follic conjunctivit|Chr follic conjunctivit
C0155147|T047|PT|372.12|ICD9CM|Chronic follicular conjunctivitis|Chronic follicular conjunctivitis
C0009773|T047|AB|372.13|ICD9CM|Vernal conjunctivitis|Vernal conjunctivitis
C0009773|T047|PT|372.13|ICD9CM|Vernal conjunctivitis|Vernal conjunctivitis
C0029543|T047|AB|372.14|ICD9CM|Chr allrg conjunctiv NEC|Chr allrg conjunctiv NEC
C0029543|T047|PT|372.14|ICD9CM|Other chronic allergic conjunctivitis|Other chronic allergic conjunctivitis
C0155148|T047|AB|372.15|ICD9CM|Parasitic conjunctivitis|Parasitic conjunctivitis
C0155148|T047|PT|372.15|ICD9CM|Parasitic conjunctivitis|Parasitic conjunctivitis
C0005743|T047|HT|372.2|ICD9CM|Blepharoconjunctivitis|Blepharoconjunctivitis
C0005743|T047|AB|372.20|ICD9CM|Blepharoconjunctivit NOS|Blepharoconjunctivit NOS
C0005743|T047|PT|372.20|ICD9CM|Blepharoconjunctivitis, unspecified|Blepharoconjunctivitis, unspecified
C0155149|T047|AB|372.21|ICD9CM|Angular blepharoconjunct|Angular blepharoconjunct
C0155149|T047|PT|372.21|ICD9CM|Angular blepharoconjunctivitis|Angular blepharoconjunctivitis
C0155150|T047|AB|372.22|ICD9CM|Contact blepharoconjunct|Contact blepharoconjunct
C0155150|T047|PT|372.22|ICD9CM|Contact blepharoconjunctivitis|Contact blepharoconjunctivitis
C0029560|T047|HT|372.3|ICD9CM|Other and unspecified conjunctivitis|Other and unspecified conjunctivitis
C0009763|T047|AB|372.30|ICD9CM|Conjunctivitis NOS|Conjunctivitis NOS
C0009763|T047|PT|372.30|ICD9CM|Conjunctivitis, unspecified|Conjunctivitis, unspecified
C0155152|T047|AB|372.31|ICD9CM|Rosacea conjunctivitis|Rosacea conjunctivitis
C0155152|T047|PT|372.31|ICD9CM|Rosacea conjunctivitis|Rosacea conjunctivitis
C0155153|T047|PT|372.33|ICD9CM|Conjunctivitis in mucocutaneous disease|Conjunctivitis in mucocutaneous disease
C0155153|T047|AB|372.33|ICD9CM|Mucocutan dis conjunctiv|Mucocutan dis conjunctiv
C1328333|T047|PT|372.34|ICD9CM|Pingueculitis|Pingueculitis
C1328333|T047|AB|372.34|ICD9CM|Pingueculitis|Pingueculitis
C0029560|T047|AB|372.39|ICD9CM|Conjunctivitis NEC|Conjunctivitis NEC
C0029560|T047|PT|372.39|ICD9CM|Other conjunctivitis|Other conjunctivitis
C4520843|T047|HT|372.4|ICD9CM|Pterygium|Pterygium
C4520843|T047|AB|372.40|ICD9CM|Pterygium NOS|Pterygium NOS
C4520843|T047|PT|372.40|ICD9CM|Pterygium, unspecified|Pterygium, unspecified
C0155154|T047|AB|372.41|ICD9CM|Periph station pterygium|Periph station pterygium
C0155154|T047|PT|372.41|ICD9CM|Peripheral pterygium, stationary|Peripheral pterygium, stationary
C0155155|T047|AB|372.42|ICD9CM|Periph progess pterygium|Periph progess pterygium
C0155155|T047|PT|372.42|ICD9CM|Peripheral pterygium, progressive|Peripheral pterygium, progressive
C0155156|T047|AB|372.43|ICD9CM|Central pterygium|Central pterygium
C0155156|T047|PT|372.43|ICD9CM|Central pterygium|Central pterygium
C0155157|T047|AB|372.44|ICD9CM|Double pterygium|Double pterygium
C0155157|T047|PT|372.44|ICD9CM|Double pterygium|Double pterygium
C0155158|T047|AB|372.45|ICD9CM|Recurrent pterygium|Recurrent pterygium
C0155158|T047|PT|372.45|ICD9CM|Recurrent pterygium|Recurrent pterygium
C0155159|T020|HT|372.5|ICD9CM|Conjunctival degenerations and deposits|Conjunctival degenerations and deposits
C0155160|T047|AB|372.50|ICD9CM|Conjunctival degen NOS|Conjunctival degen NOS
C0155160|T047|PT|372.50|ICD9CM|Conjunctival degeneration, unspecified|Conjunctival degeneration, unspecified
C0152255|T047|AB|372.51|ICD9CM|Pinguecula|Pinguecula
C0152255|T047|PT|372.51|ICD9CM|Pinguecula|Pinguecula
C0155161|T047|AB|372.52|ICD9CM|Pseudopterygium|Pseudopterygium
C0155161|T047|PT|372.52|ICD9CM|Pseudopterygium|Pseudopterygium
C3665609|T047|AB|372.53|ICD9CM|Conjunctival xerosis|Conjunctival xerosis
C3665609|T047|PT|372.53|ICD9CM|Conjunctival xerosis|Conjunctival xerosis
C0155162|T020|AB|372.54|ICD9CM|Conjunctival concretions|Conjunctival concretions
C0155162|T020|PT|372.54|ICD9CM|Conjunctival concretions|Conjunctival concretions
C0155163|T047|AB|372.55|ICD9CM|Conjunctiva pigmentation|Conjunctiva pigmentation
C0155163|T047|PT|372.55|ICD9CM|Conjunctival pigmentations|Conjunctival pigmentations
C0162280|T047|AB|372.56|ICD9CM|Conjunctival deposits|Conjunctival deposits
C0162280|T047|PT|372.56|ICD9CM|Conjunctival deposits|Conjunctival deposits
C0155164|T020|HT|372.6|ICD9CM|Conjunctival scars|Conjunctival scars
C0155165|T047|AB|372.61|ICD9CM|Granuloma of conjunctiva|Granuloma of conjunctiva
C0155165|T047|PT|372.61|ICD9CM|Granuloma of conjunctiva|Granuloma of conjunctiva
C0155166|T047|AB|372.62|ICD9CM|Local conjunctiva adhes|Local conjunctiva adhes
C0155166|T047|PT|372.62|ICD9CM|Localized adhesions and strands of conjunctiva|Localized adhesions and strands of conjunctiva
C0152454|T046|AB|372.63|ICD9CM|Symblepharon|Symblepharon
C0152454|T046|PT|372.63|ICD9CM|Symblepharon|Symblepharon
C0155164|T020|AB|372.64|ICD9CM|Scarring of conjunctiva|Scarring of conjunctiva
C0155164|T020|PT|372.64|ICD9CM|Scarring of conjunctiva|Scarring of conjunctiva
C0155168|T047|HT|372.7|ICD9CM|Conjunctival vascular disorders and cysts|Conjunctival vascular disorders and cysts
C1761613|T033|AB|372.71|ICD9CM|Hyperemia of conjunctiva|Hyperemia of conjunctiva
C1761613|T033|PT|372.71|ICD9CM|Hyperemia of conjunctiva|Hyperemia of conjunctiva
C0009760|T046|AB|372.72|ICD9CM|Conjunctival hemorrhage|Conjunctival hemorrhage
C0009760|T046|PT|372.72|ICD9CM|Conjunctival hemorrhage|Conjunctival hemorrhage
C0151601|T046|AB|372.73|ICD9CM|Conjunctival edema|Conjunctival edema
C0151601|T046|PT|372.73|ICD9CM|Conjunctival edema|Conjunctival edema
C0042370|T190|AB|372.74|ICD9CM|Conjunctiva vasc anomaly|Conjunctiva vasc anomaly
C0042370|T190|PT|372.74|ICD9CM|Vascular abnormalities of conjunctiva|Vascular abnormalities of conjunctiva
C0155170|T047|AB|372.75|ICD9CM|Conjunctival cysts|Conjunctival cysts
C0155170|T047|PT|372.75|ICD9CM|Conjunctival cysts|Conjunctival cysts
C0155171|T047|HT|372.8|ICD9CM|Other disorders of conjunctiva|Other disorders of conjunctiva
C0878693|T047|AB|372.81|ICD9CM|Conjunctivochalasis|Conjunctivochalasis
C0878693|T047|PT|372.81|ICD9CM|Conjunctivochalasis|Conjunctivochalasis
C0155171|T047|AB|372.89|ICD9CM|Conjunctiva disorder NEC|Conjunctiva disorder NEC
C0155171|T047|PT|372.89|ICD9CM|Other disorders of conjunctiva|Other disorders of conjunctiva
C0009759|T047|AB|372.9|ICD9CM|Conjunctiva disorder NOS|Conjunctiva disorder NOS
C0009759|T047|PT|372.9|ICD9CM|Unspecified disorder of conjunctiva|Unspecified disorder of conjunctiva
C1812623|T047|HT|373|ICD9CM|Inflammation of eyelids|Inflammation of eyelids
C0005741|T047|HT|373.0|ICD9CM|Blepharitis|Blepharitis
C0005741|T047|AB|373.00|ICD9CM|Blepharitis NOS|Blepharitis NOS
C0005741|T047|PT|373.00|ICD9CM|Blepharitis, unspecified|Blepharitis, unspecified
C0155173|T047|AB|373.01|ICD9CM|Ulcerative blepharitis|Ulcerative blepharitis
C0155173|T047|PT|373.01|ICD9CM|Ulcerative blepharitis|Ulcerative blepharitis
C0155174|T047|AB|373.02|ICD9CM|Squamous blepharitis|Squamous blepharitis
C0155174|T047|PT|373.02|ICD9CM|Squamous blepharitis|Squamous blepharitis
C0019918|T047|HT|373.1|ICD9CM|Hordeolum and other deep inflammation of eyelid|Hordeolum and other deep inflammation of eyelid
C0019919|T047|AB|373.11|ICD9CM|Hordeolum externum|Hordeolum externum
C0019919|T047|PT|373.11|ICD9CM|Hordeolum externum|Hordeolum externum
C0085690|T047|AB|373.12|ICD9CM|Hordeolum internum|Hordeolum internum
C0085690|T047|PT|373.12|ICD9CM|Hordeolum internum|Hordeolum internum
C0155175|T047|AB|373.13|ICD9CM|Abscess of eyelid|Abscess of eyelid
C0155175|T047|PT|373.13|ICD9CM|Abscess of eyelid|Abscess of eyelid
C0007933|T047|AB|373.2|ICD9CM|Chalazion|Chalazion
C0007933|T047|PT|373.2|ICD9CM|Chalazion|Chalazion
C0155176|T047|HT|373.3|ICD9CM|Noninfectious dermatoses of eyelid|Noninfectious dermatoses of eyelid
C0155177|T047|AB|373.31|ICD9CM|Eczem dermatitis eyelid|Eczem dermatitis eyelid
C0155177|T047|PT|373.31|ICD9CM|Eczematous dermatitis of eyelid|Eczematous dermatitis of eyelid
C0155178|T047|PT|373.32|ICD9CM|Contact and allergic dermatitis of eyelid|Contact and allergic dermatitis of eyelid
C0155178|T047|AB|373.32|ICD9CM|Contact dermatit eyelid|Contact dermatit eyelid
C0155179|T047|AB|373.33|ICD9CM|Xeroderma of eyelid|Xeroderma of eyelid
C0155179|T047|PT|373.33|ICD9CM|Xeroderma of eyelid|Xeroderma of eyelid
C0155180|T047|AB|373.34|ICD9CM|Disc lup erythematos lid|Disc lup erythematos lid
C0155180|T047|PT|373.34|ICD9CM|Discoid lupus erythematosus of eyelid|Discoid lupus erythematosus of eyelid
C0155181|T047|AB|373.4|ICD9CM|Infect derm lid w deform|Infect derm lid w deform
C0155181|T047|PT|373.4|ICD9CM|Infective dermatitis of eyelid of types resulting in deformity|Infective dermatitis of eyelid of types resulting in deformity
C0155182|T047|AB|373.5|ICD9CM|Infec dermatitis lid NEC|Infec dermatitis lid NEC
C0155182|T047|PT|373.5|ICD9CM|Other infective dermatitis of eyelid|Other infective dermatitis of eyelid
C0155183|T047|AB|373.6|ICD9CM|Parasitic infest eyelid|Parasitic infest eyelid
C0155183|T047|PT|373.6|ICD9CM|Parasitic infestation of eyelid|Parasitic infestation of eyelid
C0155184|T047|AB|373.8|ICD9CM|Inflammation eyelid NEC|Inflammation eyelid NEC
C0155184|T047|PT|373.8|ICD9CM|Other inflammations of eyelids|Other inflammations of eyelids
C0005741|T047|AB|373.9|ICD9CM|Inflammation eyelid NOS|Inflammation eyelid NOS
C0005741|T047|PT|373.9|ICD9CM|Unspecified inflammation of eyelid|Unspecified inflammation of eyelid
C0155186|T047|HT|374|ICD9CM|Other disorders of eyelids|Other disorders of eyelids
C0339058|T047|HT|374.0|ICD9CM|Entropion and trichiasis of eyelid|Entropion and trichiasis of eyelid
C0014390|T047|AB|374.00|ICD9CM|Entropion NOS|Entropion NOS
C0014390|T047|PT|374.00|ICD9CM|Entropion, unspecified|Entropion, unspecified
C0155188|T047|AB|374.01|ICD9CM|Senile entropion|Senile entropion
C0155188|T047|PT|374.01|ICD9CM|Senile entropion|Senile entropion
C0155189|T047|AB|374.02|ICD9CM|Mechanical entropion|Mechanical entropion
C0155189|T047|PT|374.02|ICD9CM|Mechanical entropion|Mechanical entropion
C0155190|T047|AB|374.03|ICD9CM|Spastic entropion|Spastic entropion
C0155190|T047|PT|374.03|ICD9CM|Spastic entropion|Spastic entropion
C0155191|T047|AB|374.04|ICD9CM|Cicatricial entropion|Cicatricial entropion
C0155191|T047|PT|374.04|ICD9CM|Cicatricial entropion|Cicatricial entropion
C0271311|T047|PT|374.05|ICD9CM|Trichiasis of eyelid without entropion|Trichiasis of eyelid without entropion
C0271311|T047|AB|374.05|ICD9CM|Trichiasis w/o entropion|Trichiasis w/o entropion
C0013592|T047|HT|374.1|ICD9CM|Ectropion|Ectropion
C0013592|T047|AB|374.10|ICD9CM|Ectropion NOS|Ectropion NOS
C0013592|T047|PT|374.10|ICD9CM|Ectropion, unspecified|Ectropion, unspecified
C0155193|T047|AB|374.11|ICD9CM|Senile ectropion|Senile ectropion
C0155193|T047|PT|374.11|ICD9CM|Senile ectropion|Senile ectropion
C0155194|T047|AB|374.12|ICD9CM|Mechanical ectropion|Mechanical ectropion
C0155194|T047|PT|374.12|ICD9CM|Mechanical ectropion|Mechanical ectropion
C0155195|T047|AB|374.13|ICD9CM|Spastic ectropion|Spastic ectropion
C0155195|T047|PT|374.13|ICD9CM|Spastic ectropion|Spastic ectropion
C0155196|T047|AB|374.14|ICD9CM|Cicatricial ectropion|Cicatricial ectropion
C0155196|T047|PT|374.14|ICD9CM|Cicatricial ectropion|Cicatricial ectropion
C0152226|T047|HT|374.2|ICD9CM|Lagophthalmos|Lagophthalmos
C0152226|T047|AB|374.20|ICD9CM|Lagophthalmos NOS|Lagophthalmos NOS
C0152226|T047|PT|374.20|ICD9CM|Lagophthalmos, unspecified|Lagophthalmos, unspecified
C0155197|T047|AB|374.21|ICD9CM|Paralytic lagophthalmos|Paralytic lagophthalmos
C0155197|T047|PT|374.21|ICD9CM|Paralytic lagophthalmos|Paralytic lagophthalmos
C0155198|T047|AB|374.22|ICD9CM|Mechanical lagophthalmos|Mechanical lagophthalmos
C0155198|T047|PT|374.22|ICD9CM|Mechanical lagophthalmos|Mechanical lagophthalmos
C0155199|T047|AB|374.23|ICD9CM|Cicatricial lagophthalm|Cicatricial lagophthalm
C0155199|T047|PT|374.23|ICD9CM|Cicatricial lagophthalmos|Cicatricial lagophthalmos
C0005745|T047|HT|374.3|ICD9CM|Ptosis of eyelid|Ptosis of eyelid
C0005745|T047|AB|374.30|ICD9CM|Ptosis of eyelid NOS|Ptosis of eyelid NOS
C0005745|T047|PT|374.30|ICD9CM|Ptosis of eyelid, unspecified|Ptosis of eyelid, unspecified
C0392587|T033|AB|374.31|ICD9CM|Paralytic ptosis|Paralytic ptosis
C0392587|T033|PT|374.31|ICD9CM|Paralytic ptosis|Paralytic ptosis
C0155201|T046|AB|374.32|ICD9CM|Myogenic ptosis|Myogenic ptosis
C0155201|T046|PT|374.32|ICD9CM|Myogenic ptosis|Myogenic ptosis
C0155202|T020|AB|374.33|ICD9CM|Mechanical ptosis|Mechanical ptosis
C0155202|T020|PT|374.33|ICD9CM|Mechanical ptosis|Mechanical ptosis
C0005742|T047|AB|374.34|ICD9CM|Blepharochalasis|Blepharochalasis
C0005742|T047|PT|374.34|ICD9CM|Blepharochalasis|Blepharochalasis
C0155203|T047|HT|374.4|ICD9CM|Other disorders affecting eyelid function|Other disorders affecting eyelid function
C0155204|T184|AB|374.41|ICD9CM|Lid retraction or lag|Lid retraction or lag
C0155204|T184|PT|374.41|ICD9CM|Lid retraction or lag|Lid retraction or lag
C0266521|T047|AB|374.43|ICD9CM|Abnorm innervation synd|Abnorm innervation synd
C0266521|T047|PT|374.43|ICD9CM|Abnormal innervation syndrome of eyelid|Abnormal innervation syndrome of eyelid
C0155206|T047|PT|374.44|ICD9CM|Sensory disorders of eyelid|Sensory disorders of eyelid
C0155206|T047|AB|374.44|ICD9CM|Sensory disorders, lid|Sensory disorders, lid
C0155207|T047|PT|374.45|ICD9CM|Other sensorimotor disorders of eyelid|Other sensorimotor disorders of eyelid
C0155207|T047|AB|374.45|ICD9CM|Sensormotr disor lid NEC|Sensormotr disor lid NEC
C0005744|T019|AB|374.46|ICD9CM|Blepharophimosis|Blepharophimosis
C0005744|T019|PT|374.46|ICD9CM|Blepharophimosis|Blepharophimosis
C0155208|T046|HT|374.5|ICD9CM|Degenerative disorders of eyelid and periocular area|Degenerative disorders of eyelid and periocular area
C0155209|T047|AB|374.50|ICD9CM|Degen disorder NOS, lid|Degen disorder NOS, lid
C0155209|T047|PT|374.50|ICD9CM|Degenerative disorder of eyelid, unspecified|Degenerative disorder of eyelid, unspecified
C0155210|T047|AB|374.51|ICD9CM|Xanthelasma|Xanthelasma
C0155210|T047|PT|374.51|ICD9CM|Xanthelasma of eyelid|Xanthelasma of eyelid
C0155211|T047|AB|374.52|ICD9CM|Hyperpigmentation lid|Hyperpigmentation lid
C0155211|T047|PT|374.52|ICD9CM|Hyperpigmentation of eyelid|Hyperpigmentation of eyelid
C0155212|T047|AB|374.53|ICD9CM|Hypopigmentation lid|Hypopigmentation lid
C0155212|T047|PT|374.53|ICD9CM|Hypopigmentation of eyelid|Hypopigmentation of eyelid
C0155213|T047|AB|374.54|ICD9CM|Hypertrichosis of eyelid|Hypertrichosis of eyelid
C0155213|T047|PT|374.54|ICD9CM|Hypertrichosis of eyelid|Hypertrichosis of eyelid
C0155214|T047|AB|374.55|ICD9CM|Hypotrichosis of eyelid|Hypotrichosis of eyelid
C0155214|T047|PT|374.55|ICD9CM|Hypotrichosis of eyelid|Hypotrichosis of eyelid
C0155215|T047|AB|374.56|ICD9CM|Degen dis eyelid NEC|Degen dis eyelid NEC
C0155215|T047|PT|374.56|ICD9CM|Other degenerative disorders of skin affecting eyelid|Other degenerative disorders of skin affecting eyelid
C0155186|T047|HT|374.8|ICD9CM|Other disorders of eyelid|Other disorders of eyelid
C0155216|T046|AB|374.81|ICD9CM|Hemorrhage of eyelid|Hemorrhage of eyelid
C0155216|T046|PT|374.81|ICD9CM|Hemorrhage of eyelid|Hemorrhage of eyelid
C0162285|T046|AB|374.82|ICD9CM|Edema of eyelid|Edema of eyelid
C0162285|T046|PT|374.82|ICD9CM|Edema of eyelid|Edema of eyelid
C0155217|T047|AB|374.83|ICD9CM|Elephantiasis of eyelid|Elephantiasis of eyelid
C0155217|T047|PT|374.83|ICD9CM|Elephantiasis of eyelid|Elephantiasis of eyelid
C0155218|T047|AB|374.84|ICD9CM|Cysts of eyelids|Cysts of eyelids
C0155218|T047|PT|374.84|ICD9CM|Cysts of eyelids|Cysts of eyelids
C0155219|T190|PT|374.85|ICD9CM|Vascular anomalies of eyelid|Vascular anomalies of eyelid
C0155219|T190|AB|374.85|ICD9CM|Vascular anomaly, eyelid|Vascular anomaly, eyelid
C0339097|T047|AB|374.86|ICD9CM|Old foreign body, eyelid|Old foreign body, eyelid
C0339097|T047|PT|374.86|ICD9CM|Retained foreign body of eyelid|Retained foreign body of eyelid
C0423124|T033|AB|374.87|ICD9CM|Dermatochalasis|Dermatochalasis
C0423124|T033|PT|374.87|ICD9CM|Dermatochalasis|Dermatochalasis
C0155186|T047|AB|374.89|ICD9CM|Disorders of eyelid NEC|Disorders of eyelid NEC
C0155186|T047|PT|374.89|ICD9CM|Other disorders of eyelid|Other disorders of eyelid
C0015423|T047|AB|374.9|ICD9CM|Disorder of eyelid NOS|Disorder of eyelid NOS
C0015423|T047|PT|374.9|ICD9CM|Unspecified disorder of eyelid|Unspecified disorder of eyelid
C0022904|T047|HT|375|ICD9CM|Disorders of lacrimal system|Disorders of lacrimal system
C0155223|T047|HT|375.0|ICD9CM|Dacryoadenitis|Dacryoadenitis
C0155223|T047|AB|375.00|ICD9CM|Dacryoadenitis NOS|Dacryoadenitis NOS
C0155223|T047|PT|375.00|ICD9CM|Dacryoadenitis, unspecified|Dacryoadenitis, unspecified
C0149505|T047|AB|375.01|ICD9CM|Acute dacryoadenitis|Acute dacryoadenitis
C0149505|T047|PT|375.01|ICD9CM|Acute dacryoadenitis|Acute dacryoadenitis
C0155224|T047|AB|375.02|ICD9CM|Chronic dacryoadenitis|Chronic dacryoadenitis
C0155224|T047|PT|375.02|ICD9CM|Chronic dacryoadenitis|Chronic dacryoadenitis
C1300133|T047|AB|375.03|ICD9CM|Ch enlargmnt lacrim glnd|Ch enlargmnt lacrim glnd
C1300133|T047|PT|375.03|ICD9CM|Chronic enlargement of lacrimal gland|Chronic enlargement of lacrimal gland
C0155226|T047|HT|375.1|ICD9CM|Other disorders of lacrimal gland|Other disorders of lacrimal gland
C0155227|T184|AB|375.11|ICD9CM|Dacryops|Dacryops
C0155227|T184|PT|375.11|ICD9CM|Dacryops|Dacryops
C0155228|T047|AB|375.12|ICD9CM|Lacrimal gland cyst NEC|Lacrimal gland cyst NEC
C0155228|T047|PT|375.12|ICD9CM|Other lacrimal cysts and cystic degeneration|Other lacrimal cysts and cystic degeneration
C0155229|T047|AB|375.13|ICD9CM|Primary lacrimal atrophy|Primary lacrimal atrophy
C0155229|T047|PT|375.13|ICD9CM|Primary lacrimal atrophy|Primary lacrimal atrophy
C0339121|T020|AB|375.14|ICD9CM|Secondary lacrim atrophy|Secondary lacrim atrophy
C0339121|T020|PT|375.14|ICD9CM|Secondary lacrimal atrophy|Secondary lacrimal atrophy
C0043349|T047|AB|375.15|ICD9CM|Tear film insuffic NOS|Tear film insuffic NOS
C0043349|T047|PT|375.15|ICD9CM|Tear film insufficiency, unspecified|Tear film insufficiency, unspecified
C0155231|T047|PT|375.16|ICD9CM|Dislocation of lacrimal gland|Dislocation of lacrimal gland
C0155231|T047|AB|375.16|ICD9CM|Lacrimal gland dislocat|Lacrimal gland dislocat
C0152227|T047|HT|375.2|ICD9CM|Epiphora|Epiphora
C0152227|T047|AB|375.20|ICD9CM|Epiphora NOS|Epiphora NOS
C0152227|T047|PT|375.20|ICD9CM|Epiphora, unspecified as to cause|Epiphora, unspecified as to cause
C0155233|T047|AB|375.21|ICD9CM|Epiphora d/t excess tear|Epiphora d/t excess tear
C0155233|T047|PT|375.21|ICD9CM|Epiphora due to excess lacrimation|Epiphora due to excess lacrimation
C0155234|T047|AB|375.22|ICD9CM|Epiphora d/t insuf drain|Epiphora d/t insuf drain
C0155234|T047|PT|375.22|ICD9CM|Epiphora due to insufficient drainage|Epiphora due to insufficient drainage
C0339129|T047|HT|375.3|ICD9CM|Acute and unspecified inflammation of lacrimal passages|Acute and unspecified inflammation of lacrimal passages
C0010930|T047|AB|375.30|ICD9CM|Dacryocystitis NOS|Dacryocystitis NOS
C0010930|T047|PT|375.30|ICD9CM|Dacryocystitis, unspecified|Dacryocystitis, unspecified
C0339130|T047|AB|375.31|ICD9CM|Acute canaliculitis|Acute canaliculitis
C0339130|T047|PT|375.31|ICD9CM|Acute canaliculitis, lacrimal|Acute canaliculitis, lacrimal
C0155237|T047|AB|375.32|ICD9CM|Acute dacryocystitis|Acute dacryocystitis
C0155237|T047|PT|375.32|ICD9CM|Acute dacryocystitis|Acute dacryocystitis
C0155238|T047|AB|375.33|ICD9CM|Phlegmon dacryocystitis|Phlegmon dacryocystitis
C0155238|T047|PT|375.33|ICD9CM|Phlegmonous dacryocystitis|Phlegmonous dacryocystitis
C0155239|T047|HT|375.4|ICD9CM|Chronic inflammation of lacrimal passages|Chronic inflammation of lacrimal passages
C0155240|T047|AB|375.41|ICD9CM|Chronic canaliculitis|Chronic canaliculitis
C0155240|T047|PT|375.41|ICD9CM|Chronic canaliculitis|Chronic canaliculitis
C0149506|T047|AB|375.42|ICD9CM|Chronic dacryocystitis|Chronic dacryocystitis
C0149506|T047|PT|375.42|ICD9CM|Chronic dacryocystitis|Chronic dacryocystitis
C0155241|T047|AB|375.43|ICD9CM|Lacrimal mucocele|Lacrimal mucocele
C0155241|T047|PT|375.43|ICD9CM|Lacrimal mucocele|Lacrimal mucocele
C0155242|T047|HT|375.5|ICD9CM|Stenosis and insufficiency of lacrimal passages|Stenosis and insufficiency of lacrimal passages
C0155242|T190|HT|375.5|ICD9CM|Stenosis and insufficiency of lacrimal passages|Stenosis and insufficiency of lacrimal passages
C0155243|T047|PT|375.51|ICD9CM|Eversion of lacrimal punctum|Eversion of lacrimal punctum
C0155243|T047|AB|375.51|ICD9CM|Lacriml punctum eversion|Lacriml punctum eversion
C0155244|T047|AB|375.52|ICD9CM|Lacriml punctum stenosis|Lacriml punctum stenosis
C0155244|T047|PT|375.52|ICD9CM|Stenosis of lacrimal punctum|Stenosis of lacrimal punctum
C0155245|T190|AB|375.53|ICD9CM|Lacrim canalic stenosis|Lacrim canalic stenosis
C0155245|T190|PT|375.53|ICD9CM|Stenosis of lacrimal canaliculi|Stenosis of lacrimal canaliculi
C0155246|T190|AB|375.54|ICD9CM|Lacrimal sac stenosis|Lacrimal sac stenosis
C0155246|T190|PT|375.54|ICD9CM|Stenosis of lacrimal sac|Stenosis of lacrimal sac
C2745960|T047|AB|375.55|ICD9CM|Neonatal nasolacrml obst|Neonatal nasolacrml obst
C2745960|T047|PT|375.55|ICD9CM|Obstruction of nasolacrimal duct, neonatal|Obstruction of nasolacrimal duct, neonatal
C0155248|T020|AB|375.56|ICD9CM|Acq nasolacrml stenosis|Acq nasolacrml stenosis
C0155248|T020|PT|375.56|ICD9CM|Stenosis of nasolacrimal duct, acquired|Stenosis of nasolacrimal duct, acquired
C0155249|T047|AB|375.57|ICD9CM|Dacryolith|Dacryolith
C0155249|T047|PT|375.57|ICD9CM|Dacryolith|Dacryolith
C0155250|T020|HT|375.6|ICD9CM|Other changes of lacrimal passages|Other changes of lacrimal passages
C0155251|T190|AB|375.61|ICD9CM|Lacrimal fistula|Lacrimal fistula
C0155251|T190|PT|375.61|ICD9CM|Lacrimal fistula|Lacrimal fistula
C0155250|T020|AB|375.69|ICD9CM|Lacrim passge change NEC|Lacrim passge change NEC
C0155250|T020|PT|375.69|ICD9CM|Other changes of lacrimal passages|Other changes of lacrimal passages
C0155252|T047|HT|375.8|ICD9CM|Other disorders of lacrimal system|Other disorders of lacrimal system
C0155253|T047|PT|375.81|ICD9CM|Granuloma of lacrimal passages|Granuloma of lacrimal passages
C0155253|T047|AB|375.81|ICD9CM|Lacrim passage granuloma|Lacrim passage granuloma
C0155252|T047|AB|375.89|ICD9CM|Lacrimal syst dis NEC|Lacrimal syst dis NEC
C0155252|T047|PT|375.89|ICD9CM|Other disorders of lacrimal system|Other disorders of lacrimal system
C0022904|T047|AB|375.9|ICD9CM|Lacrimal syst dis NOS|Lacrimal syst dis NOS
C0022904|T047|PT|375.9|ICD9CM|Unspecified disorder of lacrimal system|Unspecified disorder of lacrimal system
C0029182|T047|HT|376|ICD9CM|Disorders of the orbit|Disorders of the orbit
C0155256|T033|HT|376.0|ICD9CM|Acute inflammation of orbit|Acute inflammation of orbit
C0155256|T033|AB|376.00|ICD9CM|Acute inflam NOS, orbit|Acute inflam NOS, orbit
C0155256|T033|PT|376.00|ICD9CM|Acute inflammation of orbit, unspecified|Acute inflammation of orbit, unspecified
C0149507|T047|AB|376.01|ICD9CM|Orbital cellulitis|Orbital cellulitis
C0149507|T047|PT|376.01|ICD9CM|Orbital cellulitis|Orbital cellulitis
C0155257|T047|AB|376.02|ICD9CM|Orbital periostitis|Orbital periostitis
C0155257|T047|PT|376.02|ICD9CM|Orbital periostitis|Orbital periostitis
C0155258|T047|AB|376.03|ICD9CM|Orbital osteomyelitis|Orbital osteomyelitis
C0155258|T047|PT|376.03|ICD9CM|Orbital osteomyelitis|Orbital osteomyelitis
C0155259|T047|AB|376.04|ICD9CM|Orbital tenonitis|Orbital tenonitis
C0155259|T047|PT|376.04|ICD9CM|Orbital tenonitis|Orbital tenonitis
C0155261|T047|HT|376.1|ICD9CM|Chronic inflammatory disorders of orbit|Chronic inflammatory disorders of orbit
C0155261|T047|AB|376.10|ICD9CM|Chr inflam NOS, orbit|Chr inflam NOS, orbit
C0155261|T047|PT|376.10|ICD9CM|Chronic inflammation of orbit, unspecified|Chronic inflammation of orbit, unspecified
C0155262|T047|AB|376.11|ICD9CM|Orbital granuloma|Orbital granuloma
C0155262|T047|PT|376.11|ICD9CM|Orbital granuloma|Orbital granuloma
C2350476|T047|AB|376.12|ICD9CM|Orbital myositis|Orbital myositis
C2350476|T047|PT|376.12|ICD9CM|Orbital myositis|Orbital myositis
C0155263|T047|AB|376.13|ICD9CM|Parasite infest, orbit|Parasite infest, orbit
C0155263|T047|PT|376.13|ICD9CM|Parasitic infestation of orbit|Parasitic infestation of orbit
C0155264|T047|HT|376.2|ICD9CM|Endocrine exophthalmos|Endocrine exophthalmos
C0155265|T047|AB|376.21|ICD9CM|Thyrotoxic exophthalmos|Thyrotoxic exophthalmos
C0155265|T047|PT|376.21|ICD9CM|Thyrotoxic exophthalmos|Thyrotoxic exophthalmos
C0152135|T047|AB|376.22|ICD9CM|Exophthalm ophthalmopleg|Exophthalm ophthalmopleg
C0152135|T047|PT|376.22|ICD9CM|Exophthalmic ophthalmoplegia|Exophthalmic ophthalmoplegia
C0155266|T047|HT|376.3|ICD9CM|Other exophthalmic conditions|Other exophthalmic conditions
C0015300|T047|AB|376.30|ICD9CM|Exophthalmos NOS|Exophthalmos NOS
C0015300|T047|PT|376.30|ICD9CM|Exophthalmos, unspecified|Exophthalmos, unspecified
C0155267|T047|AB|376.31|ICD9CM|Constant exophthalmos|Constant exophthalmos
C0155267|T047|PT|376.31|ICD9CM|Constant exophthalmos|Constant exophthalmos
C0155268|T046|AB|376.32|ICD9CM|Orbital hemorrhage|Orbital hemorrhage
C0155268|T046|PT|376.32|ICD9CM|Orbital hemorrhage|Orbital hemorrhage
C0424813|T046|AB|376.33|ICD9CM|Orbital edema|Orbital edema
C0424813|T046|PT|376.33|ICD9CM|Orbital edema or congestion|Orbital edema or congestion
C0155270|T047|PT|376.34|ICD9CM|Intermittent exophthalmos|Intermittent exophthalmos
C0155270|T047|AB|376.34|ICD9CM|Intermittnt exophthalmos|Intermittnt exophthalmos
C0155271|T047|AB|376.35|ICD9CM|Pulsating exophthalmos|Pulsating exophthalmos
C0155271|T047|PT|376.35|ICD9CM|Pulsating exophthalmos|Pulsating exophthalmos
C0155272|T047|PT|376.36|ICD9CM|Lateral displacement of globe|Lateral displacement of globe
C0155272|T047|AB|376.36|ICD9CM|Lateral globe displacmnt|Lateral globe displacmnt
C0162019|T190|HT|376.4|ICD9CM|Deformity of orbit|Deformity of orbit
C0162019|T190|AB|376.40|ICD9CM|Deformity of orbit NOS|Deformity of orbit NOS
C0162019|T190|PT|376.40|ICD9CM|Deformity of orbit, unspecified|Deformity of orbit, unspecified
C0020534|T033|AB|376.41|ICD9CM|Hypertelorism of orbit|Hypertelorism of orbit
C0020534|T033|PT|376.41|ICD9CM|Hypertelorism of orbit|Hypertelorism of orbit
C0155275|T047|AB|376.42|ICD9CM|Exostosis of orbit|Exostosis of orbit
C0155275|T047|PT|376.42|ICD9CM|Exostosis of orbit|Exostosis of orbit
C0155276|T020|PT|376.43|ICD9CM|Local deformities of orbit due to bone disease|Local deformities of orbit due to bone disease
C0155276|T020|AB|376.43|ICD9CM|Orbt deform d/t bone dis|Orbt deform d/t bone dis
C0155277|T190|AB|376.44|ICD9CM|Craniofacial-orbit defor|Craniofacial-orbit defor
C0155277|T190|PT|376.44|ICD9CM|Orbital deformities associated with craniofacial deformities|Orbital deformities associated with craniofacial deformities
C0155278|T046|AB|376.45|ICD9CM|Atrophy of orbit|Atrophy of orbit
C0155278|T046|PT|376.45|ICD9CM|Atrophy of orbit|Atrophy of orbit
C0155279|T047|AB|376.46|ICD9CM|Enlargement of orbit|Enlargement of orbit
C0155279|T047|PT|376.46|ICD9CM|Enlargement of orbit|Enlargement of orbit
C0155280|T020|PT|376.47|ICD9CM|Deformity of orbit due to trauma or surgery|Deformity of orbit due to trauma or surgery
C0155280|T020|AB|376.47|ICD9CM|Orbit deform d/t trauma|Orbit deform d/t trauma
C0014306|T047|HT|376.5|ICD9CM|Enophthalmos|Enophthalmos
C0014306|T047|AB|376.50|ICD9CM|Enophthalmos NOS|Enophthalmos NOS
C0014306|T047|PT|376.50|ICD9CM|Enophthalmos, unspecified as to cause|Enophthalmos, unspecified as to cause
C0155281|T047|AB|376.51|ICD9CM|Enophth d/t orbit atrphy|Enophth d/t orbit atrphy
C0155281|T047|PT|376.51|ICD9CM|Enophthalmos due to atrophy of orbital tissue|Enophthalmos due to atrophy of orbital tissue
C0155282|T020|AB|376.52|ICD9CM|Enophthalmos d/t trauma|Enophthalmos d/t trauma
C0155282|T020|PT|376.52|ICD9CM|Enophthalmos due to trauma or surgery|Enophthalmos due to trauma or surgery
C0155283|T020|AB|376.6|ICD9CM|Old foreign body, orbit|Old foreign body, orbit
C0155283|T020|PT|376.6|ICD9CM|Retained (old) foreign body following penetrating wound of orbit|Retained (old) foreign body following penetrating wound of orbit
C0155284|T047|HT|376.8|ICD9CM|Other orbital disorders|Other orbital disorders
C0155285|T047|AB|376.81|ICD9CM|Orbital cysts|Orbital cysts
C0155285|T047|PT|376.81|ICD9CM|Orbital cysts|Orbital cysts
C0155286|T047|AB|376.82|ICD9CM|Extraocul muscl myopathy|Extraocul muscl myopathy
C0155286|T047|PT|376.82|ICD9CM|Myopathy of extraocular muscles|Myopathy of extraocular muscles
C2609444|T047|AB|376.89|ICD9CM|Orbital disorders NEC|Orbital disorders NEC
C2609444|T047|PT|376.89|ICD9CM|Other orbital disorders|Other orbital disorders
C0029182|T047|AB|376.9|ICD9CM|Orbital disorder NOS|Orbital disorder NOS
C0029182|T047|PT|376.9|ICD9CM|Unspecified disorder of orbit|Unspecified disorder of orbit
C1533675|T047|HT|377|ICD9CM|Disorders of optic nerve and visual pathways|Disorders of optic nerve and visual pathways
C0030353|T047|HT|377.0|ICD9CM|Papilledema|Papilledema
C0030353|T047|AB|377.00|ICD9CM|Papilledema NOS|Papilledema NOS
C0030353|T047|PT|377.00|ICD9CM|Papilledema, unspecified|Papilledema, unspecified
C0155288|T047|PT|377.01|ICD9CM|Papilledema associated with increased intracranial pressure|Papilledema associated with increased intracranial pressure
C0155288|T047|AB|377.01|ICD9CM|Papilledema w incr press|Papilledema w incr press
C1827466|T047|PT|377.02|ICD9CM|Papilledema associated with decreased ocular pressure|Papilledema associated with decreased ocular pressure
C1827466|T047|AB|377.02|ICD9CM|Papilledema w decr press|Papilledema w decr press
C0155290|T047|PT|377.03|ICD9CM|Papilledema associated with retinal disorder|Papilledema associated with retinal disorder
C0155290|T047|AB|377.03|ICD9CM|Papilledema w retina dis|Papilledema w retina dis
C0152112|T047|PT|377.04|ICD9CM|Foster-Kennedy syndrome|Foster-Kennedy syndrome
C0152112|T047|AB|377.04|ICD9CM|Foster-kennedy syndrome|Foster-kennedy syndrome
C0029124|T047|HT|377.1|ICD9CM|Optic atrophy|Optic atrophy
C0029124|T047|AB|377.10|ICD9CM|Optic atrophy NOS|Optic atrophy NOS
C0029124|T047|PT|377.10|ICD9CM|Optic atrophy, unspecified|Optic atrophy, unspecified
C0155291|T047|AB|377.11|ICD9CM|Primary optic atrophy|Primary optic atrophy
C0155291|T047|PT|377.11|ICD9CM|Primary optic atrophy|Primary optic atrophy
C0155292|T047|AB|377.12|ICD9CM|Postinflam optic atrophy|Postinflam optic atrophy
C0155292|T047|PT|377.12|ICD9CM|Postinflammatory optic atrophy|Postinflammatory optic atrophy
C0155293|T047|PT|377.13|ICD9CM|Optic atrophy associated with retinal dystrophies|Optic atrophy associated with retinal dystrophies
C0155293|T047|AB|377.13|ICD9CM|Optic atrph w retin dyst|Optic atrph w retin dyst
C0271342|T047|AB|377.14|ICD9CM|Cupping of optic disc|Cupping of optic disc
C0271342|T047|PT|377.14|ICD9CM|Glaucomatous atrophy [cupping] of optic disc|Glaucomatous atrophy [cupping] of optic disc
C0155295|T047|AB|377.15|ICD9CM|Partial optic atrophy|Partial optic atrophy
C0155295|T047|PT|377.15|ICD9CM|Partial optic atrophy|Partial optic atrophy
C0029125|T047|AB|377.16|ICD9CM|Hereditary optic atrophy|Hereditary optic atrophy
C0029125|T047|PT|377.16|ICD9CM|Hereditary optic atrophy|Hereditary optic atrophy
C0155296|T047|HT|377.2|ICD9CM|Other disorders of optic disc|Other disorders of optic disc
C0029128|T047|AB|377.21|ICD9CM|Drusen of optic disc|Drusen of optic disc
C0029128|T047|PT|377.21|ICD9CM|Drusen of optic disc|Drusen of optic disc
C0155298|T047|AB|377.22|ICD9CM|Crater-like hole op disc|Crater-like hole op disc
C0155298|T047|PT|377.22|ICD9CM|Crater-like holes of optic disc|Crater-like holes of optic disc
C0155299|T047|AB|377.23|ICD9CM|Coloboma of optic disc|Coloboma of optic disc
C0155299|T047|PT|377.23|ICD9CM|Coloboma of optic disc|Coloboma of optic disc
C0155300|T047|AB|377.24|ICD9CM|Pseudopapilledema|Pseudopapilledema
C0155300|T047|PT|377.24|ICD9CM|Pseudopapilledema|Pseudopapilledema
C0029134|T047|HT|377.3|ICD9CM|Optic neuritis|Optic neuritis
C0029134|T047|AB|377.30|ICD9CM|Optic neuritis NOS|Optic neuritis NOS
C0029134|T047|PT|377.30|ICD9CM|Optic neuritis, unspecified|Optic neuritis, unspecified
C0030353|T047|AB|377.31|ICD9CM|Optic papillitis|Optic papillitis
C0030353|T047|PT|377.31|ICD9CM|Optic papillitis|Optic papillitis
C0155301|T047|AB|377.32|ICD9CM|Retrobulbar neuritis|Retrobulbar neuritis
C0155301|T047|PT|377.32|ICD9CM|Retrobulbar neuritis (acute)|Retrobulbar neuritis (acute)
C0155302|T047|AB|377.33|ICD9CM|Nutrition optc neuropthy|Nutrition optc neuropthy
C0155302|T047|PT|377.33|ICD9CM|Nutritional optic neuropathy|Nutritional optic neuropathy
C0155303|T047|AB|377.34|ICD9CM|Toxic optic neuropathy|Toxic optic neuropathy
C0155303|T047|PT|377.34|ICD9CM|Toxic optic neuropathy|Toxic optic neuropathy
C0029681|T047|AB|377.39|ICD9CM|Optic neuritis NEC|Optic neuritis NEC
C0029681|T047|PT|377.39|ICD9CM|Other optic neuritis|Other optic neuritis
C0155304|T047|HT|377.4|ICD9CM|Other disorders of optic nerve|Other disorders of optic nerve
C0155305|T047|PT|377.41|ICD9CM|Ischemic optic neuropathy|Ischemic optic neuropathy
C0155305|T047|AB|377.41|ICD9CM|Ischemic optic neuropthy|Ischemic optic neuropthy
C0155306|T046|PT|377.42|ICD9CM|Hemorrhage in optic nerve sheaths|Hemorrhage in optic nerve sheaths
C0155306|T046|AB|377.42|ICD9CM|Optic nerve sheath hemor|Optic nerve sheath hemor
C0338502|T047|PT|377.43|ICD9CM|Optic nerve hypoplasia|Optic nerve hypoplasia
C0338502|T047|AB|377.43|ICD9CM|Optic nerve hypoplasia|Optic nerve hypoplasia
C0155304|T047|AB|377.49|ICD9CM|Optic nerve disorder NEC|Optic nerve disorder NEC
C0155304|T047|PT|377.49|ICD9CM|Other disorders of optic nerve|Other disorders of optic nerve
C0155307|T047|HT|377.5|ICD9CM|Disorders of optic chiasm|Disorders of optic chiasm
C0155308|T047|PT|377.51|ICD9CM|Disorders of optic chiasm associated with pituitary neoplasms and disorders|Disorders of optic chiasm associated with pituitary neoplasms and disorders
C0155308|T047|AB|377.51|ICD9CM|Opt chiasm w pituit dis|Opt chiasm w pituit dis
C2004477|T047|PT|377.52|ICD9CM|Disorders of optic chiasm associated with other neoplasms|Disorders of optic chiasm associated with other neoplasms
C2004477|T047|AB|377.52|ICD9CM|Opt chiasm dis/neopl NEC|Opt chiasm dis/neopl NEC
C3665440|T047|PT|377.53|ICD9CM|Disorders of optic chiasm associated with vascular disorders|Disorders of optic chiasm associated with vascular disorders
C3665440|T047|AB|377.53|ICD9CM|Opt chiasm w vascul dis|Opt chiasm w vascul dis
C0155311|T047|PT|377.54|ICD9CM|Disorders of optic chiasm associated with inflammatory disorders|Disorders of optic chiasm associated with inflammatory disorders
C0155311|T047|AB|377.54|ICD9CM|Op chiasm dis w infl dis|Op chiasm dis w infl dis
C0155312|T047|HT|377.6|ICD9CM|Disorders of other visual pathways|Disorders of other visual pathways
C0155313|T047|PT|377.61|ICD9CM|Disorders of other visual pathways associated with neoplasms|Disorders of other visual pathways associated with neoplasms
C0155313|T047|AB|377.61|ICD9CM|Vis path dis w neoplasms|Vis path dis w neoplasms
C0155314|T047|PT|377.62|ICD9CM|Disorders of other visual pathways associated with vascular disorders|Disorders of other visual pathways associated with vascular disorders
C0155314|T047|AB|377.62|ICD9CM|Vis path dis w vasc dis|Vis path dis w vasc dis
C0155315|T047|PT|377.63|ICD9CM|Disorders of other visual pathways associated with inflammatory disorders|Disorders of other visual pathways associated with inflammatory disorders
C0155315|T047|AB|377.63|ICD9CM|Vis path dis w infl dis|Vis path dis w infl dis
C0234398|T047|HT|377.7|ICD9CM|Disorders of visual cortex|Disorders of visual cortex
C3665441|T047|PT|377.71|ICD9CM|Disorders of visual cortex associated with neoplasms|Disorders of visual cortex associated with neoplasms
C3665441|T047|AB|377.71|ICD9CM|Vis cortx dis w neoplasm|Vis cortx dis w neoplasm
C3665442|T047|PT|377.72|ICD9CM|Disorders of visual cortex associated with vascular disorders|Disorders of visual cortex associated with vascular disorders
C3665442|T047|AB|377.72|ICD9CM|Vis cortx dis w vasc dis|Vis cortx dis w vasc dis
C3665443|T047|PT|377.73|ICD9CM|Disorders of visual cortex associated with inflammatory disorders|Disorders of visual cortex associated with inflammatory disorders
C3665443|T047|AB|377.73|ICD9CM|Vis cortex dis w inflam|Vis cortex dis w inflam
C0155320|T047|AB|377.75|ICD9CM|Cortical blindness|Cortical blindness
C0155320|T047|PT|377.75|ICD9CM|Cortical blindness|Cortical blindness
C1533675|T047|AB|377.9|ICD9CM|Optic nerve disorder NOS|Optic nerve disorder NOS
C1533675|T047|PT|377.9|ICD9CM|Unspecified disorder of optic nerve and visual pathways|Unspecified disorder of optic nerve and visual pathways
C0038380|T047|HT|378|ICD9CM|Strabismus and other disorders of binocular eye movements|Strabismus and other disorders of binocular eye movements
C0014877|T047|HT|378.0|ICD9CM|Esotropia|Esotropia
C0014877|T047|AB|378.00|ICD9CM|Esotropia NOS|Esotropia NOS
C0014877|T047|PT|378.00|ICD9CM|Esotropia, unspecified|Esotropia, unspecified
C0152204|T047|AB|378.01|ICD9CM|Monocular esotropia|Monocular esotropia
C0152204|T047|PT|378.01|ICD9CM|Monocular esotropia|Monocular esotropia
C0155322|T047|AB|378.02|ICD9CM|Monoc esotrop w a pattrn|Monoc esotrop w a pattrn
C0155322|T047|PT|378.02|ICD9CM|Monocular esotropia with A pattern|Monocular esotropia with A pattern
C0155323|T047|AB|378.03|ICD9CM|Monoc esotrop w v pattrn|Monoc esotrop w v pattrn
C0155323|T047|PT|378.03|ICD9CM|Monocular esotropia with V pattern|Monocular esotropia with V pattern
C0155324|T047|AB|378.04|ICD9CM|Monoc esotrop w x/y pat|Monoc esotrop w x/y pat
C0155324|T047|PT|378.04|ICD9CM|Monocular esotropia with other noncomitancies|Monocular esotropia with other noncomitancies
C0152205|T047|AB|378.05|ICD9CM|Alternating esotropia|Alternating esotropia
C0152205|T047|PT|378.05|ICD9CM|Alternating esotropia|Alternating esotropia
C0155325|T047|AB|378.06|ICD9CM|Alt esotropia w a pattrn|Alt esotropia w a pattrn
C0155325|T047|PT|378.06|ICD9CM|Alternating esotropia with A pattern|Alternating esotropia with A pattern
C0155326|T047|AB|378.07|ICD9CM|Alt esotropia w v pattrn|Alt esotropia w v pattrn
C0155326|T047|PT|378.07|ICD9CM|Alternating esotropia with V pattern|Alternating esotropia with V pattern
C0155327|T047|AB|378.08|ICD9CM|Alt esotrop w x/y pattrn|Alt esotrop w x/y pattrn
C0155327|T047|PT|378.08|ICD9CM|Alternating esotropia with other noncomitancies|Alternating esotropia with other noncomitancies
C0015310|T047|HT|378.1|ICD9CM|Exotropia|Exotropia
C0015310|T047|AB|378.10|ICD9CM|Exotropia NOS|Exotropia NOS
C0015310|T047|PT|378.10|ICD9CM|Exotropia, unspecified|Exotropia, unspecified
C0152206|T047|AB|378.11|ICD9CM|Monocular exotropia|Monocular exotropia
C0152206|T047|PT|378.11|ICD9CM|Monocular exotropia|Monocular exotropia
C0155328|T047|AB|378.12|ICD9CM|Monoc exotrop w a pattrn|Monoc exotrop w a pattrn
C0155328|T047|PT|378.12|ICD9CM|Monocular exotropia with A pattern|Monocular exotropia with A pattern
C0155329|T047|AB|378.13|ICD9CM|Monoc exotrop w v pattrn|Monoc exotrop w v pattrn
C0155329|T047|PT|378.13|ICD9CM|Monocular exotropia with V pattern|Monocular exotropia with V pattern
C0155330|T047|AB|378.14|ICD9CM|Monoc exotrop w x/y pat|Monoc exotrop w x/y pat
C0155330|T047|PT|378.14|ICD9CM|Monocular exotropia with other noncomitancies|Monocular exotropia with other noncomitancies
C0152207|T047|AB|378.15|ICD9CM|Alternating exotropia|Alternating exotropia
C0152207|T047|PT|378.15|ICD9CM|Alternating exotropia|Alternating exotropia
C0155331|T047|AB|378.16|ICD9CM|Alt exotropia w a pattrn|Alt exotropia w a pattrn
C0155331|T047|PT|378.16|ICD9CM|Alternating exotropia with A pattern|Alternating exotropia with A pattern
C0155332|T047|AB|378.17|ICD9CM|Alt exotropia w v pattrn|Alt exotropia w v pattrn
C0155332|T047|PT|378.17|ICD9CM|Alternating exotropia with V pattern|Alternating exotropia with V pattern
C0155333|T047|AB|378.18|ICD9CM|Alt exotrop w x/y pattrn|Alt exotrop w x/y pattrn
C0155333|T047|PT|378.18|ICD9CM|Alternating exotropia with other noncomitancies|Alternating exotropia with other noncomitancies
C0152210|T047|HT|378.2|ICD9CM|Intermittent heterotropia|Intermittent heterotropia
C0152210|T047|AB|378.20|ICD9CM|Intermit heterotrop NOS|Intermit heterotrop NOS
C0152210|T047|PT|378.20|ICD9CM|Intermittent heterotropia, unspecified|Intermittent heterotropia, unspecified
C0152211|T047|AB|378.21|ICD9CM|Intermit monoc esotropia|Intermit monoc esotropia
C0152211|T047|PT|378.21|ICD9CM|Intermittent esotropia, monocular|Intermittent esotropia, monocular
C0152212|T047|AB|378.22|ICD9CM|Intermit altrn esotropia|Intermit altrn esotropia
C0152212|T047|PT|378.22|ICD9CM|Intermittent esotropia, alternating|Intermittent esotropia, alternating
C0152213|T047|AB|378.23|ICD9CM|Intermit monoc exotropia|Intermit monoc exotropia
C0152213|T047|PT|378.23|ICD9CM|Intermittent exotropia, monocular|Intermittent exotropia, monocular
C0152214|T047|AB|378.24|ICD9CM|Intermit altrn exotropia|Intermit altrn exotropia
C0152214|T047|PT|378.24|ICD9CM|Intermittent exotropia, alternating|Intermittent exotropia, alternating
C0155334|T047|HT|378.3|ICD9CM|Other and unspecified heterotropia|Other and unspecified heterotropia
C0038379|T047|AB|378.30|ICD9CM|Heterotropia NOS|Heterotropia NOS
C0038379|T047|PT|378.30|ICD9CM|Heterotropia, unspecified|Heterotropia, unspecified
C0020575|T047|AB|378.31|ICD9CM|Hypertropia|Hypertropia
C0020575|T047|PT|378.31|ICD9CM|Hypertropia|Hypertropia
C0152208|T047|AB|378.32|ICD9CM|Hypotropia|Hypotropia
C0152208|T047|PT|378.32|ICD9CM|Hypotropia|Hypotropia
C0152209|T047|AB|378.33|ICD9CM|Cyclotropia|Cyclotropia
C0152209|T047|PT|378.33|ICD9CM|Cyclotropia|Cyclotropia
C0339611|T047|AB|378.34|ICD9CM|Monofixation syndrome|Monofixation syndrome
C0339611|T047|PT|378.34|ICD9CM|Monofixation syndrome|Monofixation syndrome
C0155336|T047|PT|378.35|ICD9CM|Accommodative component in esotropia|Accommodative component in esotropia
C0155336|T047|AB|378.35|ICD9CM|Accommodative esotropia|Accommodative esotropia
C4721400|T047|HT|378.4|ICD9CM|Heterophoria|Heterophoria
C4721400|T047|AB|378.40|ICD9CM|Heterophoria NOS|Heterophoria NOS
C4721400|T047|PT|378.40|ICD9CM|Heterophoria, unspecified|Heterophoria, unspecified
C0152216|T047|AB|378.41|ICD9CM|Esophoria|Esophoria
C0152216|T047|PT|378.41|ICD9CM|Esophoria|Esophoria
C0152217|T047|AB|378.42|ICD9CM|Exophoria|Exophoria
C0152217|T047|PT|378.42|ICD9CM|Exophoria|Exophoria
C0152218|T047|AB|378.43|ICD9CM|Vertical heterophoria|Vertical heterophoria
C0152218|T047|PT|378.43|ICD9CM|Vertical heterophoria|Vertical heterophoria
C0152219|T047|AB|378.44|ICD9CM|Cyclophoria|Cyclophoria
C0152219|T047|PT|378.44|ICD9CM|Cyclophoria|Cyclophoria
C0152220|T047|AB|378.45|ICD9CM|Alternating hyperphoria|Alternating hyperphoria
C0152220|T047|PT|378.45|ICD9CM|Alternating hyperphoria|Alternating hyperphoria
C0152221|T047|HT|378.5|ICD9CM|Paralytic strabismus|Paralytic strabismus
C0152221|T047|AB|378.50|ICD9CM|Paralytic strabismus NOS|Paralytic strabismus NOS
C0152221|T047|PT|378.50|ICD9CM|Paralytic strabismus, unspecified|Paralytic strabismus, unspecified
C0271370|T047|AB|378.51|ICD9CM|Partial third nerv palsy|Partial third nerv palsy
C0271370|T047|PT|378.51|ICD9CM|Third or oculomotor nerve palsy, partial|Third or oculomotor nerve palsy, partial
C0271371|T047|PT|378.52|ICD9CM|Third or oculomotor nerve palsy, total|Third or oculomotor nerve palsy, total
C0271371|T047|AB|378.52|ICD9CM|Total third nerve palsy|Total third nerve palsy
C0271375|T047|AB|378.53|ICD9CM|Fourth nerve palsy|Fourth nerve palsy
C0271375|T047|PT|378.53|ICD9CM|Fourth or trochlear nerve palsy|Fourth or trochlear nerve palsy
C4551519|T047|AB|378.54|ICD9CM|Sixth nerve palsy|Sixth nerve palsy
C4551519|T047|PT|378.54|ICD9CM|Sixth or abducens nerve palsy|Sixth or abducens nerve palsy
C0162292|T047|AB|378.55|ICD9CM|External ophthalmoplegia|External ophthalmoplegia
C0162292|T047|PT|378.55|ICD9CM|External ophthalmoplegia|External ophthalmoplegia
C0155338|T047|AB|378.56|ICD9CM|Total ophthalmoplegia|Total ophthalmoplegia
C0155338|T047|PT|378.56|ICD9CM|Total ophthalmoplegia|Total ophthalmoplegia
C0152223|T047|HT|378.6|ICD9CM|Mechanical strabismus|Mechanical strabismus
C0152223|T047|AB|378.60|ICD9CM|Mechanical strabism NOS|Mechanical strabism NOS
C0152223|T047|PT|378.60|ICD9CM|Mechanical strabismus, unspecified|Mechanical strabismus, unspecified
C0155339|T047|PT|378.61|ICD9CM|Brown's (tendon) sheath syndrome|Brown's (tendon) sheath syndrome
C0155339|T047|AB|378.61|ICD9CM|Brown's sheath syndrome|Brown's sheath syndrome
C0155340|T047|AB|378.62|ICD9CM|Mech strab d/t muscl dis|Mech strab d/t muscl dis
C0155340|T047|PT|378.62|ICD9CM|Mechanical strabismus from other musculofascial disorders|Mechanical strabismus from other musculofascial disorders
C0155341|T047|PT|378.63|ICD9CM|Limited duction associated with other conditions|Limited duction associated with other conditions
C0155341|T047|AB|378.63|ICD9CM|Mech strab w oth conditn|Mech strab w oth conditn
C0029831|T047|HT|378.7|ICD9CM|Other specified strabismus|Other specified strabismus
C0013261|T047|AB|378.71|ICD9CM|Duane's syndrome|Duane's syndrome
C0013261|T047|PT|378.71|ICD9CM|Duane's syndrome|Duane's syndrome
C0162674|T047|AB|378.72|ICD9CM|Prog ext ophthalmoplegia|Prog ext ophthalmoplegia
C0162674|T047|PT|378.72|ICD9CM|Progressive external ophthalmoplegia|Progressive external ophthalmoplegia
C0155342|T047|AB|378.73|ICD9CM|Neuromuscle dis strabism|Neuromuscle dis strabism
C0155342|T047|PT|378.73|ICD9CM|Strabismus in other neuromuscular disorders|Strabismus in other neuromuscular disorders
C0155343|T047|HT|378.8|ICD9CM|Other disorders of binocular eye movements|Other disorders of binocular eye movements
C0702143|T047|AB|378.81|ICD9CM|Palsy of conjugate gaze|Palsy of conjugate gaze
C0702143|T047|PT|378.81|ICD9CM|Palsy of conjugate gaze|Palsy of conjugate gaze
C0155344|T184|AB|378.82|ICD9CM|Spasm of conjugate gaze|Spasm of conjugate gaze
C0155344|T184|PT|378.82|ICD9CM|Spasm of conjugate gaze|Spasm of conjugate gaze
C0155345|T047|AB|378.83|ICD9CM|Convergenc insufficiency|Convergenc insufficiency
C0155345|T047|PT|378.83|ICD9CM|Convergence insufficiency or palsy|Convergence insufficiency or palsy
C0155346|T047|AB|378.84|ICD9CM|Convergence excess|Convergence excess
C0155346|T047|PT|378.84|ICD9CM|Convergence excess or spasm|Convergence excess or spasm
C0155347|T184|AB|378.85|ICD9CM|Anomalies of divergence|Anomalies of divergence
C0155347|T184|PT|378.85|ICD9CM|Anomalies of divergence|Anomalies of divergence
C0152134|T047|AB|378.86|ICD9CM|Internucl ophthalmopleg|Internucl ophthalmopleg
C0152134|T047|PT|378.86|ICD9CM|Internuclear ophthalmoplegia|Internuclear ophthalmoplegia
C0733455|T047|PT|378.87|ICD9CM|Other dissociated deviation of eye movements|Other dissociated deviation of eye movements
C0733455|T047|AB|378.87|ICD9CM|Skew deviation, eye|Skew deviation, eye
C0028850|T047|AB|378.9|ICD9CM|Eye movemnt disorder NOS|Eye movemnt disorder NOS
C0028850|T047|PT|378.9|ICD9CM|Unspecified disorder of eye movements|Unspecified disorder of eye movements
C0497217|T047|HT|379|ICD9CM|Other disorders of eye|Other disorders of eye
C1971635|T047|HT|379.0|ICD9CM|Scleritis and episcleritis|Scleritis and episcleritis
C0036416|T047|AB|379.00|ICD9CM|Scleritis NOS|Scleritis NOS
C0036416|T047|PT|379.00|ICD9CM|Scleritis, unspecified|Scleritis, unspecified
C0155351|T047|AB|379.01|ICD9CM|Episclerit periodic fugx|Episclerit periodic fugx
C0155351|T047|PT|379.01|ICD9CM|Episcleritis periodica fugax|Episcleritis periodica fugax
C0155352|T047|AB|379.02|ICD9CM|Nodular episcleritis|Nodular episcleritis
C0155352|T047|PT|379.02|ICD9CM|Nodular episcleritis|Nodular episcleritis
C0155353|T047|AB|379.03|ICD9CM|Anterior scleritis|Anterior scleritis
C0155353|T047|PT|379.03|ICD9CM|Anterior scleritis|Anterior scleritis
C0155354|T047|AB|379.04|ICD9CM|Scleromalacia perforans|Scleromalacia perforans
C0155354|T047|PT|379.04|ICD9CM|Scleromalacia perforans|Scleromalacia perforans
C0155355|T047|AB|379.05|ICD9CM|Scleritis w cornea invol|Scleritis w cornea invol
C0155355|T047|PT|379.05|ICD9CM|Scleritis with corneal involvement|Scleritis with corneal involvement
C0155356|T047|AB|379.06|ICD9CM|Brawny scleritis|Brawny scleritis
C0155356|T047|PT|379.06|ICD9CM|Brawny scleritis|Brawny scleritis
C0155357|T047|AB|379.07|ICD9CM|Posterior scleritis|Posterior scleritis
C0155357|T047|PT|379.07|ICD9CM|Posterior scleritis|Posterior scleritis
C0029734|T047|PT|379.09|ICD9CM|Other scleritis and episcleritis|Other scleritis and episcleritis
C0029734|T047|AB|379.09|ICD9CM|Scleritis NEC|Scleritis NEC
C0155358|T047|HT|379.1|ICD9CM|Other disorders of sclera|Other disorders of sclera
C0155359|T047|AB|379.11|ICD9CM|Scleral ectasia|Scleral ectasia
C0155359|T047|PT|379.11|ICD9CM|Scleral ectasia|Scleral ectasia
C0155360|T047|AB|379.12|ICD9CM|Staphyloma posticum|Staphyloma posticum
C0155360|T047|PT|379.12|ICD9CM|Staphyloma posticum|Staphyloma posticum
C0155361|T047|AB|379.13|ICD9CM|Equatorial staphyloma|Equatorial staphyloma
C0155361|T047|PT|379.13|ICD9CM|Equatorial staphyloma|Equatorial staphyloma
C0155362|T047|PT|379.14|ICD9CM|Anterior staphyloma, localized|Anterior staphyloma, localized
C0155362|T047|AB|379.14|ICD9CM|Local anterior staphylma|Local anterior staphylma
C0155363|T047|AB|379.15|ICD9CM|Ring staphyloma|Ring staphyloma
C0155363|T047|PT|379.15|ICD9CM|Ring staphyloma|Ring staphyloma
C0155364|T047|PT|379.16|ICD9CM|Other degenerative disorders of sclera|Other degenerative disorders of sclera
C0155364|T047|AB|379.16|ICD9CM|Scleral degen dis NEC|Scleral degen dis NEC
C0155358|T047|AB|379.19|ICD9CM|Disorder of sclera NEC|Disorder of sclera NEC
C0155358|T047|PT|379.19|ICD9CM|Other disorders of sclera|Other disorders of sclera
C0155365|T047|HT|379.2|ICD9CM|Disorders of vitreous body|Disorders of vitreous body
C0155366|T047|AB|379.21|ICD9CM|Vitreous degeneration|Vitreous degeneration
C0155366|T047|PT|379.21|ICD9CM|Vitreous degeneration|Vitreous degeneration
C0155367|T047|AB|379.22|ICD9CM|Crystal deposit vitreous|Crystal deposit vitreous
C0155367|T047|PT|379.22|ICD9CM|Crystalline deposits in vitreous|Crystalline deposits in vitreous
C0042909|T046|AB|379.23|ICD9CM|Vitreous hemorrhage|Vitreous hemorrhage
C0042909|T046|PT|379.23|ICD9CM|Vitreous hemorrhage|Vitreous hemorrhage
C0029872|T047|PT|379.24|ICD9CM|Other vitreous opacities|Other vitreous opacities
C0029872|T047|AB|379.24|ICD9CM|Vitreous opacities NEC|Vitreous opacities NEC
C0155368|T047|AB|379.25|ICD9CM|Vitreous membranes|Vitreous membranes
C0155368|T047|PT|379.25|ICD9CM|Vitreous membranes and strands|Vitreous membranes and strands
C0155369|T190|AB|379.26|ICD9CM|Vitreous prolapse|Vitreous prolapse
C0155369|T190|PT|379.26|ICD9CM|Vitreous prolapse|Vitreous prolapse
C2748203|T190|PT|379.27|ICD9CM|Vitreomacular adhesion|Vitreomacular adhesion
C2748203|T190|AB|379.27|ICD9CM|Vitreomacular adhesion|Vitreomacular adhesion
C0155370|T047|PT|379.29|ICD9CM|Other disorders of vitreous|Other disorders of vitreous
C0155370|T047|AB|379.29|ICD9CM|Vitreous disorders NEC|Vitreous disorders NEC
C0155371|T047|HT|379.3|ICD9CM|Aphakia and other disorders of lens|Aphakia and other disorders of lens
C0003534|T190|AB|379.31|ICD9CM|Aphakia|Aphakia
C0003534|T190|PT|379.31|ICD9CM|Aphakia|Aphakia
C0023316|T047|AB|379.32|ICD9CM|Subluxation of lens|Subluxation of lens
C0023316|T047|PT|379.32|ICD9CM|Subluxation of lens|Subluxation of lens
C0155372|T047|AB|379.33|ICD9CM|Ant dislocation of lens|Ant dislocation of lens
C0155372|T047|PT|379.33|ICD9CM|Anterior dislocation of lens|Anterior dislocation of lens
C0155373|T047|AB|379.34|ICD9CM|Post dislocation of lens|Post dislocation of lens
C0155373|T047|PT|379.34|ICD9CM|Posterior dislocation of lens|Posterior dislocation of lens
C0029590|T047|AB|379.39|ICD9CM|Disorders of lens NEC|Disorders of lens NEC
C0029590|T047|PT|379.39|ICD9CM|Other disorders of lens|Other disorders of lens
C0917967|T033|HT|379.4|ICD9CM|Anomalies of pupillary function|Anomalies of pupillary function
C0917967|T033|AB|379.40|ICD9CM|Abn pupil function NOS|Abn pupil function NOS
C0917967|T033|PT|379.40|ICD9CM|Abnormal pupillary function, unspecified|Abnormal pupillary function, unspecified
C0003079|T033|AB|379.41|ICD9CM|Anisocoria|Anisocoria
C0003079|T033|PT|379.41|ICD9CM|Anisocoria|Anisocoria
C0026205|T047|PT|379.42|ICD9CM|Miosis (persistent), not due to miotics|Miosis (persistent), not due to miotics
C0026205|T047|AB|379.42|ICD9CM|Miosis not d/t miotics|Miosis not d/t miotics
C0026962|T046|PT|379.43|ICD9CM|Mydriasis (persistent), not due to mydriatics|Mydriasis (persistent), not due to mydriatics
C0026962|T046|AB|379.43|ICD9CM|Mydriasis not d/t mydrtc|Mydriasis not d/t mydrtc
C0155375|T047|AB|379.45|ICD9CM|Argyll robertson pupil|Argyll robertson pupil
C0155375|T047|PT|379.45|ICD9CM|Argyll Robertson pupil, atypical|Argyll Robertson pupil, atypical
C0040416|T184|AB|379.46|ICD9CM|Tonic pupillary reaction|Tonic pupillary reaction
C0040416|T184|PT|379.46|ICD9CM|Tonic pupillary reaction|Tonic pupillary reaction
C0155376|T047|PT|379.49|ICD9CM|Other anomalies of pupillary function|Other anomalies of pupillary function
C0155376|T047|AB|379.49|ICD9CM|Pupil funct anomaly NEC|Pupil funct anomaly NEC
C0339666|T033|HT|379.5|ICD9CM|Nystagmus and other irregular eye movements|Nystagmus and other irregular eye movements
C0028738|T047|AB|379.50|ICD9CM|Nystagmus NOS|Nystagmus NOS
C0028738|T047|PT|379.50|ICD9CM|Nystagmus, unspecified|Nystagmus, unspecified
C0700501|T019|AB|379.51|ICD9CM|Congenital nystagmus|Congenital nystagmus
C0700501|T019|PT|379.51|ICD9CM|Congenital nystagmus|Congenital nystagmus
C0152225|T047|AB|379.52|ICD9CM|Latent nystagmus|Latent nystagmus
C0152225|T047|PT|379.52|ICD9CM|Latent nystagmus|Latent nystagmus
C0271384|T047|PT|379.53|ICD9CM|Visual deprivation nystagmus|Visual deprivation nystagmus
C0271384|T047|AB|379.53|ICD9CM|Visual deprivatn nystagm|Visual deprivatn nystagm
C0155379|T047|AB|379.54|ICD9CM|Nystagms w vestibulr dis|Nystagms w vestibulr dis
C0155379|T047|PT|379.54|ICD9CM|Nystagmus associated with disorders of the vestibular system|Nystagmus associated with disorders of the vestibular system
C0155380|T047|AB|379.55|ICD9CM|Dissociated nystagmus|Dissociated nystagmus
C0155380|T047|PT|379.55|ICD9CM|Dissociated nystagmus|Dissociated nystagmus
C0029620|T047|AB|379.56|ICD9CM|Nystagmus NEC|Nystagmus NEC
C0029620|T047|PT|379.56|ICD9CM|Other forms of nystagmus|Other forms of nystagmus
C0595983|T033|PT|379.57|ICD9CM|Deficiencies of saccadic eye movements|Deficiencies of saccadic eye movements
C0595983|T033|AB|379.57|ICD9CM|Saccadic eye movmnt def|Saccadic eye movmnt def
C0155382|T184|PT|379.58|ICD9CM|Deficiencies of smooth pursuit movements|Deficiencies of smooth pursuit movements
C0155382|T184|AB|379.58|ICD9CM|Smooth pursuit mvmnt def|Smooth pursuit mvmnt def
C0155383|T047|AB|379.59|ICD9CM|Irregular eye mvmnts NEC|Irregular eye mvmnts NEC
C0155383|T047|PT|379.59|ICD9CM|Other irregularities of eye movements|Other irregularities of eye movements
C1719449|T046|HT|379.6|ICD9CM|Inflammation (infection) of postprocedural bleb|Inflammation (infection) of postprocedural bleb
C1719445|T047|AB|379.60|ICD9CM|Inflam postproc bleb NOS|Inflam postproc bleb NOS
C1719445|T047|PT|379.60|ICD9CM|Inflammation (infection) of postprocedural bleb, unspecified|Inflammation (infection) of postprocedural bleb, unspecified
C1719446|T047|AB|379.61|ICD9CM|Inflam postproc bleb, 1|Inflam postproc bleb, 1
C1719446|T047|PT|379.61|ICD9CM|Inflammation (infection) of postprocedural bleb, stage 1|Inflammation (infection) of postprocedural bleb, stage 1
C1719447|T047|AB|379.62|ICD9CM|Inflam postproc bleb, 2|Inflam postproc bleb, 2
C1719447|T047|PT|379.62|ICD9CM|Inflammation (infection) of postprocedural bleb, stage 2|Inflammation (infection) of postprocedural bleb, stage 2
C1719448|T047|AB|379.63|ICD9CM|Inflam postproc bleb, 3|Inflam postproc bleb, 3
C1719448|T047|PT|379.63|ICD9CM|Inflammation (infection) of postprocedural bleb, stage 3|Inflammation (infection) of postprocedural bleb, stage 3
C0155384|T047|AB|379.8|ICD9CM|Eye disorders NEC|Eye disorders NEC
C0155384|T047|PT|379.8|ICD9CM|Other specified disorders of eye and adnexa|Other specified disorders of eye and adnexa
C1314803|T047|HT|379.9|ICD9CM|Unspecified disorder of eye and adnexa|Unspecified disorder of eye and adnexa
C0015397|T047|PT|379.90|ICD9CM|Disorder of eye, unspecified|Disorder of eye, unspecified
C0015397|T047|AB|379.90|ICD9CM|Eye disorder NOS|Eye disorder NOS
C0030197|T184|AB|379.91|ICD9CM|Pain in or around eye|Pain in or around eye
C0030197|T184|PT|379.91|ICD9CM|Pain in or around eye|Pain in or around eye
C0155386|T047|AB|379.92|ICD9CM|Swelling or mass of eye|Swelling or mass of eye
C0155386|T047|PT|379.92|ICD9CM|Swelling or mass of eye|Swelling or mass of eye
C0034915|T184|PT|379.93|ICD9CM|Redness or discharge of eye|Redness or discharge of eye
C0034915|T184|AB|379.93|ICD9CM|Redness/discharge of eye|Redness/discharge of eye
C0155387|T047|AB|379.99|ICD9CM|Ill-defined eye dis NEC|Ill-defined eye dis NEC
C0155387|T047|PT|379.99|ICD9CM|Other ill-defined disorders of eye|Other ill-defined disorders of eye
C0155388|T047|HT|380|ICD9CM|Disorders of external ear|Disorders of external ear
C0178269|T047|HT|380-389.99|ICD9CM|DISEASES OF THE EAR AND MASTOID PROCESS|DISEASES OF THE EAR AND MASTOID PROCESS
C0155389|T047|HT|380.0|ICD9CM|Perichondritis and chondritis of pinna|Perichondritis and chondritis of pinna
C0155389|T047|PT|380.00|ICD9CM|Perichondritis of pinna, unspecified|Perichondritis of pinna, unspecified
C0155389|T047|AB|380.00|ICD9CM|Perichondritis pinna NOS|Perichondritis pinna NOS
C0155390|T047|AB|380.01|ICD9CM|Ac perichondritis pinna|Ac perichondritis pinna
C0155390|T047|PT|380.01|ICD9CM|Acute perichondritis of pinna|Acute perichondritis of pinna
C0155391|T047|AB|380.02|ICD9CM|Chr perichondritis pinna|Chr perichondritis pinna
C0155391|T047|PT|380.02|ICD9CM|Chronic perichondritis of pinna|Chronic perichondritis of pinna
C0741305|T046|AB|380.03|ICD9CM|Chondritis of pinna|Chondritis of pinna
C0741305|T046|PT|380.03|ICD9CM|Chondritis of pinna|Chondritis of pinna
C0021355|T047|HT|380.1|ICD9CM|Infective otitis externa|Infective otitis externa
C0021355|T047|AB|380.10|ICD9CM|Infec otitis externa NOS|Infec otitis externa NOS
C0021355|T047|PT|380.10|ICD9CM|Infective otitis externa, unspecified|Infective otitis externa, unspecified
C0155392|T047|AB|380.11|ICD9CM|Acute infection of pinna|Acute infection of pinna
C0155392|T047|PT|380.11|ICD9CM|Acute infection of pinna|Acute infection of pinna
C0155393|T047|AB|380.12|ICD9CM|Acute swimmers' ear|Acute swimmers' ear
C0155393|T047|PT|380.12|ICD9CM|Acute swimmers' ear|Acute swimmers' ear
C0155394|T047|AB|380.13|ICD9CM|Ac infect extern ear NEC|Ac infect extern ear NEC
C0155394|T047|PT|380.13|ICD9CM|Other acute infections of external ear|Other acute infections of external ear
C0155395|T047|AB|380.14|ICD9CM|Malignant otitis externa|Malignant otitis externa
C0155395|T047|PT|380.14|ICD9CM|Malignant otitis externa|Malignant otitis externa
C0155396|T047|AB|380.15|ICD9CM|Chr mycot otitis externa|Chr mycot otitis externa
C0155396|T047|PT|380.15|ICD9CM|Chronic mycotic otitis externa|Chronic mycotic otitis externa
C0155397|T047|AB|380.16|ICD9CM|Chr inf otit externa NEC|Chr inf otit externa NEC
C0155397|T047|PT|380.16|ICD9CM|Other chronic infective otitis externa|Other chronic infective otitis externa
C0029695|T047|HT|380.2|ICD9CM|Other otitis externa|Other otitis externa
C0155398|T047|AB|380.21|ICD9CM|Cholesteatoma extern ear|Cholesteatoma extern ear
C0155398|T047|PT|380.21|ICD9CM|Cholesteatoma of external ear|Cholesteatoma of external ear
C0155399|T047|AB|380.22|ICD9CM|Acute otitis externa NEC|Acute otitis externa NEC
C0155399|T047|PT|380.22|ICD9CM|Other acute otitis externa|Other acute otitis externa
C0155400|T047|AB|380.23|ICD9CM|Chr otitis externa NEC|Chr otitis externa NEC
C0155400|T047|PT|380.23|ICD9CM|Other chronic otitis externa|Other chronic otitis externa
C0494553|T047|HT|380.3|ICD9CM|Noninfectious disorders of pinna|Noninfectious disorders of pinna
C0155402|T047|AB|380.30|ICD9CM|Disorder of pinna NOS|Disorder of pinna NOS
C0155402|T047|PT|380.30|ICD9CM|Disorder of pinna, unspecified|Disorder of pinna, unspecified
C0271413|T046|AB|380.31|ICD9CM|Hematoma auricle/pinna|Hematoma auricle/pinna
C0271413|T046|PT|380.31|ICD9CM|Hematoma of auricle or pinna|Hematoma of auricle or pinna
C0001170|T020|AB|380.32|ICD9CM|Acq deform auricle/pinna|Acq deform auricle/pinna
C0001170|T020|PT|380.32|ICD9CM|Acquired deformities of auricle or pinna|Acquired deformities of auricle or pinna
C0155404|T047|AB|380.39|ICD9CM|Noninfect dis pinna NEC|Noninfect dis pinna NEC
C0155404|T047|PT|380.39|ICD9CM|Other noninfectious disorders of pinna|Other noninfectious disorders of pinna
C0021092|T033|AB|380.4|ICD9CM|Impacted cerumen|Impacted cerumen
C0021092|T033|PT|380.4|ICD9CM|Impacted cerumen|Impacted cerumen
C0155405|T047|HT|380.5|ICD9CM|Acquired stenosis of external ear canal|Acquired stenosis of external ear canal
C0155405|T047|AB|380.50|ICD9CM|Acq stenos ear canal NOS|Acq stenos ear canal NOS
C0155405|T047|PT|380.50|ICD9CM|Acquired stenosis of external ear canal, unspecified as to cause|Acquired stenosis of external ear canal, unspecified as to cause
C0395839|T020|PT|380.51|ICD9CM|Acquired stenosis of external ear canal secondary to trauma|Acquired stenosis of external ear canal secondary to trauma
C0395839|T020|AB|380.51|ICD9CM|Stenosis ear d/t trauma|Stenosis ear d/t trauma
C0395841|T020|PT|380.52|ICD9CM|Acquired stenosis of external ear canal secondary to surgery|Acquired stenosis of external ear canal secondary to surgery
C0395841|T020|AB|380.52|ICD9CM|Stenosis ear d/t surgery|Stenosis ear d/t surgery
C0395842|T020|PT|380.53|ICD9CM|Acquired stenosis of external ear canal secondary to inflammation|Acquired stenosis of external ear canal secondary to inflammation
C0395842|T020|AB|380.53|ICD9CM|Stenosis ear d/t inflam|Stenosis ear d/t inflam
C0155410|T047|HT|380.8|ICD9CM|Other disorders of external ear|Other disorders of external ear
C0155411|T047|AB|380.81|ICD9CM|Exostosis ext ear canal|Exostosis ext ear canal
C0155411|T047|PT|380.81|ICD9CM|Exostosis of external ear canal|Exostosis of external ear canal
C0155410|T047|AB|380.89|ICD9CM|Dis external ear NEC|Dis external ear NEC
C0155410|T047|PT|380.89|ICD9CM|Other disorders of external ear|Other disorders of external ear
C0155388|T047|AB|380.9|ICD9CM|Dis external ear NOS|Dis external ear NOS
C0155388|T047|PT|380.9|ICD9CM|Unspecified disorder of external ear|Unspecified disorder of external ear
C0155413|T047|HT|381|ICD9CM|Nonsuppurative otitis media and Eustachian tube disorders|Nonsuppurative otitis media and Eustachian tube disorders
C0271432|T047|HT|381.0|ICD9CM|Acute nonsuppurative otitis media|Acute nonsuppurative otitis media
C0271432|T047|AB|381.00|ICD9CM|Ac nonsup otitis med NOS|Ac nonsup otitis med NOS
C0271432|T047|PT|381.00|ICD9CM|Acute nonsuppurative otitis media, unspecified|Acute nonsuppurative otitis media, unspecified
C0155415|T047|AB|381.01|ICD9CM|Ac serous otitis media|Ac serous otitis media
C0155415|T047|PT|381.01|ICD9CM|Acute serous otitis media|Acute serous otitis media
C0395863|T047|AB|381.02|ICD9CM|Ac mucoid otitis media|Ac mucoid otitis media
C0395863|T047|PT|381.02|ICD9CM|Acute mucoid otitis media|Acute mucoid otitis media
C0395865|T047|AB|381.03|ICD9CM|Ac sanguin otitis media|Ac sanguin otitis media
C0395865|T047|PT|381.03|ICD9CM|Acute sanguinous otitis media|Acute sanguinous otitis media
C0155418|T047|AB|381.04|ICD9CM|Ac allergic serous OM|Ac allergic serous OM
C0155418|T047|PT|381.04|ICD9CM|Acute allergic serous otitis media|Acute allergic serous otitis media
C0155419|T047|AB|381.05|ICD9CM|Ac allergic mucoid OM|Ac allergic mucoid OM
C0155419|T047|PT|381.05|ICD9CM|Acute allergic mucoid otitis media|Acute allergic mucoid otitis media
C0155420|T047|AB|381.06|ICD9CM|Ac allerg sanguinous OM|Ac allerg sanguinous OM
C0155420|T047|PT|381.06|ICD9CM|Acute allergic sanguinous otitis media|Acute allergic sanguinous otitis media
C0155421|T047|HT|381.1|ICD9CM|Chronic serous otitis media|Chronic serous otitis media
C0155422|T047|AB|381.10|ICD9CM|Chr serous OM simp/NOS|Chr serous OM simp/NOS
C0155422|T047|PT|381.10|ICD9CM|Chronic serous otitis media, simple or unspecified|Chronic serous otitis media, simple or unspecified
C0155423|T047|AB|381.19|ICD9CM|Chr serous OM NEC|Chr serous OM NEC
C0155423|T047|PT|381.19|ICD9CM|Other chronic serous otitis media|Other chronic serous otitis media
C1455742|T047|HT|381.2|ICD9CM|Chronic mucoid otitis media|Chronic mucoid otitis media
C1455742|T047|AB|381.20|ICD9CM|Chr mucoid OM simp/NOS|Chr mucoid OM simp/NOS
C1455742|T047|PT|381.20|ICD9CM|Chronic mucoid otitis media, simple or unspecified|Chronic mucoid otitis media, simple or unspecified
C0155426|T047|AB|381.29|ICD9CM|Chr mucoid OM NEC|Chr mucoid OM NEC
C0155426|T047|PT|381.29|ICD9CM|Other chronic mucoid otitis media|Other chronic mucoid otitis media
C0155427|T047|AB|381.3|ICD9CM|Chr nonsup OM NOS/NEC|Chr nonsup OM NOS/NEC
C0155427|T047|PT|381.3|ICD9CM|Other and unspecified chronic nonsuppurative otitis media|Other and unspecified chronic nonsuppurative otitis media
C0271446|T047|AB|381.4|ICD9CM|Nonsupp otitis media NOS|Nonsupp otitis media NOS
C0271446|T047|PT|381.4|ICD9CM|Nonsuppurative otitis media, not specified as acute or chronic|Nonsuppurative otitis media, not specified as acute or chronic
C0155428|T047|HT|381.5|ICD9CM|Eustachian salpingitis|Eustachian salpingitis
C0155428|T047|AB|381.50|ICD9CM|Eustachian salping NOS|Eustachian salping NOS
C0155428|T047|PT|381.50|ICD9CM|Eustachian salpingitis, unspecified|Eustachian salpingitis, unspecified
C0155429|T047|AB|381.51|ICD9CM|Ac eustachian salping|Ac eustachian salping
C0155429|T047|PT|381.51|ICD9CM|Acute Eustachian salpingitis|Acute Eustachian salpingitis
C0155430|T047|AB|381.52|ICD9CM|Chr eustachian salping|Chr eustachian salping
C0155430|T047|PT|381.52|ICD9CM|Chronic Eustachian salpingitis|Chronic Eustachian salpingitis
C0149508|T033|HT|381.6|ICD9CM|Obstruction of Eustachian tube|Obstruction of Eustachian tube
C0149508|T033|AB|381.60|ICD9CM|Obstr eustach tube NOS|Obstr eustach tube NOS
C0149508|T033|PT|381.60|ICD9CM|Obstruction of Eustachian tube, unspecified|Obstruction of Eustachian tube, unspecified
C0155431|T047|AB|381.61|ICD9CM|Osseous eustachian obstr|Osseous eustachian obstr
C0155431|T047|PT|381.61|ICD9CM|Osseous obstruction of Eustachian tube|Osseous obstruction of Eustachian tube
C0271471|T047|PT|381.62|ICD9CM|Intrinsic cartilagenous obstruction of Eustachian tube|Intrinsic cartilagenous obstruction of Eustachian tube
C0271471|T047|AB|381.62|ICD9CM|Intrinsic eustach obstr|Intrinsic eustach obstr
C0155433|T047|PT|381.63|ICD9CM|Extrinsic cartilagenous obstruction of Eustachian tube|Extrinsic cartilagenous obstruction of Eustachian tube
C0155433|T047|AB|381.63|ICD9CM|Extrinsic eustach obstr|Extrinsic eustach obstr
C0155434|T047|AB|381.7|ICD9CM|Patulous eustachian tube|Patulous eustachian tube
C0155434|T047|PT|381.7|ICD9CM|Patulous Eustachian tube|Patulous Eustachian tube
C0155435|T047|HT|381.8|ICD9CM|Other disorders of Eustachian tube|Other disorders of Eustachian tube
C0271468|T047|AB|381.81|ICD9CM|Dysfunct eustachian tube|Dysfunct eustachian tube
C0271468|T047|PT|381.81|ICD9CM|Dysfunction of Eustachian tube|Dysfunction of Eustachian tube
C0155435|T047|AB|381.89|ICD9CM|Eustachian tube dis NEC|Eustachian tube dis NEC
C0155435|T047|PT|381.89|ICD9CM|Other disorders of Eustachian tube|Other disorders of Eustachian tube
C0271468|T047|AB|381.9|ICD9CM|Eustachian tube dis NOS|Eustachian tube dis NOS
C0271468|T047|PT|381.9|ICD9CM|Unspecified Eustachian tube disorder|Unspecified Eustachian tube disorder
C0029888|T047|HT|382|ICD9CM|Suppurative and unspecified otitis media|Suppurative and unspecified otitis media
C0271431|T047|HT|382.0|ICD9CM|Acute suppurative otitis media|Acute suppurative otitis media
C0395861|T047|AB|382.00|ICD9CM|Ac supp otitis media NOS|Ac supp otitis media NOS
C0395861|T047|PT|382.00|ICD9CM|Acute suppurative otitis media without spontaneous rupture of eardrum|Acute suppurative otitis media without spontaneous rupture of eardrum
C0395862|T047|AB|382.01|ICD9CM|Ac supp OM w drum rupt|Ac supp OM w drum rupt
C0395862|T047|PT|382.01|ICD9CM|Acute suppurative otitis media with spontaneous rupture of eardrum|Acute suppurative otitis media with spontaneous rupture of eardrum
C0155439|T047|AB|382.02|ICD9CM|Ac supp OM in oth dis|Ac supp OM in oth dis
C0155439|T047|PT|382.02|ICD9CM|Acute suppurative otitis media in diseases classified elsewhere|Acute suppurative otitis media in diseases classified elsewhere
C0155440|T047|AB|382.1|ICD9CM|Chr tubotympan suppur OM|Chr tubotympan suppur OM
C0155440|T047|PT|382.1|ICD9CM|Chronic tubotympanic suppurative otitis media|Chronic tubotympanic suppurative otitis media
C0155441|T047|AB|382.2|ICD9CM|Chr atticoantral sup OM|Chr atticoantral sup OM
C0155441|T047|PT|382.2|ICD9CM|Chronic atticoantral suppurative otitis media|Chronic atticoantral suppurative otitis media
C0271454|T047|AB|382.3|ICD9CM|Chr sup otitis media NOS|Chr sup otitis media NOS
C0271454|T047|PT|382.3|ICD9CM|Unspecified chronic suppurative otitis media|Unspecified chronic suppurative otitis media
C0029888|T047|AB|382.4|ICD9CM|Suppur otitis media NOS|Suppur otitis media NOS
C0029888|T047|PT|382.4|ICD9CM|Unspecified suppurative otitis media|Unspecified suppurative otitis media
C0029882|T047|AB|382.9|ICD9CM|Otitis media NOS|Otitis media NOS
C0029882|T047|PT|382.9|ICD9CM|Unspecified otitis media|Unspecified otitis media
C0155442|T047|HT|383|ICD9CM|Mastoiditis and related conditions|Mastoiditis and related conditions
C0701825|T047|HT|383.0|ICD9CM|Acute mastoiditis|Acute mastoiditis
C0795702|T047|AB|383.00|ICD9CM|Ac mastoiditis w/o compl|Ac mastoiditis w/o compl
C0795702|T047|PT|383.00|ICD9CM|Acute mastoiditis without complications|Acute mastoiditis without complications
C0155445|T047|AB|383.01|ICD9CM|Subperi mastoid abscess|Subperi mastoid abscess
C0155445|T047|PT|383.01|ICD9CM|Subperiosteal abscess of mastoid|Subperiosteal abscess of mastoid
C0155446|T047|AB|383.02|ICD9CM|Ac mastoiditis-compl NEC|Ac mastoiditis-compl NEC
C0155446|T047|PT|383.02|ICD9CM|Acute mastoiditis with other complications|Acute mastoiditis with other complications
C0155447|T047|AB|383.1|ICD9CM|Chronic mastoiditis|Chronic mastoiditis
C0155447|T047|PT|383.1|ICD9CM|Chronic mastoiditis|Chronic mastoiditis
C0155448|T047|HT|383.2|ICD9CM|Petrositis|Petrositis
C0155448|T047|AB|383.20|ICD9CM|Petrositis NOS|Petrositis NOS
C0155448|T047|PT|383.20|ICD9CM|Petrositis, unspecified|Petrositis, unspecified
C0155449|T047|AB|383.21|ICD9CM|Acute petrositis|Acute petrositis
C0155449|T047|PT|383.21|ICD9CM|Acute petrositis|Acute petrositis
C0155450|T047|AB|383.22|ICD9CM|Chronic petrositis|Chronic petrositis
C0155450|T047|PT|383.22|ICD9CM|Chronic petrositis|Chronic petrositis
C0155452|T046|HT|383.3|ICD9CM|Complications following mastoidectomy|Complications following mastoidectomy
C0155452|T046|AB|383.30|ICD9CM|Postmastoid compl NOS|Postmastoid compl NOS
C0155452|T046|PT|383.30|ICD9CM|Postmastoidectomy complication, unspecified|Postmastoidectomy complication, unspecified
C0155453|T047|PT|383.31|ICD9CM|Mucosal cyst of postmastoidectomy cavity|Mucosal cyst of postmastoidectomy cavity
C0155453|T047|AB|383.31|ICD9CM|Postmastoid mucosal cyst|Postmastoid mucosal cyst
C0155454|T047|AB|383.32|ICD9CM|Postmastoid cholesteatma|Postmastoid cholesteatma
C0155454|T047|PT|383.32|ICD9CM|Recurrent cholesteatoma of postmastoidectomy cavity|Recurrent cholesteatoma of postmastoidectomy cavity
C0155455|T046|PT|383.33|ICD9CM|Granulations of postmastoidectomy cavity|Granulations of postmastoidectomy cavity
C0155455|T046|AB|383.33|ICD9CM|Postmastoid granulations|Postmastoid granulations
C0155456|T047|HT|383.8|ICD9CM|Other disorders of mastoid|Other disorders of mastoid
C0395905|T020|AB|383.81|ICD9CM|Postauricular fistula|Postauricular fistula
C0395905|T020|PT|383.81|ICD9CM|Postauricular fistula|Postauricular fistula
C0155456|T047|AB|383.89|ICD9CM|Disorders of mastoid NEC|Disorders of mastoid NEC
C0155456|T047|PT|383.89|ICD9CM|Other disorders of mastoid|Other disorders of mastoid
C0024904|T047|AB|383.9|ICD9CM|Mastoiditis NOS|Mastoiditis NOS
C0024904|T047|PT|383.9|ICD9CM|Unspecified mastoiditis|Unspecified mastoiditis
C0155458|T047|HT|384|ICD9CM|Other disorders of tympanic membrane|Other disorders of tympanic membrane
C0155459|T047|HT|384.0|ICD9CM|Acute myringitis without mention of otitis media|Acute myringitis without mention of otitis media
C0155460|T047|AB|384.00|ICD9CM|Acute myringitis NOS|Acute myringitis NOS
C0155460|T047|PT|384.00|ICD9CM|Acute myringitis, unspecified|Acute myringitis, unspecified
C0155461|T047|AB|384.01|ICD9CM|Bullous myringitis|Bullous myringitis
C0155461|T047|PT|384.01|ICD9CM|Bullous myringitis|Bullous myringitis
C0155462|T047|AB|384.09|ICD9CM|Acute myringitis NEC|Acute myringitis NEC
C0155462|T047|PT|384.09|ICD9CM|Other acute myringitis without mention of otitis media|Other acute myringitis without mention of otitis media
C0395849|T047|AB|384.1|ICD9CM|Chronic myringitis|Chronic myringitis
C0395849|T047|PT|384.1|ICD9CM|Chronic myringitis without mention of otitis media|Chronic myringitis without mention of otitis media
C0206504|T037|HT|384.2|ICD9CM|Perforation of tympanic membrane|Perforation of tympanic membrane
C0206504|T037|AB|384.20|ICD9CM|Perforat tympan memb NOS|Perforat tympan memb NOS
C0206504|T037|PT|384.20|ICD9CM|Perforation of tympanic membrane, unspecified|Perforation of tympanic membrane, unspecified
C0155464|T020|AB|384.21|ICD9CM|Cent perf tympanic memb|Cent perf tympanic memb
C0155464|T020|PT|384.21|ICD9CM|Central perforation of tympanic membrane|Central perforation of tympanic membrane
C0155465|T033|AB|384.22|ICD9CM|Attic perf tympanic memb|Attic perf tympanic memb
C0155465|T033|PT|384.22|ICD9CM|Attic perforation of tympanic membrane|Attic perforation of tympanic membrane
C0155466|T047|AB|384.23|ICD9CM|Marginal perf tymp NEC|Marginal perf tymp NEC
C0155466|T047|PT|384.23|ICD9CM|Other marginal perforation of tympanic membrane|Other marginal perforation of tympanic membrane
C0155467|T047|AB|384.24|ICD9CM|Mult perf tympanic memb|Mult perf tympanic memb
C0155467|T047|PT|384.24|ICD9CM|Multiple perforations of tympanic membrane|Multiple perforations of tympanic membrane
C0155468|T047|AB|384.25|ICD9CM|Total perf tympanic memb|Total perf tympanic memb
C0155468|T047|PT|384.25|ICD9CM|Total perforation of tympanic membrane|Total perforation of tympanic membrane
C0155469|T047|HT|384.8|ICD9CM|Other specified disorders of tympanic membrane|Other specified disorders of tympanic membrane
C0155470|T047|AB|384.81|ICD9CM|Atrophic flaccid tympan|Atrophic flaccid tympan
C0155470|T047|PT|384.81|ICD9CM|Atrophic flaccid tympanic membrane|Atrophic flaccid tympanic membrane
C0155471|T047|AB|384.82|ICD9CM|Atrophic nonflaccid tymp|Atrophic nonflaccid tymp
C0155471|T047|PT|384.82|ICD9CM|Atrophic nonflaccid tympanic membrane|Atrophic nonflaccid tympanic membrane
C0041825|T047|AB|384.9|ICD9CM|Dis tympanic memb NOS|Dis tympanic memb NOS
C0041825|T047|PT|384.9|ICD9CM|Unspecified disorder of tympanic membrane|Unspecified disorder of tympanic membrane
C0155472|T047|HT|385|ICD9CM|Other disorders of middle ear and mastoid|Other disorders of middle ear and mastoid
C0395887|T047|HT|385.0|ICD9CM|Tympanosclerosis|Tympanosclerosis
C0395887|T047|AB|385.00|ICD9CM|Tympanosclerosis NOS|Tympanosclerosis NOS
C0395887|T047|PT|385.00|ICD9CM|Tympanosclerosis, unspecified as to involvement|Tympanosclerosis, unspecified as to involvement
C0395888|T047|AB|385.01|ICD9CM|Tympanoscl-tympanic memb|Tympanoscl-tympanic memb
C0395888|T047|PT|385.01|ICD9CM|Tympanosclerosis involving tympanic membrane only|Tympanosclerosis involving tympanic membrane only
C0395889|T047|PT|385.02|ICD9CM|Tympanosclerosis involving tympanic membrane and ear ossicles|Tympanosclerosis involving tympanic membrane and ear ossicles
C0395889|T047|AB|385.02|ICD9CM|Tympnoscler-tymp/ossicle|Tympnoscler-tymp/ossicle
C0395890|T047|AB|385.03|ICD9CM|Tympanoscler-all parts|Tympanoscler-all parts
C0395890|T047|PT|385.03|ICD9CM|Tympanosclerosis involving tympanic membrane, ear ossicles, and middle ear|Tympanosclerosis involving tympanic membrane, ear ossicles, and middle ear
C0155477|T047|PT|385.09|ICD9CM|Tympanosclerosis involving other combination of structures|Tympanosclerosis involving other combination of structures
C0155477|T047|AB|385.09|ICD9CM|Tympnsclr-oth site comb|Tympnsclr-oth site comb
C0155478|T047|HT|385.1|ICD9CM|Adhesive middle ear disease|Adhesive middle ear disease
C0155478|T047|AB|385.10|ICD9CM|Adhesive mid ear dis NOS|Adhesive mid ear dis NOS
C0155478|T047|PT|385.10|ICD9CM|Adhesive middle ear disease, unspecified as to involvement|Adhesive middle ear disease, unspecified as to involvement
C0155480|T047|AB|385.11|ICD9CM|Adhesion tympanum-incus|Adhesion tympanum-incus
C0155480|T047|PT|385.11|ICD9CM|Adhesions of drum head to incus|Adhesions of drum head to incus
C0155481|T047|AB|385.12|ICD9CM|Adhesion tympanum-stapes|Adhesion tympanum-stapes
C0155481|T047|PT|385.12|ICD9CM|Adhesions of drum head to stapes|Adhesions of drum head to stapes
C0155482|T047|AB|385.13|ICD9CM|Adhesion tymp-promontor|Adhesion tymp-promontor
C0155482|T047|PT|385.13|ICD9CM|Adhesions of drum head to promontorium|Adhesions of drum head to promontorium
C0155483|T047|AB|385.19|ICD9CM|Adhesive mid ear dis NEC|Adhesive mid ear dis NEC
C0155483|T047|PT|385.19|ICD9CM|Other middle ear adhesions and combinations|Other middle ear adhesions and combinations
C0155484|T020|HT|385.2|ICD9CM|Other acquired abnormality of ear ossicles|Other acquired abnormality of ear ossicles
C0584793|T033|AB|385.21|ICD9CM|Ankylosis malleus|Ankylosis malleus
C0584793|T033|PT|385.21|ICD9CM|Impaired mobility of malleus|Impaired mobility of malleus
C0155486|T047|AB|385.22|ICD9CM|Ankylosis ear ossicl NEC|Ankylosis ear ossicl NEC
C0155486|T047|PT|385.22|ICD9CM|Impaired mobility of other ear ossicles|Impaired mobility of other ear ossicles
C0155487|T020|PT|385.23|ICD9CM|Discontinuity or dislocation of ear ossicles|Discontinuity or dislocation of ear ossicles
C0155487|T020|AB|385.23|ICD9CM|Dislocation ear ossicle|Dislocation ear ossicle
C0155488|T047|AB|385.24|ICD9CM|Partial loss ear ossicle|Partial loss ear ossicle
C0155488|T047|PT|385.24|ICD9CM|Partial loss or necrosis of ear ossicles|Partial loss or necrosis of ear ossicles
C0008374|T047|HT|385.3|ICD9CM|Cholesteatoma of middle ear and mastoid|Cholesteatoma of middle ear and mastoid
C0008373|T047|AB|385.30|ICD9CM|Cholesteatoma NOS|Cholesteatoma NOS
C0008373|T047|PT|385.30|ICD9CM|Cholesteatoma, unspecified|Cholesteatoma, unspecified
C0155489|T047|AB|385.31|ICD9CM|Cholesteatoma of attic|Cholesteatoma of attic
C0155489|T047|PT|385.31|ICD9CM|Cholesteatoma of attic|Cholesteatoma of attic
C0155490|T047|AB|385.32|ICD9CM|Cholesteatoma middle ear|Cholesteatoma middle ear
C0155490|T047|PT|385.32|ICD9CM|Cholesteatoma of middle ear|Cholesteatoma of middle ear
C0008374|T047|PT|385.33|ICD9CM|Cholesteatoma of middle ear and mastoid|Cholesteatoma of middle ear and mastoid
C0008374|T047|AB|385.33|ICD9CM|Cholestma mid ear/mstoid|Cholestma mid ear/mstoid
C0155491|T047|AB|385.35|ICD9CM|Diffuse cholesteatosis|Diffuse cholesteatosis
C0155491|T047|PT|385.35|ICD9CM|Diffuse cholesteatosis of middle ear and mastoid|Diffuse cholesteatosis of middle ear and mastoid
C0155472|T047|HT|385.8|ICD9CM|Other disorders of middle ear and mastoid|Other disorders of middle ear and mastoid
C0155492|T047|AB|385.82|ICD9CM|Cholesterin granuloma|Cholesterin granuloma
C0155492|T047|PT|385.82|ICD9CM|Cholesterin granuloma of middle ear and mastoid|Cholesterin granuloma of middle ear and mastoid
C0155493|T047|AB|385.83|ICD9CM|Foreign body middle ear|Foreign body middle ear
C0155493|T047|PT|385.83|ICD9CM|Retained foreign body of middle ear|Retained foreign body of middle ear
C0155472|T047|AB|385.89|ICD9CM|Dis mid ear/mastoid NEC|Dis mid ear/mastoid NEC
C0155472|T047|PT|385.89|ICD9CM|Other disorders of middle ear and mastoid|Other disorders of middle ear and mastoid
C0155494|T047|AB|385.9|ICD9CM|Dis mid ear/mastoid NOS|Dis mid ear/mastoid NOS
C0155494|T047|PT|385.9|ICD9CM|Unspecified disorder of middle ear and mastoid|Unspecified disorder of middle ear and mastoid
C0155523|T047|HT|386|ICD9CM|Vertiginous syndromes and other disorders of vestibular system|Vertiginous syndromes and other disorders of vestibular system
C0025281|T047|HT|386.0|ICD9CM|Meniere's disease|Meniere's disease
C0025281|T047|AB|386.00|ICD9CM|Meniere's disease NOS|Meniere's disease NOS
C0025281|T047|PT|386.00|ICD9CM|Ménière's disease, unspecified|Ménière's disease, unspecified
C0155496|T047|PT|386.01|ICD9CM|Active Ménière's disease, cochleovestibular|Active Ménière's disease, cochleovestibular
C0155496|T047|AB|386.01|ICD9CM|Actv Meniere,cochlvestib|Actv Meniere,cochlvestib
C0155497|T047|AB|386.02|ICD9CM|Active Meniere, cochlear|Active Meniere, cochlear
C0155497|T047|PT|386.02|ICD9CM|Active Ménière's disease, cochlear|Active Ménière's disease, cochlear
C0155498|T047|PT|386.03|ICD9CM|Active Ménière's disease, vestibular|Active Ménière's disease, vestibular
C0155498|T047|AB|386.03|ICD9CM|Actv Meniere, vestibular|Actv Meniere, vestibular
C0155499|T047|AB|386.04|ICD9CM|Inactive Meniere's dis|Inactive Meniere's dis
C0155499|T047|PT|386.04|ICD9CM|Inactive Ménière's disease|Inactive Ménière's disease
C0029706|T047|HT|386.1|ICD9CM|Other and unspecified peripheral vertigo|Other and unspecified peripheral vertigo
C0155501|T047|AB|386.10|ICD9CM|Peripheral vertigo NOS|Peripheral vertigo NOS
C0155501|T047|PT|386.10|ICD9CM|Peripheral vertigo, unspecified|Peripheral vertigo, unspecified
C0155502|T047|PT|386.11|ICD9CM|Benign paroxysmal positional vertigo|Benign paroxysmal positional vertigo
C0155502|T047|AB|386.11|ICD9CM|Benign parxysmal vertigo|Benign parxysmal vertigo
C0751908|T047|AB|386.12|ICD9CM|Vestibular neuronitis|Vestibular neuronitis
C0751908|T047|PT|386.12|ICD9CM|Vestibular neuronitis|Vestibular neuronitis
C0029706|T047|PT|386.19|ICD9CM|Other peripheral vertigo|Other peripheral vertigo
C0029706|T047|AB|386.19|ICD9CM|Peripheral vertigo NEC|Peripheral vertigo NEC
C0155503|T047|AB|386.2|ICD9CM|Central origin vertigo|Central origin vertigo
C0155503|T047|PT|386.2|ICD9CM|Vertigo of central origin|Vertigo of central origin
C0022893|T047|HT|386.3|ICD9CM|Labyrinthitis|Labyrinthitis
C0022893|T047|AB|386.30|ICD9CM|Labyrinthitis NOS|Labyrinthitis NOS
C0022893|T047|PT|386.30|ICD9CM|Labyrinthitis, unspecified|Labyrinthitis, unspecified
C0155504|T047|AB|386.31|ICD9CM|Serous labyrinthitis|Serous labyrinthitis
C0155504|T047|PT|386.31|ICD9CM|Serous labyrinthitis|Serous labyrinthitis
C0155505|T047|AB|386.32|ICD9CM|Circumscri labyrinthitis|Circumscri labyrinthitis
C0155505|T047|PT|386.32|ICD9CM|Circumscribed labyrinthitis|Circumscribed labyrinthitis
C0155506|T047|AB|386.33|ICD9CM|Suppurativ labyrinthitis|Suppurativ labyrinthitis
C0155506|T047|PT|386.33|ICD9CM|Suppurative labyrinthitis|Suppurative labyrinthitis
C0155507|T047|AB|386.34|ICD9CM|Toxic labyrinthitis|Toxic labyrinthitis
C0155507|T047|PT|386.34|ICD9CM|Toxic labyrinthitis|Toxic labyrinthitis
C0155508|T047|AB|386.35|ICD9CM|Viral labyrinthitis|Viral labyrinthitis
C0155508|T047|PT|386.35|ICD9CM|Viral labyrinthitis|Viral labyrinthitis
C0155509|T190|HT|386.4|ICD9CM|Labyrinthine fistula|Labyrinthine fistula
C0155509|T190|AB|386.40|ICD9CM|Labyrinthine fistula NOS|Labyrinthine fistula NOS
C0155509|T190|PT|386.40|ICD9CM|Labyrinthine fistula, unspecified|Labyrinthine fistula, unspecified
C0339781|T020|AB|386.41|ICD9CM|Round window fistula|Round window fistula
C0339781|T020|PT|386.41|ICD9CM|Round window fistula|Round window fistula
C0339782|T020|AB|386.42|ICD9CM|Oval window fistula|Oval window fistula
C0339782|T020|PT|386.42|ICD9CM|Oval window fistula|Oval window fistula
C0155512|T190|AB|386.43|ICD9CM|Semicircul canal fistula|Semicircul canal fistula
C0155512|T190|PT|386.43|ICD9CM|Semicircular canal fistula|Semicircular canal fistula
C0155513|T190|AB|386.48|ICD9CM|Labyrinth fistula comb|Labyrinth fistula comb
C0155513|T190|PT|386.48|ICD9CM|Labyrinthine fistula of combined sites|Labyrinthine fistula of combined sites
C0155514|T047|HT|386.5|ICD9CM|Labyrinthine dysfunction|Labyrinthine dysfunction
C0155514|T047|AB|386.50|ICD9CM|Labyrinthine dysfunc NOS|Labyrinthine dysfunc NOS
C0155514|T047|PT|386.50|ICD9CM|Labyrinthine dysfunction, unspecified|Labyrinthine dysfunction, unspecified
C0155515|T047|PT|386.51|ICD9CM|Hyperactive labyrinth, unilateral|Hyperactive labyrinth, unilateral
C0155515|T047|AB|386.51|ICD9CM|Hypract labyrinth unilat|Hypract labyrinth unilat
C0155516|T047|AB|386.52|ICD9CM|Hyperact labyrinth bilat|Hyperact labyrinth bilat
C0155516|T047|PT|386.52|ICD9CM|Hyperactive labyrinth, bilateral|Hyperactive labyrinth, bilateral
C0155517|T047|AB|386.53|ICD9CM|Hypoact labyrinth unilat|Hypoact labyrinth unilat
C0155517|T047|PT|386.53|ICD9CM|Hypoactive labyrinth, unilateral|Hypoactive labyrinth, unilateral
C0155518|T047|AB|386.54|ICD9CM|Hypoact labyrinth bilat|Hypoact labyrinth bilat
C0155518|T047|PT|386.54|ICD9CM|Hypoactive labyrinth, bilateral|Hypoactive labyrinth, bilateral
C0155519|T047|AB|386.55|ICD9CM|Loss labyrn react unilat|Loss labyrn react unilat
C0155519|T047|PT|386.55|ICD9CM|Loss of labyrinthine reactivity, unilateral|Loss of labyrinthine reactivity, unilateral
C0155520|T047|AB|386.56|ICD9CM|Loss labyrin react bilat|Loss labyrin react bilat
C0155520|T047|PT|386.56|ICD9CM|Loss of labyrinthine reactivity, bilateral|Loss of labyrinthine reactivity, bilateral
C0155521|T047|AB|386.58|ICD9CM|Labyrinthine dysfunc NEC|Labyrinthine dysfunc NEC
C0155521|T047|PT|386.58|ICD9CM|Other forms and combinations of labyrinthine dysfunction|Other forms and combinations of labyrinthine dysfunction
C0155522|T047|AB|386.8|ICD9CM|Disorders labyrinth NEC|Disorders labyrinth NEC
C0155522|T047|PT|386.8|ICD9CM|Other disorders of labyrinth|Other disorders of labyrinth
C0155523|T047|PT|386.9|ICD9CM|Unspecified vertiginous syndromes and labyrinthine disorders|Unspecified vertiginous syndromes and labyrinthine disorders
C0155523|T047|AB|386.9|ICD9CM|Vertiginous synd NOS|Vertiginous synd NOS
C0029899|T047|HT|387|ICD9CM|Otosclerosis|Otosclerosis
C0155524|T047|AB|387.0|ICD9CM|Otoscler-oval wnd nonobl|Otoscler-oval wnd nonobl
C0155524|T047|PT|387.0|ICD9CM|Otosclerosis involving oval window, nonobliterative|Otosclerosis involving oval window, nonobliterative
C0155525|T047|AB|387.1|ICD9CM|Otoscler-oval wndw oblit|Otoscler-oval wndw oblit
C0155525|T047|PT|387.1|ICD9CM|Otosclerosis involving oval window, obliterative|Otosclerosis involving oval window, obliterative
C0155526|T020|AB|387.2|ICD9CM|Cochlear otosclerosis|Cochlear otosclerosis
C0155526|T020|PT|387.2|ICD9CM|Cochlear otosclerosis|Cochlear otosclerosis
C0029696|T047|PT|387.8|ICD9CM|Other otosclerosis|Other otosclerosis
C0029696|T047|AB|387.8|ICD9CM|Otosclerosis NEC|Otosclerosis NEC
C0029899|T047|AB|387.9|ICD9CM|Otosclerosis NOS|Otosclerosis NOS
C0029899|T047|PT|387.9|ICD9CM|Otosclerosis, unspecified|Otosclerosis, unspecified
C0155527|T047|HT|388|ICD9CM|Other disorders of ear|Other disorders of ear
C0155528|T047|HT|388.0|ICD9CM|Degenerative and vascular disorders of ear|Degenerative and vascular disorders of ear
C0155528|T047|AB|388.00|ICD9CM|Degen/vascul dis ear NOS|Degen/vascul dis ear NOS
C0155528|T047|PT|388.00|ICD9CM|Degenerative and vascular disorders, unspecified|Degenerative and vascular disorders, unspecified
C0033074|T046|AB|388.01|ICD9CM|Presbyacusis|Presbyacusis
C0033074|T046|PT|388.01|ICD9CM|Presbyacusis|Presbyacusis
C0155530|T046|AB|388.02|ICD9CM|Trans ischemic deafness|Trans ischemic deafness
C0155530|T046|PT|388.02|ICD9CM|Transient ischemic deafness|Transient ischemic deafness
C0155531|T037|HT|388.1|ICD9CM|Noise effects on inner ear|Noise effects on inner ear
C0155531|T037|AB|388.10|ICD9CM|Noise effect-ear/NOS|Noise effect-ear/NOS
C0155531|T037|PT|388.10|ICD9CM|Noise effects on inner ear, unspecified|Noise effects on inner ear, unspecified
C0155532|T037|AB|388.11|ICD9CM|Acoustic trauma|Acoustic trauma
C0155532|T037|PT|388.11|ICD9CM|Acoustic trauma (explosive) to ear|Acoustic trauma (explosive) to ear
C0018781|T037|AB|388.12|ICD9CM|Hearing loss d/t noise|Hearing loss d/t noise
C0018781|T037|PT|388.12|ICD9CM|Noise-induced hearing loss|Noise-induced hearing loss
C0011057|T033|AB|388.2|ICD9CM|Sudden hearing loss NOS|Sudden hearing loss NOS
C0011057|T033|PT|388.2|ICD9CM|Sudden hearing loss, unspecified|Sudden hearing loss, unspecified
C0040264|T047|HT|388.3|ICD9CM|Tinnitus|Tinnitus
C0040264|T047|AB|388.30|ICD9CM|Tinnitus NOS|Tinnitus NOS
C0040264|T047|PT|388.30|ICD9CM|Tinnitus, unspecified|Tinnitus, unspecified
C0155533|T184|AB|388.31|ICD9CM|Subjective tinnitus|Subjective tinnitus
C0155533|T184|PT|388.31|ICD9CM|Subjective tinnitus|Subjective tinnitus
C0155534|T184|AB|388.32|ICD9CM|Objective tinnitus|Objective tinnitus
C0155534|T184|PT|388.32|ICD9CM|Objective tinnitus|Objective tinnitus
C0155535|T033|HT|388.4|ICD9CM|Other abnormal auditory perception|Other abnormal auditory perception
C0375257|T046|AB|388.40|ICD9CM|Abn auditory percept NOS|Abn auditory percept NOS
C0375257|T046|PT|388.40|ICD9CM|Abnormal auditory perception, unspecified|Abnormal auditory perception, unspecified
C0152228|T184|AB|388.41|ICD9CM|Diplacusis|Diplacusis
C0152228|T184|PT|388.41|ICD9CM|Diplacusis|Diplacusis
C0034880|T184|AB|388.42|ICD9CM|Hyperacusis|Hyperacusis
C0034880|T184|PT|388.42|ICD9CM|Hyperacusis|Hyperacusis
C0155537|T047|AB|388.43|ICD9CM|Impairm auditory discrim|Impairm auditory discrim
C0155537|T047|PT|388.43|ICD9CM|Impairment of auditory discrimination|Impairment of auditory discrimination
C0271510|T047|AB|388.44|ICD9CM|Auditory recruitment|Auditory recruitment
C0271510|T047|PT|388.44|ICD9CM|Auditory recruitment|Auditory recruitment
C1955771|T047|AB|388.45|ICD9CM|Acq auditory process dis|Acq auditory process dis
C1955771|T047|PT|388.45|ICD9CM|Acquired auditory processing disorder|Acquired auditory processing disorder
C0001163|T047|AB|388.5|ICD9CM|Acoustic nerve disorders|Acoustic nerve disorders
C0001163|T047|PT|388.5|ICD9CM|Disorders of acoustic nerve|Disorders of acoustic nerve
C0155540|T033|HT|388.6|ICD9CM|Otorrhea|Otorrhea
C0155540|T033|AB|388.60|ICD9CM|Otorrhea NOS|Otorrhea NOS
C0155540|T033|PT|388.60|ICD9CM|Otorrhea, unspecified|Otorrhea, unspecified
C0007814|T047|AB|388.61|ICD9CM|Cerebrosp fluid otorrhea|Cerebrosp fluid otorrhea
C0007814|T047|PT|388.61|ICD9CM|Cerebrospinal fluid otorrhea|Cerebrospinal fluid otorrhea
C0155541|T047|PT|388.69|ICD9CM|Other otorrhea|Other otorrhea
C0155541|T047|AB|388.69|ICD9CM|Otorrhea NEC|Otorrhea NEC
C0013456|T184|HT|388.7|ICD9CM|Otalgia|Otalgia
C0013456|T184|AB|388.70|ICD9CM|Otalgia NOS|Otalgia NOS
C0013456|T184|PT|388.70|ICD9CM|Otalgia, unspecified|Otalgia, unspecified
C0155542|T184|AB|388.71|ICD9CM|Otogenic pain|Otogenic pain
C0155542|T184|PT|388.71|ICD9CM|Otogenic pain|Otogenic pain
C0271411|T184|PT|388.72|ICD9CM|Referred otogenic pain|Referred otogenic pain
C0271411|T184|AB|388.72|ICD9CM|Referred pain of ear|Referred pain of ear
C0155527|T047|AB|388.8|ICD9CM|Disorders of ear NEC|Disorders of ear NEC
C0155527|T047|PT|388.8|ICD9CM|Other disorders of ear|Other disorders of ear
C0013447|T047|AB|388.9|ICD9CM|Disorder of ear NOS|Disorder of ear NOS
C0013447|T047|PT|388.9|ICD9CM|Unspecified disorder of ear|Unspecified disorder of ear
C1384666|T047|HT|389|ICD9CM|Hearing loss|Hearing loss
C0018777|T047|HT|389.0|ICD9CM|Conductive hearing loss|Conductive hearing loss
C0018777|T047|AB|389.00|ICD9CM|Conduct hearing loss NOS|Conduct hearing loss NOS
C0018777|T047|PT|389.00|ICD9CM|Conductive hearing loss, unspecified|Conductive hearing loss, unspecified
C0155544|T047|AB|389.01|ICD9CM|Conduc hear loss ext ear|Conduc hear loss ext ear
C0155544|T047|PT|389.01|ICD9CM|Conductive hearing loss, external ear|Conductive hearing loss, external ear
C0155545|T047|AB|389.02|ICD9CM|Conduct hear loss tympan|Conduct hear loss tympan
C0155545|T047|PT|389.02|ICD9CM|Conductive hearing loss, tympanic membrane|Conductive hearing loss, tympanic membrane
C0155546|T047|AB|389.03|ICD9CM|Conduc hear loss mid ear|Conduc hear loss mid ear
C0155546|T047|PT|389.03|ICD9CM|Conductive hearing loss, middle ear|Conductive hearing loss, middle ear
C0155547|T047|AB|389.04|ICD9CM|Cond hear loss inner ear|Cond hear loss inner ear
C0155547|T047|PT|389.04|ICD9CM|Conductive hearing loss, inner ear|Conductive hearing loss, inner ear
C1955772|T047|AB|389.05|ICD9CM|Condctv hear loss,unilat|Condctv hear loss,unilat
C1955772|T047|PT|389.05|ICD9CM|Conductive hearing loss, unilateral|Conductive hearing loss, unilateral
C0452136|T047|AB|389.06|ICD9CM|Condctv hear loss, bilat|Condctv hear loss, bilat
C0452136|T047|PT|389.06|ICD9CM|Conductive hearing loss, bilateral|Conductive hearing loss, bilateral
C0155548|T047|AB|389.08|ICD9CM|Cond hear loss comb type|Cond hear loss comb type
C0155548|T047|PT|389.08|ICD9CM|Conductive hearing loss of combined types|Conductive hearing loss of combined types
C0018784|T047|HT|389.1|ICD9CM|Sensorineural hearing loss|Sensorineural hearing loss
C0018784|T047|PT|389.10|ICD9CM|Sensorineural hearing loss, unspecified|Sensorineural hearing loss, unspecified
C0018784|T047|AB|389.10|ICD9CM|Sensorneur hear loss NOS|Sensorneur hear loss NOS
C1719452|T047|PT|389.11|ICD9CM|Sensory hearing loss, bilateral|Sensory hearing loss, bilateral
C1719452|T047|AB|389.11|ICD9CM|Sensry hearng loss,bilat|Sensry hearng loss,bilat
C2315695|T047|PT|389.12|ICD9CM|Neural hearing loss, bilateral|Neural hearing loss, bilateral
C2315695|T047|AB|389.12|ICD9CM|Neural hearng loss,bilat|Neural hearng loss,bilat
C1955773|T047|AB|389.13|ICD9CM|Neural hear loss, unilat|Neural hear loss, unilat
C1955773|T047|PT|389.13|ICD9CM|Neural hearing loss, unilateral|Neural hearing loss, unilateral
C0018776|T047|AB|389.14|ICD9CM|Central hearing loss|Central hearing loss
C0018776|T047|PT|389.14|ICD9CM|Central hearing loss|Central hearing loss
C0744667|T033|PT|389.15|ICD9CM|Sensorineural hearing loss, unilateral|Sensorineural hearing loss, unilateral
C0744667|T033|AB|389.15|ICD9CM|Sensorneur hear loss uni|Sensorneur hear loss uni
C1719455|T047|AB|389.16|ICD9CM|Sensoneur hear loss asym|Sensoneur hear loss asym
C1719455|T047|PT|389.16|ICD9CM|Sensorineural hearing loss, asymmetrical|Sensorineural hearing loss, asymmetrical
C1955774|T047|AB|389.17|ICD9CM|Sensory hear loss,unilat|Sensory hear loss,unilat
C1955774|T047|PT|389.17|ICD9CM|Sensory hearing loss, unilateral|Sensory hearing loss, unilateral
C0452138|T047|AB|389.18|ICD9CM|Sensonrl hear loss,bilat|Sensonrl hear loss,bilat
C0452138|T047|PT|389.18|ICD9CM|Sensorineural hearing loss, bilateral|Sensorineural hearing loss, bilateral
C0155552|T047|HT|389.2|ICD9CM|Mixed conductive and sensorineural hearing loss|Mixed conductive and sensorineural hearing loss
C0155552|T047|AB|389.20|ICD9CM|Mixed hearing loss NOS|Mixed hearing loss NOS
C0155552|T047|PT|389.20|ICD9CM|Mixed hearing loss, unspecified|Mixed hearing loss, unspecified
C1955775|T047|PT|389.21|ICD9CM|Mixed hearing loss, unilateral|Mixed hearing loss, unilateral
C1955775|T047|AB|389.21|ICD9CM|Mixed hearing loss,unilt|Mixed hearing loss,unilt
C0452153|T047|PT|389.22|ICD9CM|Mixed hearing loss, bilateral|Mixed hearing loss, bilateral
C0452153|T047|AB|389.22|ICD9CM|Mixed hearing loss,bilat|Mixed hearing loss,bilat
C1955777|T047|AB|389.7|ICD9CM|Deaf, nonspeaking NEC|Deaf, nonspeaking NEC
C1955777|T047|PT|389.7|ICD9CM|Deaf, nonspeaking, not elsewhere classifiable|Deaf, nonspeaking, not elsewhere classifiable
C0477458|T047|AB|389.8|ICD9CM|Hearing loss NEC|Hearing loss NEC
C0477458|T047|PT|389.8|ICD9CM|Other specified forms of hearing loss|Other specified forms of hearing loss
C1384666|T047|AB|389.9|ICD9CM|Hearing loss NOS|Hearing loss NOS
C1384666|T047|PT|389.9|ICD9CM|Unspecified hearing loss|Unspecified hearing loss
C0264743|T047|AB|390|ICD9CM|Rheum fev w/o hrt involv|Rheum fev w/o hrt involv
C0264743|T047|PT|390|ICD9CM|Rheumatic fever without mention of heart involvement|Rheumatic fever without mention of heart involvement
C0035436|T047|HT|390-392.99|ICD9CM|ACUTE RHEUMATIC FEVER|ACUTE RHEUMATIC FEVER
C0728936|T047|HT|390-459.99|ICD9CM|DISEASES OF THE CIRCULATORY SYSTEM|DISEASES OF THE CIRCULATORY SYSTEM
C3536892|T047|HT|391|ICD9CM|Rheumatic fever with heart involvement|Rheumatic fever with heart involvement
C0155555|T047|AB|391.0|ICD9CM|Acute rheumatic pericard|Acute rheumatic pericard
C0155555|T047|PT|391.0|ICD9CM|Acute rheumatic pericarditis|Acute rheumatic pericarditis
C0155556|T047|AB|391.1|ICD9CM|Acute rheumatic endocard|Acute rheumatic endocard
C0155556|T047|PT|391.1|ICD9CM|Acute rheumatic endocarditis|Acute rheumatic endocarditis
C0155557|T047|AB|391.2|ICD9CM|Ac rheumatic myocarditis|Ac rheumatic myocarditis
C0155557|T047|PT|391.2|ICD9CM|Acute rheumatic myocarditis|Acute rheumatic myocarditis
C0155558|T047|AB|391.8|ICD9CM|Ac rheumat hrt dis NEC|Ac rheumat hrt dis NEC
C0155558|T047|PT|391.8|ICD9CM|Other acute rheumatic heart disease|Other acute rheumatic heart disease
C0035440|T047|AB|391.9|ICD9CM|Ac rheumat hrt dis NOS|Ac rheumat hrt dis NOS
C0035440|T047|PT|391.9|ICD9CM|Acute rheumatic heart disease, unspecified|Acute rheumatic heart disease, unspecified
C0152113|T047|HT|392|ICD9CM|Rheumatic chorea|Rheumatic chorea
C0155559|T047|AB|392.0|ICD9CM|Rheum chorea w hrt invol|Rheum chorea w hrt invol
C0155559|T047|PT|392.0|ICD9CM|Rheumatic chorea with heart involvement|Rheumatic chorea with heart involvement
C0489958|T047|AB|392.9|ICD9CM|Rheumatic chorea NOS|Rheumatic chorea NOS
C0489958|T047|PT|392.9|ICD9CM|Rheumatic chorea without mention of heart involvement|Rheumatic chorea without mention of heart involvement
C0155561|T047|AB|393|ICD9CM|Chr rheumatic pericard|Chr rheumatic pericard
C0155561|T047|PT|393|ICD9CM|Chronic rheumatic pericarditis|Chronic rheumatic pericarditis
C0175708|T047|HT|393-398.99|ICD9CM|CHRONIC RHEUMATIC HEART DISEASE|CHRONIC RHEUMATIC HEART DISEASE
C0264765|T047|HT|394|ICD9CM|Diseases of mitral valve|Diseases of mitral valve
C0264766|T047|AB|394.0|ICD9CM|Mitral stenosis|Mitral stenosis
C0264766|T047|PT|394.0|ICD9CM|Mitral stenosis|Mitral stenosis
C0155563|T047|AB|394.1|ICD9CM|Rheumatic mitral insuff|Rheumatic mitral insuff
C0155563|T047|PT|394.1|ICD9CM|Rheumatic mitral insufficiency|Rheumatic mitral insufficiency
C0264767|T047|AB|394.2|ICD9CM|Mitral stenosis w insuff|Mitral stenosis w insuff
C0264767|T047|PT|394.2|ICD9CM|Mitral stenosis with insufficiency|Mitral stenosis with insufficiency
C0348579|T047|AB|394.9|ICD9CM|Mitral valve dis NEC/NOS|Mitral valve dis NEC/NOS
C0348579|T047|PT|394.9|ICD9CM|Other and unspecified mitral valve diseases|Other and unspecified mitral valve diseases
C1260873|T047|HT|395|ICD9CM|Diseases of aortic valve|Diseases of aortic valve
C0155567|T047|AB|395.0|ICD9CM|Rheumat aortic stenosis|Rheumat aortic stenosis
C0155567|T047|PT|395.0|ICD9CM|Rheumatic aortic stenosis|Rheumatic aortic stenosis
C0155568|T047|AB|395.1|ICD9CM|Rheumatic aortic insuff|Rheumatic aortic insuff
C0155568|T047|PT|395.1|ICD9CM|Rheumatic aortic insufficiency|Rheumatic aortic insufficiency
C0155569|T047|AB|395.2|ICD9CM|Rheum aortic sten/insuff|Rheum aortic sten/insuff
C0155569|T047|PT|395.2|ICD9CM|Rheumatic aortic stenosis with insufficiency|Rheumatic aortic stenosis with insufficiency
C0155570|T047|PT|395.9|ICD9CM|Other and unspecified rheumatic aortic diseases|Other and unspecified rheumatic aortic diseases
C0155570|T047|AB|395.9|ICD9CM|Rheum aortic dis NEC/NOS|Rheum aortic dis NEC/NOS
C0375259|T047|HT|396|ICD9CM|Diseases of mitral and aortic valves|Diseases of mitral and aortic valves
C0155572|T047|PT|396.0|ICD9CM|Mitral valve stenosis and aortic valve stenosis|Mitral valve stenosis and aortic valve stenosis
C0155572|T047|AB|396.0|ICD9CM|Mitral/aortic stenosis|Mitral/aortic stenosis
C0264772|T047|AB|396.1|ICD9CM|Mitral stenos/aort insuf|Mitral stenos/aort insuf
C0264772|T047|PT|396.1|ICD9CM|Mitral valve stenosis and aortic valve insufficiency|Mitral valve stenosis and aortic valve insufficiency
C1306822|T047|AB|396.2|ICD9CM|Mitral insuf/aort stenos|Mitral insuf/aort stenos
C1306822|T047|PT|396.2|ICD9CM|Mitral valve insufficiency and aortic valve stenosis|Mitral valve insufficiency and aortic valve stenosis
C0264774|T047|PT|396.3|ICD9CM|Mitral valve insufficiency and aortic valve insufficiency|Mitral valve insufficiency and aortic valve insufficiency
C0264774|T047|AB|396.3|ICD9CM|Mitral/aortic val insuff|Mitral/aortic val insuff
C0155576|T047|AB|396.8|ICD9CM|Mitr/aortic mult involv|Mitr/aortic mult involv
C0155576|T047|PT|396.8|ICD9CM|Multiple involvement of mitral and aortic valves|Multiple involvement of mitral and aortic valves
C0375259|T047|PT|396.9|ICD9CM|Mitral and aortic valve diseases, unspecified|Mitral and aortic valve diseases, unspecified
C0375259|T047|AB|396.9|ICD9CM|Mitral/aortic v dis NOS|Mitral/aortic v dis NOS
C0155578|T047|HT|397|ICD9CM|Diseases of other endocardial structures|Diseases of other endocardial structures
C0264776|T047|PT|397.0|ICD9CM|Diseases of tricuspid valve|Diseases of tricuspid valve
C0264776|T047|AB|397.0|ICD9CM|Tricuspid valve disease|Tricuspid valve disease
C0155579|T047|AB|397.1|ICD9CM|Rheum pulmon valve dis|Rheum pulmon valve dis
C0155579|T047|PT|397.1|ICD9CM|Rheumatic diseases of pulmonary valve|Rheumatic diseases of pulmonary valve
C0264764|T047|AB|397.9|ICD9CM|Rheum endocarditis NOS|Rheum endocarditis NOS
C0264764|T047|PT|397.9|ICD9CM|Rheumatic diseases of endocardium, valve unspecified|Rheumatic diseases of endocardium, valve unspecified
C0029730|T047|HT|398|ICD9CM|Other rheumatic heart disease|Other rheumatic heart disease
C0489959|T020|AB|398.0|ICD9CM|Rheumatic myocarditis|Rheumatic myocarditis
C0489959|T020|PT|398.0|ICD9CM|Rheumatic myocarditis|Rheumatic myocarditis
C0029730|T047|HT|398.9|ICD9CM|Other and unspecified rheumatic heart diseases|Other and unspecified rheumatic heart diseases
C0035439|T047|AB|398.90|ICD9CM|Rheumatic heart dis NOS|Rheumatic heart dis NOS
C0035439|T047|PT|398.90|ICD9CM|Rheumatic heart disease, unspecified|Rheumatic heart disease, unspecified
C0155582|T047|AB|398.91|ICD9CM|Rheumatic heart failure|Rheumatic heart failure
C0155582|T047|PT|398.91|ICD9CM|Rheumatic heart failure (congestive)|Rheumatic heart failure (congestive)
C0029730|T047|PT|398.99|ICD9CM|Other rheumatic heart diseases|Other rheumatic heart diseases
C0029730|T047|AB|398.99|ICD9CM|Rheumatic heart dis NEC|Rheumatic heart dis NEC
C0085580|T047|HT|401|ICD9CM|Essential hypertension|Essential hypertension
C0020538|T047|HT|401-405.99|ICD9CM|HYPERTENSIVE DISEASE|HYPERTENSIVE DISEASE
C0024588|T047|PT|401.0|ICD9CM|Malignant essential hypertension|Malignant essential hypertension
C0024588|T047|AB|401.0|ICD9CM|Malignant hypertension|Malignant hypertension
C0155583|T047|PT|401.1|ICD9CM|Benign essential hypertension|Benign essential hypertension
C0155583|T047|AB|401.1|ICD9CM|Benign hypertension|Benign hypertension
C0085580|T047|AB|401.9|ICD9CM|Hypertension NOS|Hypertension NOS
C0085580|T047|PT|401.9|ICD9CM|Unspecified essential hypertension|Unspecified essential hypertension
C0152105|T047|HT|402|ICD9CM|Hypertensive heart disease|Hypertensive heart disease
C0155584|T047|HT|402.0|ICD9CM|Malignant hypertensive heart disease|Malignant hypertensive heart disease
C1135328|T047|AB|402.00|ICD9CM|Mal hyp ht dis w/o hf|Mal hyp ht dis w/o hf
C1135328|T047|PT|402.00|ICD9CM|Malignant hypertensive heart disease without heart failure|Malignant hypertensive heart disease without heart failure
C1135329|T047|AB|402.01|ICD9CM|Mal hypert hrt dis w hf|Mal hypert hrt dis w hf
C1135329|T047|PT|402.01|ICD9CM|Malignant hypertensive heart disease with heart failure|Malignant hypertensive heart disease with heart failure
C0155587|T047|HT|402.1|ICD9CM|Benign hypertensive heart disease|Benign hypertensive heart disease
C1135330|T047|AB|402.10|ICD9CM|Benign hyp ht dis w/o hf|Benign hyp ht dis w/o hf
C1135330|T047|PT|402.10|ICD9CM|Benign hypertensive heart disease without heart failure|Benign hypertensive heart disease without heart failure
C1135331|T047|AB|402.11|ICD9CM|Benign hyp ht dis w hf|Benign hyp ht dis w hf
C1135331|T047|PT|402.11|ICD9CM|Benign hypertensive heart disease with heart failure|Benign hypertensive heart disease with heart failure
C0152105|T047|HT|402.9|ICD9CM|Unspecified hypertensive heart disease|Unspecified hypertensive heart disease
C1135332|T047|AB|402.90|ICD9CM|Hyp hrt dis NOS w/o hf|Hyp hrt dis NOS w/o hf
C1135332|T047|PT|402.90|ICD9CM|Unspecified hypertensive heart disease without heart failure|Unspecified hypertensive heart disease without heart failure
C1135333|T047|AB|402.91|ICD9CM|Hyp ht dis NOS w ht fail|Hyp ht dis NOS w ht fail
C1135333|T047|PT|402.91|ICD9CM|Unspecified hypertensive heart disease with heart failure|Unspecified hypertensive heart disease with heart failure
C3695318|T047|HT|403|ICD9CM|Hypertensive chronic kidney disease|Hypertensive chronic kidney disease
C1719462|T047|HT|403.0|ICD9CM|Hypertensive chronic kidney disease, malignant|Hypertensive chronic kidney disease, malignant
C1719460|T047|AB|403.00|ICD9CM|Mal hy kid w cr kid I-IV|Mal hy kid w cr kid I-IV
C1719461|T047|AB|403.01|ICD9CM|Mal hyp kid w cr kid V|Mal hyp kid w cr kid V
C0155596|T047|HT|403.1|ICD9CM|Hypertensive renal disease, benign|Hypertensive renal disease, benign
C0155596|T047|AB|403.10|ICD9CM|Ben hy kid w cr kid I-IV|Ben hy kid w cr kid I-IV
C0155598|T047|AB|403.11|ICD9CM|Ben hyp kid w cr kid V|Ben hyp kid w cr kid V
C0848548|T047|HT|403.9|ICD9CM|Hypertensive renal disease, unspecified|Hypertensive renal disease, unspecified
C0494574|T047|AB|403.90|ICD9CM|Hy kid NOS w cr kid I-IV|Hy kid NOS w cr kid I-IV
C0348860|T047|AB|403.91|ICD9CM|Hyp kid NOS w cr kid V|Hyp kid NOS w cr kid V
C1719469|T047|HT|404|ICD9CM|Hypertensive heart and chronic kidney disease|Hypertensive heart and chronic kidney disease
C1719468|T047|HT|404.0|ICD9CM|Hypertensive heart and chronic kidney disease, malignant|Hypertensive heart and chronic kidney disease, malignant
C1719464|T047|AB|404.00|ICD9CM|Mal hy ht/kd I-IV w/o hf|Mal hy ht/kd I-IV w/o hf
C1719465|T047|AB|404.01|ICD9CM|Mal hyp ht/kd I-IV w hf|Mal hyp ht/kd I-IV w hf
C1719466|T047|AB|404.02|ICD9CM|Mal hy ht/kd st V w/o hf|Mal hy ht/kd st V w/o hf
C1719467|T047|AB|404.03|ICD9CM|Mal hyp ht/kd stg V w hf|Mal hyp ht/kd stg V w hf
C0155607|T047|HT|404.1|ICD9CM|Hypertensive heart and renal disease, benign|Hypertensive heart and renal disease, benign
C0155608|T047|AB|404.10|ICD9CM|Ben hy ht/kd I-IV w/o hf|Ben hy ht/kd I-IV w/o hf
C0155609|T047|AB|404.11|ICD9CM|Ben hyp ht/kd I-IV w hf|Ben hyp ht/kd I-IV w hf
C0155610|T047|AB|404.12|ICD9CM|Ben hy ht/kd st V w/o hf|Ben hy ht/kd st V w/o hf
C0155611|T047|AB|404.13|ICD9CM|Ben hyp ht/kd stg V w hf|Ben hyp ht/kd stg V w hf
C0155601|T047|HT|404.9|ICD9CM|Hypertensive heart and renal disease, unspecified|Hypertensive heart and renal disease, unspecified
C0155612|T047|AB|404.90|ICD9CM|Hy ht/kd NOS I-IV w/o hf|Hy ht/kd NOS I-IV w/o hf
C3665458|T047|AB|404.91|ICD9CM|Hyp ht/kd NOS I-IV w hf|Hyp ht/kd NOS I-IV w hf
C0348879|T047|AB|404.92|ICD9CM|Hy ht/kd NOS st V w/o hf|Hy ht/kd NOS st V w/o hf
C0494576|T047|AB|404.93|ICD9CM|Hyp ht/kd NOS st V w hf|Hyp ht/kd NOS st V w hf
C0155616|T047|HT|405|ICD9CM|Secondary hypertension|Secondary hypertension
C0155617|T047|HT|405.0|ICD9CM|Malignant secondary hypertension|Malignant secondary hypertension
C0264643|T047|AB|405.01|ICD9CM|Mal renovasc hypertens|Mal renovasc hypertens
C0264643|T047|PT|405.01|ICD9CM|Malignant renovascular hypertension|Malignant renovascular hypertension
C0155619|T047|AB|405.09|ICD9CM|Mal second hyperten NEC|Mal second hyperten NEC
C0155619|T047|PT|405.09|ICD9CM|Other malignant secondary hypertension|Other malignant secondary hypertension
C0155620|T047|HT|405.1|ICD9CM|Benign secondary hypertension|Benign secondary hypertension
C0155621|T047|AB|405.11|ICD9CM|Benign renovasc hyperten|Benign renovasc hyperten
C0155621|T047|PT|405.11|ICD9CM|Benign renovascular hypertension|Benign renovascular hypertension
C0155622|T047|AB|405.19|ICD9CM|Benign second hypert NEC|Benign second hypert NEC
C0155622|T047|PT|405.19|ICD9CM|Other benign secondary hypertension|Other benign secondary hypertension
C0155616|T047|HT|405.9|ICD9CM|Unspecified secondary hypertension|Unspecified secondary hypertension
C0155624|T047|AB|405.91|ICD9CM|Renovasc hypertension|Renovasc hypertension
C0155624|T047|PT|405.91|ICD9CM|Unspecified renovascular hypertension|Unspecified renovascular hypertension
C0348586|T047|PT|405.99|ICD9CM|Other unspecified secondary hypertension|Other unspecified secondary hypertension
C0348586|T047|AB|405.99|ICD9CM|Second hypertension NEC|Second hypertension NEC
C0155626|T047|HT|410|ICD9CM|Acute myocardial infarction|Acute myocardial infarction
C0151744|T047|HT|410-414.99|ICD9CM|ISCHEMIC HEART DISEASE|ISCHEMIC HEART DISEASE
C0155627|T047|HT|410.0|ICD9CM|Acute myocardial infarction, of anterolateral wall|Acute myocardial infarction, of anterolateral wall
C0155628|T047|PT|410.00|ICD9CM|Acute myocardial infarction of anterolateral wall, episode of care unspecified|Acute myocardial infarction of anterolateral wall, episode of care unspecified
C0155628|T047|AB|410.00|ICD9CM|AMI anterolateral,unspec|AMI anterolateral,unspec
C0155629|T047|PT|410.01|ICD9CM|Acute myocardial infarction of anterolateral wall, initial episode of care|Acute myocardial infarction of anterolateral wall, initial episode of care
C0155629|T047|AB|410.01|ICD9CM|AMI anterolateral, init|AMI anterolateral, init
C0155630|T047|PT|410.02|ICD9CM|Acute myocardial infarction of anterolateral wall, subsequent episode of care|Acute myocardial infarction of anterolateral wall, subsequent episode of care
C0155630|T047|AB|410.02|ICD9CM|AMI anterolateral,subseq|AMI anterolateral,subseq
C0155631|T047|HT|410.1|ICD9CM|Acute myocardial infarction, of other anterior wall|Acute myocardial infarction, of other anterior wall
C0155632|T047|PT|410.10|ICD9CM|Acute myocardial infarction of other anterior wall, episode of care unspecified|Acute myocardial infarction of other anterior wall, episode of care unspecified
C0155632|T047|AB|410.10|ICD9CM|AMI anterior wall,unspec|AMI anterior wall,unspec
C0155633|T047|PT|410.11|ICD9CM|Acute myocardial infarction of other anterior wall, initial episode of care|Acute myocardial infarction of other anterior wall, initial episode of care
C0155633|T047|AB|410.11|ICD9CM|AMI anterior wall, init|AMI anterior wall, init
C0155634|T047|PT|410.12|ICD9CM|Acute myocardial infarction of other anterior wall, subsequent episode of care|Acute myocardial infarction of other anterior wall, subsequent episode of care
C0155634|T047|AB|410.12|ICD9CM|AMI anterior wall,subseq|AMI anterior wall,subseq
C0340308|T047|HT|410.2|ICD9CM|Acute myocardial infarction, of inferolateral wall|Acute myocardial infarction, of inferolateral wall
C0155636|T047|PT|410.20|ICD9CM|Acute myocardial infarction of inferolateral wall, episode of care unspecified|Acute myocardial infarction of inferolateral wall, episode of care unspecified
C0155636|T047|AB|410.20|ICD9CM|AMI inferolateral,unspec|AMI inferolateral,unspec
C0155637|T047|PT|410.21|ICD9CM|Acute myocardial infarction of inferolateral wall, initial episode of care|Acute myocardial infarction of inferolateral wall, initial episode of care
C0155637|T047|AB|410.21|ICD9CM|AMI inferolateral, init|AMI inferolateral, init
C0155638|T047|PT|410.22|ICD9CM|Acute myocardial infarction of inferolateral wall, subsequent episode of care|Acute myocardial infarction of inferolateral wall, subsequent episode of care
C0155638|T047|AB|410.22|ICD9CM|AMI inferolateral,subseq|AMI inferolateral,subseq
C0340304|T047|HT|410.3|ICD9CM|Acute myocardial infarction, of inferoposterior wall|Acute myocardial infarction, of inferoposterior wall
C0155640|T047|PT|410.30|ICD9CM|Acute myocardial infarction of inferoposterior wall, episode of care unspecified|Acute myocardial infarction of inferoposterior wall, episode of care unspecified
C0155640|T047|AB|410.30|ICD9CM|AMI inferopost, unspec|AMI inferopost, unspec
C0155641|T047|PT|410.31|ICD9CM|Acute myocardial infarction of inferoposterior wall, initial episode of care|Acute myocardial infarction of inferoposterior wall, initial episode of care
C0155641|T047|AB|410.31|ICD9CM|AMI inferopost, initial|AMI inferopost, initial
C0155642|T047|PT|410.32|ICD9CM|Acute myocardial infarction of inferoposterior wall, subsequent episode of care|Acute myocardial infarction of inferoposterior wall, subsequent episode of care
C0155642|T047|AB|410.32|ICD9CM|AMI inferopost, subseq|AMI inferopost, subseq
C0155643|T047|HT|410.4|ICD9CM|Acute myocardial infarction, of other inferior wall|Acute myocardial infarction, of other inferior wall
C0155644|T047|PT|410.40|ICD9CM|Acute myocardial infarction of other inferior wall, episode of care unspecified|Acute myocardial infarction of other inferior wall, episode of care unspecified
C0155644|T047|AB|410.40|ICD9CM|AMI inferior wall,unspec|AMI inferior wall,unspec
C0155645|T047|PT|410.41|ICD9CM|Acute myocardial infarction of other inferior wall, initial episode of care|Acute myocardial infarction of other inferior wall, initial episode of care
C0155645|T047|AB|410.41|ICD9CM|AMI inferior wall, init|AMI inferior wall, init
C0155646|T047|PT|410.42|ICD9CM|Acute myocardial infarction of other inferior wall, subsequent episode of care|Acute myocardial infarction of other inferior wall, subsequent episode of care
C0155646|T047|AB|410.42|ICD9CM|AMI inferior wall,subseq|AMI inferior wall,subseq
C0155647|T047|HT|410.5|ICD9CM|Acute myocardial infarction, of other lateral wall|Acute myocardial infarction, of other lateral wall
C0155648|T047|PT|410.50|ICD9CM|Acute myocardial infarction of other lateral wall, episode of care unspecified|Acute myocardial infarction of other lateral wall, episode of care unspecified
C0155648|T047|AB|410.50|ICD9CM|AMI lateral NEC, unspec|AMI lateral NEC, unspec
C0155649|T047|PT|410.51|ICD9CM|Acute myocardial infarction of other lateral wall, initial episode of care|Acute myocardial infarction of other lateral wall, initial episode of care
C0155649|T047|AB|410.51|ICD9CM|AMI lateral NEC, initial|AMI lateral NEC, initial
C0155650|T047|PT|410.52|ICD9CM|Acute myocardial infarction of other lateral wall, subsequent episode of care|Acute myocardial infarction of other lateral wall, subsequent episode of care
C0155650|T047|AB|410.52|ICD9CM|AMI lateral NEC, subseq|AMI lateral NEC, subseq
C0264706|T047|HT|410.6|ICD9CM|Acute myocardial infarction, true posterior wall infarction|Acute myocardial infarction, true posterior wall infarction
C0155652|T047|AB|410.60|ICD9CM|True post infarct,unspec|True post infarct,unspec
C0155652|T047|PT|410.60|ICD9CM|True posterior wall infarction, episode of care unspecified|True posterior wall infarction, episode of care unspecified
C0155653|T047|AB|410.61|ICD9CM|True post infarct, init|True post infarct, init
C0155653|T047|PT|410.61|ICD9CM|True posterior wall infarction, initial episode of care|True posterior wall infarction, initial episode of care
C0155654|T047|AB|410.62|ICD9CM|True post infarct,subseq|True post infarct,subseq
C0155654|T047|PT|410.62|ICD9CM|True posterior wall infarction, subsequent episode of care|True posterior wall infarction, subsequent episode of care
C0155655|T047|HT|410.7|ICD9CM|Acute myocardial infarction, subendocardial infarction|Acute myocardial infarction, subendocardial infarction
C0494580|T047|AB|410.70|ICD9CM|Subendo infarct, unspec|Subendo infarct, unspec
C0494580|T047|PT|410.70|ICD9CM|Subendocardial infarction, episode of care unspecified|Subendocardial infarction, episode of care unspecified
C0155657|T047|AB|410.71|ICD9CM|Subendo infarct, initial|Subendo infarct, initial
C0155657|T047|PT|410.71|ICD9CM|Subendocardial infarction, initial episode of care|Subendocardial infarction, initial episode of care
C0155658|T047|AB|410.72|ICD9CM|Subendo infarct, subseq|Subendo infarct, subseq
C0155658|T047|PT|410.72|ICD9CM|Subendocardial infarction, subsequent episode of care|Subendocardial infarction, subsequent episode of care
C0155659|T047|HT|410.8|ICD9CM|Acute myocardial infarction, of other specified sites|Acute myocardial infarction, of other specified sites
C0155660|T047|PT|410.80|ICD9CM|Acute myocardial infarction of other specified sites, episode of care unspecified|Acute myocardial infarction of other specified sites, episode of care unspecified
C0155660|T047|AB|410.80|ICD9CM|AMI NEC, unspecified|AMI NEC, unspecified
C0155661|T047|PT|410.81|ICD9CM|Acute myocardial infarction of other specified sites, initial episode of care|Acute myocardial infarction of other specified sites, initial episode of care
C0155661|T047|AB|410.81|ICD9CM|AMI NEC, initial|AMI NEC, initial
C0155662|T047|PT|410.82|ICD9CM|Acute myocardial infarction of other specified sites, subsequent episode of care|Acute myocardial infarction of other specified sites, subsequent episode of care
C0155662|T047|AB|410.82|ICD9CM|AMI NEC, subsequent|AMI NEC, subsequent
C0155626|T047|HT|410.9|ICD9CM|Acute myocardial infarction, unspecified site|Acute myocardial infarction, unspecified site
C0155626|T047|PT|410.90|ICD9CM|Acute myocardial infarction of unspecified site, episode of care unspecified|Acute myocardial infarction of unspecified site, episode of care unspecified
C0155626|T047|AB|410.90|ICD9CM|AMI NOS, unspecified|AMI NOS, unspecified
C0155664|T047|PT|410.91|ICD9CM|Acute myocardial infarction of unspecified site, initial episode of care|Acute myocardial infarction of unspecified site, initial episode of care
C0155664|T047|AB|410.91|ICD9CM|AMI NOS, initial|AMI NOS, initial
C0155665|T047|PT|410.92|ICD9CM|Acute myocardial infarction of unspecified site, subsequent episode of care|Acute myocardial infarction of unspecified site, subsequent episode of care
C0155665|T047|AB|410.92|ICD9CM|AMI NOS, subsequent|AMI NOS, subsequent
C0340283|T047|HT|411|ICD9CM|Other acute and subacute forms of ischemic heart disease|Other acute and subacute forms of ischemic heart disease
C0152107|T047|AB|411.0|ICD9CM|Post MI syndrome|Post MI syndrome
C0152107|T047|PT|411.0|ICD9CM|Postmyocardial infarction syndrome|Postmyocardial infarction syndrome
C0002965|T047|AB|411.1|ICD9CM|Intermed coronary synd|Intermed coronary synd
C0002965|T047|PT|411.1|ICD9CM|Intermediate coronary syndrome|Intermediate coronary syndrome
C0340283|T047|HT|411.8|ICD9CM|Other acute and subacute forms of ischemic heart disease|Other acute and subacute forms of ischemic heart disease
C0949167|T047|AB|411.81|ICD9CM|Acute cor occlsn w/o MI|Acute cor occlsn w/o MI
C0949167|T047|PT|411.81|ICD9CM|Acute coronary occlusion without myocardial infarction|Acute coronary occlusion without myocardial infarction
C0340283|T047|AB|411.89|ICD9CM|Ac ischemic hrt dis NEC|Ac ischemic hrt dis NEC
C0340283|T047|PT|411.89|ICD9CM|Other acute and subacute forms of ischemic heart disease, other|Other acute and subacute forms of ischemic heart disease, other
C0155668|T047|AB|412|ICD9CM|Old myocardial infarct|Old myocardial infarct
C0155668|T047|PT|412|ICD9CM|Old myocardial infarction|Old myocardial infarction
C0002962|T184|HT|413|ICD9CM|Angina pectoris|Angina pectoris
C0152172|T047|AB|413.0|ICD9CM|Angina decubitus|Angina decubitus
C0152172|T047|PT|413.0|ICD9CM|Angina decubitus|Angina decubitus
C0002963|T047|AB|413.1|ICD9CM|Prinzmetal angina|Prinzmetal angina
C0002963|T047|PT|413.1|ICD9CM|Prinzmetal angina|Prinzmetal angina
C0348588|T184|AB|413.9|ICD9CM|Angina pectoris NEC/NOS|Angina pectoris NEC/NOS
C0348588|T184|PT|413.9|ICD9CM|Other and unspecified angina pectoris|Other and unspecified angina pectoris
C0155669|T047|HT|414|ICD9CM|Other forms of chronic ischemic heart disease|Other forms of chronic ischemic heart disease
C0010054|T047|HT|414.0|ICD9CM|Coronary atherosclerosis|Coronary atherosclerosis
C0837133|T047|AB|414.00|ICD9CM|Cor ath unsp vsl ntv/gft|Cor ath unsp vsl ntv/gft
C0837133|T047|PT|414.00|ICD9CM|Coronary atherosclerosis of unspecified type of vessel, native or graft|Coronary atherosclerosis of unspecified type of vessel, native or graft
C0837134|T047|PT|414.01|ICD9CM|Coronary atherosclerosis of native coronary artery|Coronary atherosclerosis of native coronary artery
C0837134|T047|AB|414.01|ICD9CM|Crnry athrscl natve vssl|Crnry athrscl natve vssl
C0837135|T047|PT|414.02|ICD9CM|Coronary atherosclerosis of autologous vein bypass graft|Coronary atherosclerosis of autologous vein bypass graft
C0837135|T047|AB|414.02|ICD9CM|Crn ath atlg vn bps grft|Crn ath atlg vn bps grft
C0837136|T047|PT|414.03|ICD9CM|Coronary atherosclerosis of nonautologous biological bypass graft|Coronary atherosclerosis of nonautologous biological bypass graft
C0837136|T047|AB|414.03|ICD9CM|Crn ath nonatlg blg grft|Crn ath nonatlg blg grft
C0375264|T047|AB|414.04|ICD9CM|Cor ath artry bypas grft|Cor ath artry bypas grft
C0375264|T047|PT|414.04|ICD9CM|Coronary atherosclerosis of artery bypass graft|Coronary atherosclerosis of artery bypass graft
C0375265|T047|AB|414.05|ICD9CM|Cor ath bypass graft NOS|Cor ath bypass graft NOS
C0375265|T047|PT|414.05|ICD9CM|Coronary atherosclerosis of unspecified bypass graft|Coronary atherosclerosis of unspecified bypass graft
C1135190|T047|AB|414.06|ICD9CM|Cor ath natv art tp hrt|Cor ath natv art tp hrt
C1135190|T047|PT|414.06|ICD9CM|Coronary atherosclerosis of native coronary artery of transplanted heart|Coronary atherosclerosis of native coronary artery of transplanted heart
C1456095|T047|AB|414.07|ICD9CM|Cor ath bps graft tp hrt|Cor ath bps graft tp hrt
C1456095|T047|PT|414.07|ICD9CM|Coronary atherosclerosis of bypass graft (artery) (vein) of transplanted heart|Coronary atherosclerosis of bypass graft (artery) (vein) of transplanted heart
C1135334|T047|HT|414.1|ICD9CM|Aneurysm and dissection of heart|Aneurysm and dissection of heart
C1541919|T047|AB|414.10|ICD9CM|Aneurysm of heart|Aneurysm of heart
C1541919|T047|PT|414.10|ICD9CM|Aneurysm of heart (wall)|Aneurysm of heart (wall)
C0010051|T047|AB|414.11|ICD9CM|Aneurysm coronary vessel|Aneurysm coronary vessel
C0010051|T047|PT|414.11|ICD9CM|Aneurysm of coronary vessels|Aneurysm of coronary vessels
C0340648|T047|AB|414.12|ICD9CM|Dissection cor artery|Dissection cor artery
C0340648|T047|PT|414.12|ICD9CM|Dissection of coronary artery|Dissection of coronary artery
C0029519|T047|AB|414.19|ICD9CM|Aneurysm of heart NEC|Aneurysm of heart NEC
C0029519|T047|PT|414.19|ICD9CM|Other aneurysm of heart|Other aneurysm of heart
C1955779|T047|AB|414.2|ICD9CM|Chr tot occlus cor artry|Chr tot occlus cor artry
C1955779|T047|PT|414.2|ICD9CM|Chronic total occlusion of coronary artery|Chronic total occlusion of coronary artery
C2349509|T047|AB|414.3|ICD9CM|Cor ath d/t lpd rch plaq|Cor ath d/t lpd rch plaq
C2349509|T047|PT|414.3|ICD9CM|Coronary atherosclerosis due to lipid rich plaque|Coronary atherosclerosis due to lipid rich plaque
C3161090|T047|AB|414.4|ICD9CM|Cor ath d/t calc cor lsn|Cor ath d/t calc cor lsn
C3161090|T047|PT|414.4|ICD9CM|Coronary atherosclerosis due to calcified coronary lesion|Coronary atherosclerosis due to calcified coronary lesion
C0155670|T047|AB|414.8|ICD9CM|Chr ischemic hrt dis NEC|Chr ischemic hrt dis NEC
C0155670|T047|PT|414.8|ICD9CM|Other specified forms of chronic ischemic heart disease|Other specified forms of chronic ischemic heart disease
C0264694|T047|AB|414.9|ICD9CM|Chr ischemic hrt dis NOS|Chr ischemic hrt dis NOS
C0264694|T047|PT|414.9|ICD9CM|Chronic ischemic heart disease, unspecified|Chronic ischemic heart disease, unspecified
C0155671|T047|HT|415|ICD9CM|Acute pulmonary heart disease|Acute pulmonary heart disease
C0178272|T047|HT|415-417.99|ICD9CM|DISEASES OF PULMONARY CIRCULATION|DISEASES OF PULMONARY CIRCULATION
C0155672|T047|AB|415.0|ICD9CM|Acute cor pulmonale|Acute cor pulmonale
C0155672|T047|PT|415.0|ICD9CM|Acute cor pulmonale|Acute cor pulmonale
C0034066|T047|HT|415.1|ICD9CM|Pulmonary embolism and infarction|Pulmonary embolism and infarction
C2711829|T047|AB|415.11|ICD9CM|Iatrogen pulm emb/infarc|Iatrogen pulm emb/infarc
C2711829|T047|PT|415.11|ICD9CM|Iatrogenic pulmonary embolism and infarction|Iatrogenic pulmonary embolism and infarction
C1955781|T046|PT|415.12|ICD9CM|Septic pulmonary embolism|Septic pulmonary embolism
C1955781|T046|AB|415.12|ICD9CM|Septic pulmonary embolsm|Septic pulmonary embolsm
C3161091|T047|AB|415.13|ICD9CM|Saddle embol pulmon art|Saddle embol pulmon art
C3161091|T047|PT|415.13|ICD9CM|Saddle embolus of pulmonary artery|Saddle embolus of pulmonary artery
C0375267|T047|PT|415.19|ICD9CM|Other pulmonary embolism and infarction|Other pulmonary embolism and infarction
C0375267|T047|AB|415.19|ICD9CM|Pulm embol/infarct NEC|Pulm embol/infarct NEC
C0238074|T047|HT|416|ICD9CM|Chronic pulmonary heart disease|Chronic pulmonary heart disease
C0152171|T047|AB|416.0|ICD9CM|Prim pulm hypertension|Prim pulm hypertension
C0152171|T047|PT|416.0|ICD9CM|Primary pulmonary hypertension|Primary pulmonary hypertension
C0152102|T047|AB|416.1|ICD9CM|Kyphoscoliotic heart dis|Kyphoscoliotic heart dis
C0152102|T047|PT|416.1|ICD9CM|Kyphoscoliotic heart disease|Kyphoscoliotic heart disease
C0856722|T046|AB|416.2|ICD9CM|Chr pulmonary embolism|Chr pulmonary embolism
C0856722|T046|PT|416.2|ICD9CM|Chronic pulmonary embolism|Chronic pulmonary embolism
C0155673|T047|AB|416.8|ICD9CM|Chr pulmon heart dis NEC|Chr pulmon heart dis NEC
C0155673|T047|PT|416.8|ICD9CM|Other chronic pulmonary heart diseases|Other chronic pulmonary heart diseases
C0238074|T047|AB|416.9|ICD9CM|Chr pulmon heart dis NOS|Chr pulmon heart dis NOS
C0238074|T047|PT|416.9|ICD9CM|Chronic pulmonary heart disease, unspecified|Chronic pulmonary heart disease, unspecified
C0155674|T047|HT|417|ICD9CM|Other diseases of pulmonary circulation|Other diseases of pulmonary circulation
C0155675|T047|AB|417.0|ICD9CM|Arterioven fistu pul ves|Arterioven fistu pul ves
C0155675|T047|PT|417.0|ICD9CM|Arteriovenous fistula of pulmonary vessels|Arteriovenous fistula of pulmonary vessels
C0155676|T046|PT|417.1|ICD9CM|Aneurysm of pulmonary artery|Aneurysm of pulmonary artery
C0155676|T046|AB|417.1|ICD9CM|Pulmon artery aneurysm|Pulmon artery aneurysm
C0155677|T047|PT|417.8|ICD9CM|Other specified diseases of pulmonary circulation|Other specified diseases of pulmonary circulation
C0155677|T047|AB|417.8|ICD9CM|Pulmon circulat dis NEC|Pulmon circulat dis NEC
C0178272|T047|AB|417.9|ICD9CM|Pulmon circulat dis NOS|Pulmon circulat dis NOS
C0178272|T047|PT|417.9|ICD9CM|Unspecified disease of pulmonary circulation|Unspecified disease of pulmonary circulation
C0155679|T047|HT|420|ICD9CM|Acute pericarditis|Acute pericarditis
C0178273|T047|HT|420-429.99|ICD9CM|OTHER FORMS OF HEART DISEASE|OTHER FORMS OF HEART DISEASE
C0340443|T047|AB|420.0|ICD9CM|Ac pericardit in oth dis|Ac pericardit in oth dis
C0340443|T047|PT|420.0|ICD9CM|Acute pericarditis in diseases classified elsewhere|Acute pericarditis in diseases classified elsewhere
C0155680|T047|HT|420.9|ICD9CM|Other and unspecified acute pericarditis|Other and unspecified acute pericarditis
C0155679|T047|AB|420.90|ICD9CM|Acute pericarditis NOS|Acute pericarditis NOS
C0155679|T047|PT|420.90|ICD9CM|Acute pericarditis, unspecified|Acute pericarditis, unspecified
C0155681|T047|AB|420.91|ICD9CM|Ac idiopath pericarditis|Ac idiopath pericarditis
C0155681|T047|PT|420.91|ICD9CM|Acute idiopathic pericarditis|Acute idiopathic pericarditis
C0348597|T047|AB|420.99|ICD9CM|Acute pericarditis NEC|Acute pericarditis NEC
C0348597|T047|PT|420.99|ICD9CM|Other acute pericarditis|Other acute pericarditis
C0155683|T047|HT|421|ICD9CM|Acute and subacute endocarditis|Acute and subacute endocarditis
C0553977|T047|AB|421.0|ICD9CM|Ac/subac bact endocard|Ac/subac bact endocard
C0553977|T047|PT|421.0|ICD9CM|Acute and subacute bacterial endocarditis|Acute and subacute bacterial endocarditis
C0340348|T047|AB|421.1|ICD9CM|Ac endocardit in oth dis|Ac endocardit in oth dis
C0340348|T047|PT|421.1|ICD9CM|Acute and subacute infective endocarditis in diseases classified elsewhere|Acute and subacute infective endocarditis in diseases classified elsewhere
C0375268|T047|AB|421.9|ICD9CM|Ac/subac endocardit NOS|Ac/subac endocardit NOS
C0375268|T047|PT|421.9|ICD9CM|Acute endocarditis, unspecified|Acute endocarditis, unspecified
C0155686|T047|HT|422|ICD9CM|Acute myocarditis|Acute myocarditis
C0155687|T047|AB|422.0|ICD9CM|Ac myocardit in oth dis|Ac myocardit in oth dis
C0155687|T047|PT|422.0|ICD9CM|Acute myocarditis in diseases classified elsewhere|Acute myocarditis in diseases classified elsewhere
C0155692|T047|HT|422.9|ICD9CM|Other and unspecified acute myocarditis|Other and unspecified acute myocarditis
C0155686|T047|AB|422.90|ICD9CM|Acute myocarditis NOS|Acute myocarditis NOS
C0155686|T047|PT|422.90|ICD9CM|Acute myocarditis, unspecified|Acute myocarditis, unspecified
C0155689|T047|AB|422.91|ICD9CM|Idiopathic myocarditis|Idiopathic myocarditis
C0155689|T047|PT|422.91|ICD9CM|Idiopathic myocarditis|Idiopathic myocarditis
C0155690|T047|AB|422.92|ICD9CM|Septic myocarditis|Septic myocarditis
C0155690|T047|PT|422.92|ICD9CM|Septic myocarditis|Septic myocarditis
C0155691|T047|AB|422.93|ICD9CM|Toxic myocarditis|Toxic myocarditis
C0155691|T047|PT|422.93|ICD9CM|Toxic myocarditis|Toxic myocarditis
C0155692|T047|AB|422.99|ICD9CM|Acute myocarditis NEC|Acute myocarditis NEC
C0155692|T047|PT|422.99|ICD9CM|Other acute myocarditis|Other acute myocarditis
C0340442|T047|HT|423|ICD9CM|Other diseases of pericardium|Other diseases of pericardium
C0019064|T046|AB|423.0|ICD9CM|Hemopericardium|Hemopericardium
C0019064|T046|PT|423.0|ICD9CM|Hemopericardium|Hemopericardium
C0152452|T047|AB|423.1|ICD9CM|Adhesive pericarditis|Adhesive pericarditis
C0152452|T047|PT|423.1|ICD9CM|Adhesive pericarditis|Adhesive pericarditis
C0031048|T047|AB|423.2|ICD9CM|Constrictiv pericarditis|Constrictiv pericarditis
C0031048|T047|PT|423.2|ICD9CM|Constrictive pericarditis|Constrictive pericarditis
C0007177|T047|PT|423.3|ICD9CM|Cardiac tamponade|Cardiac tamponade
C0007177|T047|AB|423.3|ICD9CM|Cardiac tamponade|Cardiac tamponade
C0155694|T047|PT|423.8|ICD9CM|Other specified diseases of pericardium|Other specified diseases of pericardium
C0155694|T047|AB|423.8|ICD9CM|Pericardial disease NEC|Pericardial disease NEC
C0265122|T047|AB|423.9|ICD9CM|Pericardial disease NOS|Pericardial disease NOS
C0265122|T047|PT|423.9|ICD9CM|Unspecified disease of pericardium|Unspecified disease of pericardium
C0155695|T047|HT|424|ICD9CM|Other diseases of endocardium|Other diseases of endocardium
C0026265|T047|AB|424.0|ICD9CM|Mitral valve disorder|Mitral valve disorder
C0026265|T047|PT|424.0|ICD9CM|Mitral valve disorders|Mitral valve disorders
C1260873|T047|AB|424.1|ICD9CM|Aortic valve disorder|Aortic valve disorder
C1260873|T047|PT|424.1|ICD9CM|Aortic valve disorders|Aortic valve disorders
C0701168|T047|AB|424.2|ICD9CM|Nonrheum tricusp val dis|Nonrheum tricusp val dis
C0701168|T047|PT|424.2|ICD9CM|Tricuspid valve disorders, specified as nonrheumatic|Tricuspid valve disorders, specified as nonrheumatic
C0034087|T047|AB|424.3|ICD9CM|Pulmonary valve disorder|Pulmonary valve disorder
C0034087|T047|PT|424.3|ICD9CM|Pulmonary valve disorders|Pulmonary valve disorders
C0264865|T047|HT|424.9|ICD9CM|Endocarditis, valve unspecified|Endocarditis, valve unspecified
C0264865|T047|AB|424.90|ICD9CM|Endocarditis NOS|Endocarditis NOS
C0264865|T047|PT|424.90|ICD9CM|Endocarditis, valve unspecified, unspecified cause|Endocarditis, valve unspecified, unspecified cause
C0340345|T047|PT|424.91|ICD9CM|Endocarditis in diseases classified elsewhere|Endocarditis in diseases classified elsewhere
C0340345|T047|AB|424.91|ICD9CM|Endocarditis in oth dis|Endocarditis in oth dis
C0029609|T047|AB|424.99|ICD9CM|Endocarditis NEC|Endocarditis NEC
C0029609|T047|PT|424.99|ICD9CM|Other endocarditis, valve unspecified|Other endocarditis, valve unspecified
C0878544|T047|HT|425|ICD9CM|Cardiomyopathy|Cardiomyopathy
C0553980|T046|AB|425.0|ICD9CM|Endomyocardial fibrosis|Endomyocardial fibrosis
C0553980|T046|PT|425.0|ICD9CM|Endomyocardial fibrosis|Endomyocardial fibrosis
C0007194|T047|HT|425.1|ICD9CM|Hypertrophic cardiomyopathy|Hypertrophic cardiomyopathy
C4551472|T047|PT|425.11|ICD9CM|Hypertrophic obstructive cardiomyopathy|Hypertrophic obstructive cardiomyopathy
C4551472|T047|AB|425.11|ICD9CM|Hyprtrophc obst cardiomy|Hyprtrophc obst cardiomy
C0348615|T047|AB|425.18|ICD9CM|Oth hyprtrophic cardiomy|Oth hyprtrophic cardiomy
C0348615|T047|PT|425.18|ICD9CM|Other hypertrophic cardiomyopathy|Other hypertrophic cardiomyopathy
C1959600|T047|AB|425.2|ICD9CM|Obsc afric cardiomyopath|Obsc afric cardiomyopath
C1959600|T047|PT|425.2|ICD9CM|Obscure cardiomyopathy of Africa|Obscure cardiomyopathy of Africa
C0014117|T047|AB|425.3|ICD9CM|Endocard fibroelastosis|Endocard fibroelastosis
C0014117|T047|PT|425.3|ICD9CM|Endocardial fibroelastosis|Endocardial fibroelastosis
C0340419|T047|PT|425.4|ICD9CM|Other primary cardiomyopathies|Other primary cardiomyopathies
C0340419|T047|AB|425.4|ICD9CM|Prim cardiomyopathy NEC|Prim cardiomyopathy NEC
C0007192|T047|AB|425.5|ICD9CM|Alcoholic cardiomyopathy|Alcoholic cardiomyopathy
C0007192|T047|PT|425.5|ICD9CM|Alcoholic cardiomyopathy|Alcoholic cardiomyopathy
C0340422|T047|AB|425.7|ICD9CM|Metabolic cardiomyopathy|Metabolic cardiomyopathy
C0340422|T047|PT|425.7|ICD9CM|Nutritional and metabolic cardiomyopathy|Nutritional and metabolic cardiomyopathy
C0155699|T047|AB|425.8|ICD9CM|Cardiomyopath in oth dis|Cardiomyopath in oth dis
C0155699|T047|PT|425.8|ICD9CM|Cardiomyopathy in other diseases classified elsewhere|Cardiomyopathy in other diseases classified elsewhere
C0036529|T047|AB|425.9|ICD9CM|Second cardiomyopath NOS|Second cardiomyopath NOS
C0036529|T047|PT|425.9|ICD9CM|Secondary cardiomyopathy, unspecified|Secondary cardiomyopathy, unspecified
C0264886|T047|HT|426|ICD9CM|Conduction disorders|Conduction disorders
C0151517|T047|AB|426.0|ICD9CM|Atriovent block complete|Atriovent block complete
C0151517|T047|PT|426.0|ICD9CM|Atrioventricular block, complete|Atrioventricular block, complete
C0348621|T046|HT|426.1|ICD9CM|Atrioventricular block, other and unspecified|Atrioventricular block, other and unspecified
C0004245|T047|AB|426.10|ICD9CM|Atriovent block NOS|Atriovent block NOS
C0004245|T047|PT|426.10|ICD9CM|Atrioventricular block, unspecified|Atrioventricular block, unspecified
C0085614|T047|AB|426.11|ICD9CM|Atriovent block-1st degr|Atriovent block-1st degr
C0085614|T047|PT|426.11|ICD9CM|First degree atrioventricular block|First degree atrioventricular block
C0155700|T047|AB|426.12|ICD9CM|Atrioven block-mobitz ii|Atrioven block-mobitz ii
C0155700|T047|PT|426.12|ICD9CM|Mobitz (type) II atrioventricular block|Mobitz (type) II atrioventricular block
C0549211|T047|AB|426.13|ICD9CM|Av block-2nd degree NEC|Av block-2nd degree NEC
C0549211|T047|PT|426.13|ICD9CM|Other second degree atrioventricular block|Other second degree atrioventricular block
C0155702|T047|AB|426.2|ICD9CM|Left bb hemiblock|Left bb hemiblock
C0155702|T047|PT|426.2|ICD9CM|Left bundle branch hemiblock|Left bundle branch hemiblock
C0155703|T047|AB|426.3|ICD9CM|Left bb block NEC|Left bb block NEC
C0155703|T047|PT|426.3|ICD9CM|Other left bundle branch block|Other left bundle branch block
C0085615|T047|PT|426.4|ICD9CM|Right bundle branch block|Right bundle branch block
C0085615|T047|AB|426.4|ICD9CM|Rt bundle branch block|Rt bundle branch block
C0677586|T046|HT|426.5|ICD9CM|Bundle branch block, other and unspecified|Bundle branch block, other and unspecified
C0006384|T047|AB|426.50|ICD9CM|Bundle branch block NOS|Bundle branch block NOS
C0006384|T047|PT|426.50|ICD9CM|Bundle branch block, unspecified|Bundle branch block, unspecified
C0155704|T047|PT|426.51|ICD9CM|Right bundle branch block and left posterior fascicular block|Right bundle branch block and left posterior fascicular block
C0155704|T047|AB|426.51|ICD9CM|Rt bbb/lft post fasc blk|Rt bbb/lft post fasc blk
C0155705|T047|PT|426.52|ICD9CM|Right bundle branch block and left anterior fascicular block|Right bundle branch block and left anterior fascicular block
C0155705|T047|AB|426.52|ICD9CM|Rt bbb/lft ant fasc blk|Rt bbb/lft ant fasc blk
C0155706|T046|AB|426.53|ICD9CM|Bilat bb block NEC|Bilat bb block NEC
C0155706|T046|PT|426.53|ICD9CM|Other bilateral bundle branch block|Other bilateral bundle branch block
C0155707|T047|AB|426.54|ICD9CM|Trifascicular block|Trifascicular block
C0155707|T047|PT|426.54|ICD9CM|Trifascicular block|Trifascicular block
C0029630|T046|AB|426.6|ICD9CM|Other heart block|Other heart block
C0029630|T046|PT|426.6|ICD9CM|Other heart block|Other heart block
C0392470|T047|PT|426.7|ICD9CM|Anomalous atrioventricular excitation|Anomalous atrioventricular excitation
C0392470|T047|AB|426.7|ICD9CM|Anomalous av excitation|Anomalous av excitation
C0155708|T046|HT|426.8|ICD9CM|Other specified conduction disorders|Other specified conduction disorders
C0024054|T047|AB|426.81|ICD9CM|Lown-ganong-levine synd|Lown-ganong-levine synd
C0024054|T047|PT|426.81|ICD9CM|Lown-Ganong-Levine syndrome|Lown-Ganong-Levine syndrome
C0023976|T047|AB|426.82|ICD9CM|Long QT syndrome|Long QT syndrome
C0023976|T047|PT|426.82|ICD9CM|Long QT syndrome|Long QT syndrome
C0155708|T046|AB|426.89|ICD9CM|Conduction disorder NEC|Conduction disorder NEC
C0155708|T046|PT|426.89|ICD9CM|Other specified conduction disorders|Other specified conduction disorders
C0264886|T047|AB|426.9|ICD9CM|Conduction disorder NOS|Conduction disorder NOS
C0264886|T047|PT|426.9|ICD9CM|Conduction disorder, unspecified|Conduction disorder, unspecified
C0003811|T047|HT|427|ICD9CM|Cardiac dysrhythmias|Cardiac dysrhythmias
C0030590|T047|AB|427.0|ICD9CM|Parox atrial tachycardia|Parox atrial tachycardia
C0030590|T047|PT|427.0|ICD9CM|Paroxysmal supraventricular tachycardia|Paroxysmal supraventricular tachycardia
C0030591|T047|AB|427.1|ICD9CM|Parox ventric tachycard|Parox ventric tachycard
C0030591|T047|PT|427.1|ICD9CM|Paroxysmal ventricular tachycardia|Paroxysmal ventricular tachycardia
C0039236|T047|AB|427.2|ICD9CM|Parox tachycardia NOS|Parox tachycardia NOS
C0039236|T047|PT|427.2|ICD9CM|Paroxysmal tachycardia, unspecified|Paroxysmal tachycardia, unspecified
C0155709|T046|HT|427.3|ICD9CM|Atrial fibrillation and flutter|Atrial fibrillation and flutter
C0004238|T047|AB|427.31|ICD9CM|Atrial fibrillation|Atrial fibrillation
C0004238|T047|PT|427.31|ICD9CM|Atrial fibrillation|Atrial fibrillation
C0004239|T046|AB|427.32|ICD9CM|Atrial flutter|Atrial flutter
C0004239|T046|PT|427.32|ICD9CM|Atrial flutter|Atrial flutter
C0155710|T046|HT|427.4|ICD9CM|Ventricular fibrillation and flutter|Ventricular fibrillation and flutter
C0042510|T047|AB|427.41|ICD9CM|Ventricular fibrillation|Ventricular fibrillation
C0042510|T047|PT|427.41|ICD9CM|Ventricular fibrillation|Ventricular fibrillation
C0152173|T047|AB|427.42|ICD9CM|Ventricular flutter|Ventricular flutter
C0152173|T047|PT|427.42|ICD9CM|Ventricular flutter|Ventricular flutter
C0018790|T047|AB|427.5|ICD9CM|Cardiac arrest|Cardiac arrest
C0018790|T047|PT|427.5|ICD9CM|Cardiac arrest|Cardiac arrest
C0340464|T047|HT|427.6|ICD9CM|Premature beats|Premature beats
C0340464|T047|AB|427.60|ICD9CM|Premature beats NOS|Premature beats NOS
C0340464|T047|PT|427.60|ICD9CM|Premature beats, unspecified|Premature beats, unspecified
C0033036|T047|AB|427.61|ICD9CM|Atrial premature beats|Atrial premature beats
C0033036|T047|PT|427.61|ICD9CM|Supraventricular premature beats|Supraventricular premature beats
C0029712|T046|PT|427.69|ICD9CM|Other premature beats|Other premature beats
C0029712|T046|AB|427.69|ICD9CM|Premature beats NEC|Premature beats NEC
C0348626|T047|HT|427.8|ICD9CM|Other specified cardiac dysrhythmias|Other specified cardiac dysrhythmias
C0428908|T047|AB|427.81|ICD9CM|Sinoatrial node dysfunct|Sinoatrial node dysfunct
C0428908|T047|PT|427.81|ICD9CM|Sinoatrial node dysfunction|Sinoatrial node dysfunction
C0348626|T047|AB|427.89|ICD9CM|Cardiac dysrhythmias NEC|Cardiac dysrhythmias NEC
C0348626|T047|PT|427.89|ICD9CM|Other specified cardiac dysrhythmias|Other specified cardiac dysrhythmias
C0003811|T047|AB|427.9|ICD9CM|Cardiac dysrhythmia NOS|Cardiac dysrhythmia NOS
C0003811|T047|PT|427.9|ICD9CM|Cardiac dysrhythmia, unspecified|Cardiac dysrhythmia, unspecified
C0018801|T047|HT|428|ICD9CM|Heart failure|Heart failure
C0018802|T047|AB|428.0|ICD9CM|CHF NOS|CHF NOS
C0018802|T047|PT|428.0|ICD9CM|Congestive heart failure, unspecified|Congestive heart failure, unspecified
C0023212|T047|AB|428.1|ICD9CM|Left heart failure|Left heart failure
C0023212|T047|PT|428.1|ICD9CM|Left heart failure|Left heart failure
C1135191|T047|HT|428.2|ICD9CM|Systolic heart failure|Systolic heart failure
C1135191|T047|PT|428.20|ICD9CM|Systolic heart failure, unspecified|Systolic heart failure, unspecified
C1135191|T047|AB|428.20|ICD9CM|Systolic hrt failure NOS|Systolic hrt failure NOS
C2732748|T047|AB|428.21|ICD9CM|Ac systolic hrt failure|Ac systolic hrt failure
C2732748|T047|PT|428.21|ICD9CM|Acute systolic heart failure|Acute systolic heart failure
C1135194|T047|AB|428.22|ICD9CM|Chr systolic hrt failure|Chr systolic hrt failure
C1135194|T047|PT|428.22|ICD9CM|Chronic systolic heart failure|Chronic systolic heart failure
C2733492|T047|AB|428.23|ICD9CM|Ac on chr syst hrt fail|Ac on chr syst hrt fail
C2733492|T047|PT|428.23|ICD9CM|Acute on chronic systolic heart failure|Acute on chronic systolic heart failure
C1135196|T047|HT|428.3|ICD9CM|Diastolic heart failure|Diastolic heart failure
C1135196|T047|AB|428.30|ICD9CM|Diastolc hrt failure NOS|Diastolc hrt failure NOS
C1135196|T047|PT|428.30|ICD9CM|Diastolic heart failure, unspecified|Diastolic heart failure, unspecified
C2732951|T047|AB|428.31|ICD9CM|Ac diastolic hrt failure|Ac diastolic hrt failure
C2732951|T047|PT|428.31|ICD9CM|Acute diastolic heart failure|Acute diastolic heart failure
C2711480|T047|AB|428.32|ICD9CM|Chr diastolic hrt fail|Chr diastolic hrt fail
C2711480|T047|PT|428.32|ICD9CM|Chronic diastolic heart failure|Chronic diastolic heart failure
C2732749|T047|AB|428.33|ICD9CM|Ac on chr diast hrt fail|Ac on chr diast hrt fail
C2732749|T047|PT|428.33|ICD9CM|Acute on chronic diastolic heart failure|Acute on chronic diastolic heart failure
C2882273|T047|HT|428.4|ICD9CM|Combined systolic and diastolic heart failure|Combined systolic and diastolic heart failure
C2882273|T047|PT|428.40|ICD9CM|Combined systolic and diastolic heart failure, unspecified|Combined systolic and diastolic heart failure, unspecified
C2882273|T047|AB|428.40|ICD9CM|Syst/diast hrt fail NOS|Syst/diast hrt fail NOS
C2882274|T047|AB|428.41|ICD9CM|Ac syst/diastol hrt fail|Ac syst/diastol hrt fail
C2882274|T047|PT|428.41|ICD9CM|Acute combined systolic and diastolic heart failure|Acute combined systolic and diastolic heart failure
C2882275|T047|AB|428.42|ICD9CM|Chr syst/diastl hrt fail|Chr syst/diastl hrt fail
C2882275|T047|PT|428.42|ICD9CM|Chronic combined systolic and diastolic heart failure|Chronic combined systolic and diastolic heart failure
C2882276|T047|AB|428.43|ICD9CM|Ac/chr syst/dia hrt fail|Ac/chr syst/dia hrt fail
C2882276|T047|PT|428.43|ICD9CM|Acute on chronic combined systolic and diastolic heart failure|Acute on chronic combined systolic and diastolic heart failure
C0018801|T047|AB|428.9|ICD9CM|Heart failure NOS|Heart failure NOS
C0018801|T047|PT|428.9|ICD9CM|Heart failure, unspecified|Heart failure, unspecified
C0155711|T046|HT|429|ICD9CM|Ill-defined descriptions and complications of heart disease|Ill-defined descriptions and complications of heart disease
C0027059|T047|AB|429.0|ICD9CM|Myocarditis NOS|Myocarditis NOS
C0027059|T047|PT|429.0|ICD9CM|Myocarditis, unspecified|Myocarditis, unspecified
C0027046|T046|AB|429.1|ICD9CM|Myocardial degeneration|Myocardial degeneration
C0027046|T046|PT|429.1|ICD9CM|Myocardial degeneration|Myocardial degeneration
C0007222|T047|AB|429.2|ICD9CM|Ascvd|Ascvd
C0007222|T047|PT|429.2|ICD9CM|Cardiovascular disease, unspecified|Cardiovascular disease, unspecified
C0018800|T033|AB|429.3|ICD9CM|Cardiomegaly|Cardiomegaly
C0018800|T033|PT|429.3|ICD9CM|Cardiomegaly|Cardiomegaly
C0016809|T046|PT|429.4|ICD9CM|Functional disturbances following cardiac surgery|Functional disturbances following cardiac surgery
C0016809|T046|AB|429.4|ICD9CM|Hrt dis postcardiac surg|Hrt dis postcardiac surg
C0155712|T046|AB|429.5|ICD9CM|Chordae tendinae rupture|Chordae tendinae rupture
C0155712|T046|PT|429.5|ICD9CM|Rupture of chordae tendineae|Rupture of chordae tendineae
C0155713|T046|AB|429.6|ICD9CM|Papillary muscle rupture|Papillary muscle rupture
C0155713|T046|PT|429.6|ICD9CM|Rupture of papillary muscle|Rupture of papillary muscle
C0302375|T047|HT|429.7|ICD9CM|Certain sequelae of myocardial infarction, not elsewhere classified|Certain sequelae of myocardial infarction, not elsewhere classified
C0376115|T047|AB|429.71|ICD9CM|Acq cardiac septl defect|Acq cardiac septl defect
C0376115|T047|PT|429.71|ICD9CM|Acquired cardiac septal defect|Acquired cardiac septal defect
C0302376|T047|PT|429.79|ICD9CM|Certain sequelae of myocardial infarction, not elsewhere classified, other|Certain sequelae of myocardial infarction, not elsewhere classified, other
C0302376|T047|AB|429.79|ICD9CM|Other sequelae of MI NEC|Other sequelae of MI NEC
C0155717|T047|HT|429.8|ICD9CM|Other ill-defined heart diseases|Other ill-defined heart diseases
C0155718|T047|PT|429.81|ICD9CM|Other disorders of papillary muscle|Other disorders of papillary muscle
C0155718|T047|AB|429.81|ICD9CM|Papillary muscle dis NEC|Papillary muscle dis NEC
C0242407|T047|AB|429.82|ICD9CM|Hyperkinetic heart dis|Hyperkinetic heart dis
C0242407|T047|PT|429.82|ICD9CM|Hyperkinetic heart disease|Hyperkinetic heart disease
C1739395|T047|PT|429.83|ICD9CM|Takotsubo syndrome|Takotsubo syndrome
C1739395|T047|AB|429.83|ICD9CM|Takotsubo syndrome|Takotsubo syndrome
C0155717|T047|AB|429.89|ICD9CM|Ill-defined hrt dis NEC|Ill-defined hrt dis NEC
C0155717|T047|PT|429.89|ICD9CM|Other ill-defined heart diseases|Other ill-defined heart diseases
C0018799|T047|AB|429.9|ICD9CM|Heart disease NOS|Heart disease NOS
C0018799|T047|PT|429.9|ICD9CM|Heart disease, unspecified|Heart disease, unspecified
C0038525|T047|AB|430|ICD9CM|Subarachnoid hemorrhage|Subarachnoid hemorrhage
C0038525|T047|PT|430|ICD9CM|Subarachnoid hemorrhage|Subarachnoid hemorrhage
C0007820|T047|HT|430-438.99|ICD9CM|CEREBROVASCULAR DISEASE|CEREBROVASCULAR DISEASE
C2937358|T046|AB|431|ICD9CM|Intracerebral hemorrhage|Intracerebral hemorrhage
C2937358|T046|PT|431|ICD9CM|Intracerebral hemorrhage|Intracerebral hemorrhage
C0155719|T046|HT|432|ICD9CM|Other and unspecified intracranial hemorrhage|Other and unspecified intracranial hemorrhage
C1318552|T047|AB|432.0|ICD9CM|Nontraum extradural hem|Nontraum extradural hem
C1318552|T047|PT|432.0|ICD9CM|Nontraumatic extradural hemorrhage|Nontraumatic extradural hemorrhage
C0018946|T046|AB|432.1|ICD9CM|Subdural hemorrhage|Subdural hemorrhage
C0018946|T046|PT|432.1|ICD9CM|Subdural hemorrhage|Subdural hemorrhage
C0151699|T046|AB|432.9|ICD9CM|Intracranial hemorr NOS|Intracranial hemorr NOS
C0151699|T046|PT|432.9|ICD9CM|Unspecified intracranial hemorrhage|Unspecified intracranial hemorrhage
C0155727|T047|HT|433|ICD9CM|Occlusion and stenosis of precerebral arteries|Occlusion and stenosis of precerebral arteries
C0265098|T190|HT|433.0|ICD9CM|Occlusion and stenosis of basilar artery|Occlusion and stenosis of basilar artery
C0375273|T047|PT|433.00|ICD9CM|Occlusion and stenosis of basilar artery without mention of cerebral infarction|Occlusion and stenosis of basilar artery without mention of cerebral infarction
C0375273|T047|AB|433.00|ICD9CM|Ocl bslr art wo infrct|Ocl bslr art wo infrct
C0375274|T047|PT|433.01|ICD9CM|Occlusion and stenosis of basilar artery with cerebral infarction|Occlusion and stenosis of basilar artery with cerebral infarction
C0375274|T047|AB|433.01|ICD9CM|Ocl bslr art w infrct|Ocl bslr art w infrct
C0600126|T046|HT|433.1|ICD9CM|Occlusion and stenosis of carotid artery|Occlusion and stenosis of carotid artery
C0375275|T047|PT|433.10|ICD9CM|Occlusion and stenosis of carotid artery without mention of cerebral infarction|Occlusion and stenosis of carotid artery without mention of cerebral infarction
C0375275|T047|AB|433.10|ICD9CM|Ocl crtd art wo infrct|Ocl crtd art wo infrct
C0375276|T047|PT|433.11|ICD9CM|Occlusion and stenosis of carotid artery with cerebral infarction|Occlusion and stenosis of carotid artery with cerebral infarction
C0375276|T047|AB|433.11|ICD9CM|Ocl crtd art w infrct|Ocl crtd art w infrct
C0155724|T046|HT|433.2|ICD9CM|Occlusion and stenosis of vertebral artery|Occlusion and stenosis of vertebral artery
C0375277|T047|PT|433.20|ICD9CM|Occlusion and stenosis of vertebral artery without mention of cerebral infarction|Occlusion and stenosis of vertebral artery without mention of cerebral infarction
C0375277|T047|AB|433.20|ICD9CM|Ocl vrtb art wo infrct|Ocl vrtb art wo infrct
C0375278|T047|PT|433.21|ICD9CM|Occlusion and stenosis of vertebral artery with cerebral infarction|Occlusion and stenosis of vertebral artery with cerebral infarction
C0375278|T047|AB|433.21|ICD9CM|Ocl vrtb art w infrct|Ocl vrtb art w infrct
C0155725|T047|HT|433.3|ICD9CM|Occlusion and stenosis of multiple and bilateral precerebral arteries|Occlusion and stenosis of multiple and bilateral precerebral arteries
C0375279|T047|AB|433.30|ICD9CM|Ocl mlt bi art wo infrct|Ocl mlt bi art wo infrct
C0375280|T047|PT|433.31|ICD9CM|Occlusion and stenosis of multiple and bilateral precerebral arteries with cerebral infarction|Occlusion and stenosis of multiple and bilateral precerebral arteries with cerebral infarction
C0375280|T047|AB|433.31|ICD9CM|Ocl mlt bi art w infrct|Ocl mlt bi art w infrct
C0155726|T047|HT|433.8|ICD9CM|Occlusion and stenosis of other specified precerebral artery|Occlusion and stenosis of other specified precerebral artery
C0375281|T047|PT|433.80|ICD9CM|Occlusion and stenosis of other specified precerebral artery without mention of cerebral infarction|Occlusion and stenosis of other specified precerebral artery without mention of cerebral infarction
C0375281|T047|AB|433.80|ICD9CM|Ocl spcf art wo infrct|Ocl spcf art wo infrct
C0375282|T047|PT|433.81|ICD9CM|Occlusion and stenosis of other specified precerebral artery with cerebral infarction|Occlusion and stenosis of other specified precerebral artery with cerebral infarction
C0375282|T047|AB|433.81|ICD9CM|Ocl spcf art w infrct|Ocl spcf art w infrct
C0155727|T047|HT|433.9|ICD9CM|Occlusion and stenosis of unspecified precerebral artery|Occlusion and stenosis of unspecified precerebral artery
C0375283|T047|PT|433.90|ICD9CM|Occlusion and stenosis of unspecified precerebral artery without mention of cerebral infarction|Occlusion and stenosis of unspecified precerebral artery without mention of cerebral infarction
C0375283|T047|AB|433.90|ICD9CM|Ocl art NOS wo infrct|Ocl art NOS wo infrct
C0375284|T047|PT|433.91|ICD9CM|Occlusion and stenosis of unspecified precerebral artery with cerebral infarction|Occlusion and stenosis of unspecified precerebral artery with cerebral infarction
C0375284|T047|AB|433.91|ICD9CM|Ocl art NOS w infrct|Ocl art NOS w infrct
C0028790|T020|HT|434|ICD9CM|Occlusion of cerebral arteries|Occlusion of cerebral arteries
C0079102|T047|HT|434.0|ICD9CM|Cerebral thrombosis|Cerebral thrombosis
C0375285|T047|PT|434.00|ICD9CM|Cerebral thrombosis without mention of cerebral infarction|Cerebral thrombosis without mention of cerebral infarction
C0375285|T047|AB|434.00|ICD9CM|Crbl thrmbs wo infrct|Crbl thrmbs wo infrct
C0375286|T047|PT|434.01|ICD9CM|Cerebral thrombosis with cerebral infarction|Cerebral thrombosis with cerebral infarction
C0375286|T047|AB|434.01|ICD9CM|Crbl thrmbs w infrct|Crbl thrmbs w infrct
C0007780|T047|HT|434.1|ICD9CM|Cerebral embolism|Cerebral embolism
C0375287|T047|PT|434.10|ICD9CM|Cerebral embolism without mention of cerebral infarction|Cerebral embolism without mention of cerebral infarction
C0375287|T047|AB|434.10|ICD9CM|Crbl emblsm wo infrct|Crbl emblsm wo infrct
C0375288|T047|PT|434.11|ICD9CM|Cerebral embolism with cerebral infarction|Cerebral embolism with cerebral infarction
C0375288|T047|AB|434.11|ICD9CM|Crbl emblsm w infrct|Crbl emblsm w infrct
C0028790|T020|HT|434.9|ICD9CM|Cerebral artery occlusion, unspecified|Cerebral artery occlusion, unspecified
C0375290|T047|PT|434.90|ICD9CM|Cerebral artery occlusion, unspecified without mention of cerebral infarction|Cerebral artery occlusion, unspecified without mention of cerebral infarction
C0375290|T047|AB|434.90|ICD9CM|Crbl art oc NOS wo infrc|Crbl art oc NOS wo infrc
C0375291|T047|PT|434.91|ICD9CM|Cerebral artery occlusion, unspecified with cerebral infarction|Cerebral artery occlusion, unspecified with cerebral infarction
C0375291|T047|AB|434.91|ICD9CM|Crbl art ocl NOS w infrc|Crbl art ocl NOS w infrc
C0917805|T047|HT|435|ICD9CM|Transient cerebral ischemia|Transient cerebral ischemia
C0004812|T047|AB|435.0|ICD9CM|Basilar artery syndrome|Basilar artery syndrome
C0004812|T047|PT|435.0|ICD9CM|Basilar artery syndrome|Basilar artery syndrome
C2931914|T047|AB|435.1|ICD9CM|Vertebral artery syndrom|Vertebral artery syndrom
C2931914|T047|PT|435.1|ICD9CM|Vertebral artery syndrome|Vertebral artery syndrome
C0038531|T047|AB|435.2|ICD9CM|Subclavian steal syndrom|Subclavian steal syndrom
C0038531|T047|PT|435.2|ICD9CM|Subclavian steal syndrome|Subclavian steal syndrome
C0042568|T047|AB|435.3|ICD9CM|Vertbrobaslr artery synd|Vertbrobaslr artery synd
C0042568|T047|PT|435.3|ICD9CM|Vertebrobasilar artery syndrome|Vertebrobasilar artery syndrome
C0155728|T047|PT|435.8|ICD9CM|Other specified transient cerebral ischemias|Other specified transient cerebral ischemias
C0155728|T047|AB|435.8|ICD9CM|Trans cereb ischemia NEC|Trans cereb ischemia NEC
C0917805|T047|AB|435.9|ICD9CM|Trans cereb ischemia NOS|Trans cereb ischemia NOS
C0917805|T047|PT|435.9|ICD9CM|Unspecified transient cerebral ischemia|Unspecified transient cerebral ischemia
C0001365|T047|PT|436|ICD9CM|Acute, but ill-defined, cerebrovascular disease|Acute, but ill-defined, cerebrovascular disease
C0001365|T047|AB|436|ICD9CM|Cva|Cva
C0155729|T047|HT|437|ICD9CM|Other and ill-defined cerebrovascular disease|Other and ill-defined cerebrovascular disease
C0007775|T047|AB|437.0|ICD9CM|Cerebral atherosclerosis|Cerebral atherosclerosis
C0007775|T047|PT|437.0|ICD9CM|Cerebral atherosclerosis|Cerebral atherosclerosis
C0029626|T047|AB|437.1|ICD9CM|Ac cerebrovasc insuf NOS|Ac cerebrovasc insuf NOS
C0029626|T047|PT|437.1|ICD9CM|Other generalized ischemic cerebrovascular disease|Other generalized ischemic cerebrovascular disease
C0151620|T047|AB|437.2|ICD9CM|Hypertens encephalopathy|Hypertens encephalopathy
C0151620|T047|PT|437.2|ICD9CM|Hypertensive encephalopathy|Hypertensive encephalopathy
C0155730|T190|PT|437.3|ICD9CM|Cerebral aneurysm, nonruptured|Cerebral aneurysm, nonruptured
C0155730|T190|AB|437.3|ICD9CM|Nonrupt cerebral aneurym|Nonrupt cerebral aneurym
C0007773|T047|AB|437.4|ICD9CM|Cerebral arteritis|Cerebral arteritis
C0007773|T047|PT|437.4|ICD9CM|Cerebral arteritis|Cerebral arteritis
C0026654|T047|AB|437.5|ICD9CM|Moyamoya disease|Moyamoya disease
C0026654|T047|PT|437.5|ICD9CM|Moyamoya disease|Moyamoya disease
C0155731|T047|AB|437.6|ICD9CM|Nonpyogen thrombos sinus|Nonpyogen thrombos sinus
C0155731|T047|PT|437.6|ICD9CM|Nonpyogenic thrombosis of intracranial venous sinus|Nonpyogenic thrombosis of intracranial venous sinus
C0338591|T048|AB|437.7|ICD9CM|Transient global amnesia|Transient global amnesia
C0338591|T048|PT|437.7|ICD9CM|Transient global amnesia|Transient global amnesia
C0155729|T047|AB|437.8|ICD9CM|Cerebrovasc disease NEC|Cerebrovasc disease NEC
C0155729|T047|PT|437.8|ICD9CM|Other ill-defined cerebrovascular disease|Other ill-defined cerebrovascular disease
C0007820|T047|AB|437.9|ICD9CM|Cerebrovasc disease NOS|Cerebrovasc disease NOS
C0007820|T047|PT|437.9|ICD9CM|Unspecified cerebrovascular disease|Unspecified cerebrovascular disease
C0155732|T046|HT|438|ICD9CM|Late effects of cerebrovascular disease|Late effects of cerebrovascular disease
C0489983|T046|AB|438.0|ICD9CM|Late ef CV dis-cognf def|Late ef CV dis-cognf def
C0489983|T046|PT|438.0|ICD9CM|Late effects of cerebrovascular disease, cognitive deficits|Late effects of cerebrovascular disease, cognitive deficits
C0489984|T046|HT|438.1|ICD9CM|Speech and language deficits as late effect of cerebrovascular disease|Speech and language deficits as late effect of cerebrovascular disease
C0489984|T046|AB|438.10|ICD9CM|Late ef-spch/lng def NOS|Late ef-spch/lng def NOS
C0489984|T046|PT|438.10|ICD9CM|Late effects of cerebrovascular disease, speech and language deficit, unspecified|Late effects of cerebrovascular disease, speech and language deficit, unspecified
C0489985|T046|AB|438.11|ICD9CM|Late eff CV dis-aphasia|Late eff CV dis-aphasia
C0489985|T046|PT|438.11|ICD9CM|Late effects of cerebrovascular disease, aphasia|Late effects of cerebrovascular disease, aphasia
C0489986|T046|AB|438.12|ICD9CM|Late eff CV dis-dysphsia|Late eff CV dis-dysphsia
C0489986|T046|PT|438.12|ICD9CM|Late effects of cerebrovascular disease, dysphasia|Late effects of cerebrovascular disease, dysphasia
C0013362|T048|AB|438.13|ICD9CM|Late eff CV-dysarthria|Late eff CV-dysarthria
C0013362|T048|PT|438.13|ICD9CM|Late effects of cerebrovascular disease, dysarthria|Late effects of cerebrovascular disease, dysarthria
C0454533|T047|AB|438.14|ICD9CM|Late eff CV-fluency dis|Late eff CV-fluency dis
C0454533|T047|PT|438.14|ICD9CM|Late effects of cerebrovascular disease, fluency disorder|Late effects of cerebrovascular disease, fluency disorder
C0489987|T047|AB|438.19|ICD9CM|Late ef-spch/lang df NEC|Late ef-spch/lang df NEC
C0489987|T047|PT|438.19|ICD9CM|Late effects of cerebrovascular disease, other speech and language deficits|Late effects of cerebrovascular disease, other speech and language deficits
C0489988|T047|HT|438.2|ICD9CM|Hemiplegia/hemiparesis as late effect of cerebrovascular disease|Hemiplegia/hemiparesis as late effect of cerebrovascular disease
C0489989|T047|AB|438.20|ICD9CM|Late ef-hemplga side NOS|Late ef-hemplga side NOS
C0489989|T047|PT|438.20|ICD9CM|Late effects of cerebrovascular disease, hemiplegia affecting unspecified side|Late effects of cerebrovascular disease, hemiplegia affecting unspecified side
C0489990|T046|AB|438.21|ICD9CM|Late ef-hemplga dom side|Late ef-hemplga dom side
C0489990|T046|PT|438.21|ICD9CM|Late effects of cerebrovascular disease, hemiplegia affecting dominant side|Late effects of cerebrovascular disease, hemiplegia affecting dominant side
C0489991|T046|AB|438.22|ICD9CM|Late ef-hemiplga non-dom|Late ef-hemiplga non-dom
C0489991|T046|PT|438.22|ICD9CM|Late effects of cerebrovascular disease, hemiplegia affecting nondominant side|Late effects of cerebrovascular disease, hemiplegia affecting nondominant side
C0489992|T046|HT|438.3|ICD9CM|Monoplegia of upper limb as late effect of cerebrovascular disease|Monoplegia of upper limb as late effect of cerebrovascular disease
C0489993|T047|AB|438.30|ICD9CM|Late ef-mplga up lmb NOS|Late ef-mplga up lmb NOS
C0489993|T047|PT|438.30|ICD9CM|Late effects of cerebrovascular disease, monoplegia of upper limb affecting unspecified side|Late effects of cerebrovascular disease, monoplegia of upper limb affecting unspecified side
C0489994|T046|AB|438.31|ICD9CM|Late ef-mplga up lmb dom|Late ef-mplga up lmb dom
C0489994|T046|PT|438.31|ICD9CM|Late effects of cerebrovascular disease, monoplegia of upper limb affecting dominant side|Late effects of cerebrovascular disease, monoplegia of upper limb affecting dominant side
C0489995|T046|PT|438.32|ICD9CM|Late effects of cerebrovascular disease, monoplegia of upper limb affecting nondominant side|Late effects of cerebrovascular disease, monoplegia of upper limb affecting nondominant side
C0489995|T046|AB|438.32|ICD9CM|Lt ef-mplga uplmb nondom|Lt ef-mplga uplmb nondom
C0489996|T046|HT|438.4|ICD9CM|Monoplegia of lower limb as late effect of cerebrovascular disease|Monoplegia of lower limb as late effect of cerebrovascular disease
C0489997|T047|PT|438.40|ICD9CM|Late effects of cerebrovascular disease, monoplegia of lower limb affecting unspecified side|Late effects of cerebrovascular disease, monoplegia of lower limb affecting unspecified side
C0489997|T047|AB|438.40|ICD9CM|Lte ef-mplga low lmb NOS|Lte ef-mplga low lmb NOS
C0489998|T046|PT|438.41|ICD9CM|Late effects of cerebrovascular disease, monoplegia of lower limb affecting dominant side|Late effects of cerebrovascular disease, monoplegia of lower limb affecting dominant side
C0489998|T046|AB|438.41|ICD9CM|Lte ef-mplga low lmb dom|Lte ef-mplga low lmb dom
C0489999|T046|PT|438.42|ICD9CM|Late effects of cerebrovascular disease, monoplegia of lower limb affecting nondominant side|Late effects of cerebrovascular disease, monoplegia of lower limb affecting nondominant side
C0489999|T046|AB|438.42|ICD9CM|Lt ef-mplga lowlmb nondm|Lt ef-mplga lowlmb nondm
C0490000|T047|HT|438.5|ICD9CM|Other paralytic syndrome as late effect of cerebrovascular disease|Other paralytic syndrome as late effect of cerebrovascular disease
C0490001|T047|PT|438.50|ICD9CM|Late effects of cerebrovascular disease, other paralytic syndrome affecting unspecified side|Late effects of cerebrovascular disease, other paralytic syndrome affecting unspecified side
C0490001|T047|AB|438.50|ICD9CM|Lt ef oth paral side NOS|Lt ef oth paral side NOS
C0490002|T047|PT|438.51|ICD9CM|Late effects of cerebrovascular disease, other paralytic syndrome affecting dominant side|Late effects of cerebrovascular disease, other paralytic syndrome affecting dominant side
C0490002|T047|AB|438.51|ICD9CM|Lt ef oth paral dom side|Lt ef oth paral dom side
C0490003|T047|PT|438.52|ICD9CM|Late effects of cerebrovascular disease, other paralytic syndrome affecting nondominant side|Late effects of cerebrovascular disease, other paralytic syndrome affecting nondominant side
C0490003|T047|AB|438.52|ICD9CM|Lt ef oth parals non-dom|Lt ef oth parals non-dom
C0695232|T047|PT|438.53|ICD9CM|Late effects of cerebrovascular disease, other paralytic syndrome, bilateral|Late effects of cerebrovascular disease, other paralytic syndrome, bilateral
C0695232|T047|AB|438.53|ICD9CM|Lt ef oth parals-bilat|Lt ef oth parals-bilat
C1135206|T046|AB|438.6|ICD9CM|Alteration of sensations|Alteration of sensations
C1135206|T046|PT|438.6|ICD9CM|Late effects of cerebrovascular disease, alterations of sensations|Late effects of cerebrovascular disease, alterations of sensations
C3665387|T046|AB|438.7|ICD9CM|Disturbances of vision|Disturbances of vision
C3665387|T046|PT|438.7|ICD9CM|Late effects of cerebrovascular disease, disturbances of vision|Late effects of cerebrovascular disease, disturbances of vision
C0490004|T046|HT|438.8|ICD9CM|Other late effects of cerebrovascular disease|Other late effects of cerebrovascular disease
C0490005|T046|AB|438.81|ICD9CM|Late eff CV dis-apraxia|Late eff CV dis-apraxia
C0490005|T046|PT|438.81|ICD9CM|Other late effects of cerebrovascular disease, apraxia|Other late effects of cerebrovascular disease, apraxia
C0490006|T046|AB|438.82|ICD9CM|Late ef CV dis dysphagia|Late ef CV dis dysphagia
C0490006|T046|PT|438.82|ICD9CM|Other late effects of cerebrovascular disease, dysphagia|Other late effects of cerebrovascular disease, dysphagia
C0427055|T047|AB|438.83|ICD9CM|Facial weakness|Facial weakness
C0427055|T047|PT|438.83|ICD9CM|Other late effects of cerebrovascular disease, facial weakness|Other late effects of cerebrovascular disease, facial weakness
C1135207|T046|AB|438.84|ICD9CM|Ataxia|Ataxia
C1135207|T046|PT|438.84|ICD9CM|Other late effects of cerebrovascular disease, ataxia|Other late effects of cerebrovascular disease, ataxia
C1135208|T047|PT|438.85|ICD9CM|Other late effects of cerebrovascular disease, vertigo|Other late effects of cerebrovascular disease, vertigo
C1135208|T047|AB|438.85|ICD9CM|Vertigo|Vertigo
C0490004|T046|AB|438.89|ICD9CM|Late effect CV dis NEC|Late effect CV dis NEC
C0490004|T046|PT|438.89|ICD9CM|Other late effects of cerebrovascular disease|Other late effects of cerebrovascular disease
C0155732|T046|AB|438.9|ICD9CM|Late effect CV dis NOS|Late effect CV dis NOS
C0155732|T046|PT|438.9|ICD9CM|Unspecified late effects of cerebrovascular disease|Unspecified late effects of cerebrovascular disease
C0004153|T047|HT|440|ICD9CM|Atherosclerosis|Atherosclerosis
C0178274|T047|HT|440-449.99|ICD9CM|DISEASES OF ARTERIES, ARTERIOLES, AND CAPILLARIES|DISEASES OF ARTERIES, ARTERIOLES, AND CAPILLARIES
C0155733|T047|AB|440.0|ICD9CM|Aortic atherosclerosis|Aortic atherosclerosis
C0155733|T047|PT|440.0|ICD9CM|Atherosclerosis of aorta|Atherosclerosis of aorta
C0155734|T047|PT|440.1|ICD9CM|Atherosclerosis of renal artery|Atherosclerosis of renal artery
C0155734|T047|AB|440.1|ICD9CM|Renal artery atheroscler|Renal artery atheroscler
C3495604|T047|HT|440.2|ICD9CM|Atherosclerosis of native arteries of the extremities|Atherosclerosis of native arteries of the extremities
C0375294|T047|PT|440.20|ICD9CM|Atherosclerosis of native arteries of the extremities, unspecified|Atherosclerosis of native arteries of the extremities, unspecified
C0375294|T047|AB|440.20|ICD9CM|Athscl extrm ntv art NOS|Athscl extrm ntv art NOS
C0375295|T047|AB|440.21|ICD9CM|Ath ext ntv at w claudct|Ath ext ntv at w claudct
C0375295|T047|PT|440.21|ICD9CM|Atherosclerosis of native arteries of the extremities with intermittent claudication|Atherosclerosis of native arteries of the extremities with intermittent claudication
C2882703|T047|AB|440.22|ICD9CM|Ath ext ntv at w rst pn|Ath ext ntv at w rst pn
C2882703|T047|PT|440.22|ICD9CM|Atherosclerosis of native arteries of the extremities with rest pain|Atherosclerosis of native arteries of the extremities with rest pain
C0375297|T047|AB|440.23|ICD9CM|Ath ext ntv art ulcrtion|Ath ext ntv art ulcrtion
C0375297|T047|PT|440.23|ICD9CM|Atherosclerosis of native arteries of the extremities with ulceration|Atherosclerosis of native arteries of the extremities with ulceration
C0375298|T047|AB|440.24|ICD9CM|Ath ext ntv art gngrene|Ath ext ntv art gngrene
C0375298|T047|PT|440.24|ICD9CM|Atherosclerosis of native arteries of the extremities with gangrene|Atherosclerosis of native arteries of the extremities with gangrene
C0375299|T047|AB|440.29|ICD9CM|Athrsc extrm ntv art oth|Athrsc extrm ntv art oth
C0375299|T047|PT|440.29|ICD9CM|Other atherosclerosis of native arteries of the extremities|Other atherosclerosis of native arteries of the extremities
C0375300|T047|HT|440.3|ICD9CM|Of bypass graft of the extremities|Of bypass graft of the extremities
C0375301|T047|PT|440.30|ICD9CM|Atherosclerosis of unspecified bypass graft of the extremities|Atherosclerosis of unspecified bypass graft of the extremities
C0375301|T047|AB|440.30|ICD9CM|Athscl extrm bps gft NOS|Athscl extrm bps gft NOS
C0375302|T047|AB|440.31|ICD9CM|Ath ext autologs bps gft|Ath ext autologs bps gft
C0375302|T047|PT|440.31|ICD9CM|Atherosclerosis of autologous vein bypass graft of the extremities|Atherosclerosis of autologous vein bypass graft of the extremities
C1112691|T047|AB|440.32|ICD9CM|Ath ext nonautlg bps gft|Ath ext nonautlg bps gft
C1112691|T047|PT|440.32|ICD9CM|Atherosclerosis of nonautologous biological bypass graft of the extremities|Atherosclerosis of nonautologous biological bypass graft of the extremities
C1955783|T047|AB|440.4|ICD9CM|Chr tot occl art extrem|Chr tot occl art extrem
C1955783|T047|PT|440.4|ICD9CM|Chronic total occlusion of artery of the extremities|Chronic total occlusion of artery of the extremities
C0004155|T047|AB|440.8|ICD9CM|Atherosclerosis NEC|Atherosclerosis NEC
C0004155|T047|PT|440.8|ICD9CM|Atherosclerosis of other specified arteries|Atherosclerosis of other specified arteries
C0017327|T047|AB|440.9|ICD9CM|Atherosclerosis NOS|Atherosclerosis NOS
C0017327|T047|PT|440.9|ICD9CM|Generalized and unspecified atherosclerosis|Generalized and unspecified atherosclerosis
C1812607|T047|HT|441|ICD9CM|Aortic aneurysm and dissection|Aortic aneurysm and dissection
C0012736|T047|HT|441.0|ICD9CM|Dissecting aneurysm of aorta|Dissecting aneurysm of aorta
C0340643|T047|PT|441.00|ICD9CM|Dissection of aorta, unspecified site|Dissection of aorta, unspecified site
C0340643|T047|AB|441.00|ICD9CM|Dsct of aorta unsp site|Dsct of aorta unsp site
C0729233|T047|PT|441.01|ICD9CM|Dissection of aorta, thoracic|Dissection of aorta, thoracic
C0729233|T047|AB|441.01|ICD9CM|Dsct of thoracic aorta|Dsct of thoracic aorta
C0302465|T047|PT|441.02|ICD9CM|Dissection of aorta, abdominal|Dissection of aorta, abdominal
C0302465|T047|AB|441.02|ICD9CM|Dsct of abdominal aorta|Dsct of abdominal aorta
C0375305|T047|PT|441.03|ICD9CM|Dissection of aorta, thoracoabdominal|Dissection of aorta, thoracoabdominal
C0375305|T047|AB|441.03|ICD9CM|Dsct of thoracoabd aorta|Dsct of thoracoabd aorta
C0265010|T047|AB|441.1|ICD9CM|Ruptur thoracic aneurysm|Ruptur thoracic aneurysm
C0265010|T047|PT|441.1|ICD9CM|Thoracic aneurysm, ruptured|Thoracic aneurysm, ruptured
C3251816|T020|PT|441.2|ICD9CM|Thoracic aneurysm without mention of rupture|Thoracic aneurysm without mention of rupture
C3251816|T020|AB|441.2|ICD9CM|Thoracic aortic aneurysm|Thoracic aortic aneurysm
C0265012|T047|PT|441.3|ICD9CM|Abdominal aneurysm, ruptured|Abdominal aneurysm, ruptured
C0265012|T047|AB|441.3|ICD9CM|Rupt abd aortic aneurysm|Rupt abd aortic aneurysm
C0265011|T020|AB|441.4|ICD9CM|Abdom aortic aneurysm|Abdom aortic aneurysm
C0265011|T020|PT|441.4|ICD9CM|Abdominal aneurysm without mention of rupture|Abdominal aneurysm without mention of rupture
C0741160|T047|PT|441.5|ICD9CM|Aortic aneurysm of unspecified site, ruptured|Aortic aneurysm of unspecified site, ruptured
C0741160|T047|AB|441.5|ICD9CM|Rupt aortic aneurysm NOS|Rupt aortic aneurysm NOS
C1305122|T047|AB|441.6|ICD9CM|Thoracoabd aneurysm rupt|Thoracoabd aneurysm rupt
C1305122|T047|PT|441.6|ICD9CM|Thoracoabdominal aneurysm, ruptured|Thoracoabdominal aneurysm, ruptured
C0375306|T020|PT|441.7|ICD9CM|Thoracoabdominal aneurysm, without mention of rupture|Thoracoabdominal aneurysm, without mention of rupture
C0375306|T020|AB|441.7|ICD9CM|Thracabd anurysm wo rupt|Thracabd anurysm wo rupt
C0340629|T047|AB|441.9|ICD9CM|Aortic aneurysm NOS|Aortic aneurysm NOS
C0340629|T047|PT|441.9|ICD9CM|Aortic aneurysm of unspecified site without mention of rupture|Aortic aneurysm of unspecified site without mention of rupture
C0155740|T190|HT|442|ICD9CM|Other aneurysm|Other aneurysm
C0155741|T190|PT|442.0|ICD9CM|Aneurysm of artery of upper extremity|Aneurysm of artery of upper extremity
C0155741|T190|AB|442.0|ICD9CM|Upper extremity aneurysm|Upper extremity aneurysm
C0155742|T190|PT|442.1|ICD9CM|Aneurysm of renal artery|Aneurysm of renal artery
C0155742|T190|AB|442.1|ICD9CM|Renal artery aneurysm|Renal artery aneurysm
C0162870|T190|PT|442.2|ICD9CM|Aneurysm of iliac artery|Aneurysm of iliac artery
C0162870|T190|AB|442.2|ICD9CM|Iliac artery aneurysm|Iliac artery aneurysm
C0155744|T190|PT|442.3|ICD9CM|Aneurysm of artery of lower extremity|Aneurysm of artery of lower extremity
C0155744|T190|AB|442.3|ICD9CM|Lower extremity aneurysm|Lower extremity aneurysm
C0002945|T190|HT|442.8|ICD9CM|Aneurysm of other specified artery|Aneurysm of other specified artery
C0155745|T190|PT|442.81|ICD9CM|Aneurysm of artery of neck|Aneurysm of artery of neck
C0155745|T190|AB|442.81|ICD9CM|Aneurysm of neck|Aneurysm of neck
C0155746|T047|PT|442.82|ICD9CM|Aneurysm of subclavian artery|Aneurysm of subclavian artery
C0155746|T047|AB|442.82|ICD9CM|Subclavian aneurysm|Subclavian aneurysm
C0155747|T047|PT|442.83|ICD9CM|Aneurysm of splenic artery|Aneurysm of splenic artery
C0155747|T047|AB|442.83|ICD9CM|Splenic artery aneurysm|Splenic artery aneurysm
C0155748|T020|PT|442.84|ICD9CM|Aneurysm of other visceral artery|Aneurysm of other visceral artery
C0155748|T020|AB|442.84|ICD9CM|Visceral aneurysm NEC|Visceral aneurysm NEC
C0002946|T033|AB|442.89|ICD9CM|Aneurysm NEC|Aneurysm NEC
C0002946|T033|PT|442.89|ICD9CM|Aneurysm of other specified artery|Aneurysm of other specified artery
C0002940|T046|AB|442.9|ICD9CM|Aneurysm NOS|Aneurysm NOS
C0002940|T046|PT|442.9|ICD9CM|Aneurysm of unspecified site|Aneurysm of unspecified site
C0553983|T047|HT|443|ICD9CM|Other peripheral vascular disease|Other peripheral vascular disease
C0034735|T047|AB|443.0|ICD9CM|Raynaud's syndrome|Raynaud's syndrome
C0034735|T047|PT|443.0|ICD9CM|Raynaud's syndrome|Raynaud's syndrome
C0040021|T047|AB|443.1|ICD9CM|Thromboangiit obliterans|Thromboangiit obliterans
C0040021|T047|PT|443.1|ICD9CM|Thromboangiitis obliterans [Buerger's disease]|Thromboangiitis obliterans [Buerger's disease]
C1135209|T047|HT|443.2|ICD9CM|Other arterial dissection|Other arterial dissection
C0338585|T047|AB|443.21|ICD9CM|Dissect carotid artery|Dissect carotid artery
C0338585|T047|PT|443.21|ICD9CM|Dissection of carotid artery|Dissection of carotid artery
C0340649|T047|AB|443.22|ICD9CM|Dissection iliac artery|Dissection iliac artery
C0340649|T047|PT|443.22|ICD9CM|Dissection of iliac artery|Dissection of iliac artery
C0919563|T047|PT|443.23|ICD9CM|Dissection of renal artery|Dissection of renal artery
C0919563|T047|AB|443.23|ICD9CM|Dissection renal artery|Dissection renal artery
C0338586|T047|AB|443.24|ICD9CM|Dissect vertebral artery|Dissect vertebral artery
C0338586|T047|PT|443.24|ICD9CM|Dissection of vertebral artery|Dissection of vertebral artery
C1135210|T047|AB|443.29|ICD9CM|Dissection artery NEC|Dissection artery NEC
C1135210|T047|PT|443.29|ICD9CM|Dissection of other artery|Dissection of other artery
C0029822|T047|HT|443.8|ICD9CM|Other specified peripheral vascular diseases|Other specified peripheral vascular diseases
C0031115|T047|AB|443.81|ICD9CM|Angiopathy in other dis|Angiopathy in other dis
C0031115|T047|PT|443.81|ICD9CM|Peripheral angiopathy in diseases classified elsewhere|Peripheral angiopathy in diseases classified elsewhere
C0014804|T047|AB|443.82|ICD9CM|Erythromelalgia|Erythromelalgia
C0014804|T047|PT|443.82|ICD9CM|Erythromelalgia|Erythromelalgia
C0553983|T047|PT|443.89|ICD9CM|Other specified peripheral vascular diseases|Other specified peripheral vascular diseases
C0553983|T047|AB|443.89|ICD9CM|Periph vascular dis NEC|Periph vascular dis NEC
C0085096|T047|AB|443.9|ICD9CM|Periph vascular dis NOS|Periph vascular dis NOS
C0085096|T047|PT|443.9|ICD9CM|Peripheral vascular disease, unspecified|Peripheral vascular disease, unspecified
C0155749|T046|HT|444|ICD9CM|Arterial embolism and thrombosis|Arterial embolism and thrombosis
C0013923|T046|HT|444.0|ICD9CM|Embolism and thrombosis of abdominal aorta|Embolism and thrombosis of abdominal aorta
C0023370|T047|AB|444.01|ICD9CM|Saddle embolus abd aorta|Saddle embolus abd aorta
C0023370|T047|PT|444.01|ICD9CM|Saddle embolus of abdominal aorta|Saddle embolus of abdominal aorta
C3161092|T047|AB|444.09|ICD9CM|Ot art emb/thrm abd aort|Ot art emb/thrm abd aort
C3161092|T047|PT|444.09|ICD9CM|Other arterial embolism and thrombosis of abdominal aorta|Other arterial embolism and thrombosis of abdominal aorta
C0155750|T046|PT|444.1|ICD9CM|Embolism and thrombosis of thoracic aorta|Embolism and thrombosis of thoracic aorta
C0155750|T046|AB|444.1|ICD9CM|Thoracic aortic embolism|Thoracic aortic embolism
C0340579|T046|HT|444.2|ICD9CM|Embolism and thrombosis of arteries of the extremities|Embolism and thrombosis of arteries of the extremities
C0494620|T046|PT|444.21|ICD9CM|Arterial embolism and thrombosis of upper extremity|Arterial embolism and thrombosis of upper extremity
C0494620|T046|AB|444.21|ICD9CM|Upper extremity embolism|Upper extremity embolism
C0340589|T046|PT|444.22|ICD9CM|Arterial embolism and thrombosis of lower extremity|Arterial embolism and thrombosis of lower extremity
C0340589|T046|AB|444.22|ICD9CM|Lower extremity embolism|Lower extremity embolism
C0155754|T047|HT|444.8|ICD9CM|Embolism and thrombosis of other specified artery|Embolism and thrombosis of other specified artery
C0155755|T046|PT|444.81|ICD9CM|Embolism and thrombosis of iliac artery|Embolism and thrombosis of iliac artery
C0155755|T046|AB|444.81|ICD9CM|Iliac artery embolism|Iliac artery embolism
C0348650|T047|AB|444.89|ICD9CM|Arterial embolism NEC|Arterial embolism NEC
C0348650|T047|PT|444.89|ICD9CM|Embolism and thrombosis of other specified artery|Embolism and thrombosis of other specified artery
C0013924|T046|AB|444.9|ICD9CM|Arterial embolism NOS|Arterial embolism NOS
C0013924|T046|PT|444.9|ICD9CM|Embolism and thrombosis of unspecified artery|Embolism and thrombosis of unspecified artery
C0149649|T047|HT|445|ICD9CM|Atheroembolism|Atheroembolism
C1135211|T047|HT|445.0|ICD9CM|Atheroembolism Of extremities|Atheroembolism Of extremities
C1135212|T047|PT|445.01|ICD9CM|Atheroembolism of upper extremity|Atheroembolism of upper extremity
C1135212|T047|AB|445.01|ICD9CM|Atheroembolism,upper ext|Atheroembolism,upper ext
C1135213|T047|PT|445.02|ICD9CM|Atheroembolism of lower extremity|Atheroembolism of lower extremity
C1135213|T047|AB|445.02|ICD9CM|Atheroembolism,lower ext|Atheroembolism,lower ext
C1135216|T047|HT|445.8|ICD9CM|Atheroembolism of other sites|Atheroembolism of other sites
C0268792|T047|PT|445.81|ICD9CM|Atheroembolism of kidney|Atheroembolism of kidney
C0268792|T047|AB|445.81|ICD9CM|Atheroembolism, kidney|Atheroembolism, kidney
C1135216|T047|PT|445.89|ICD9CM|Atheroembolism of other site|Atheroembolism of other site
C1135216|T047|AB|445.89|ICD9CM|Atheroembolism, site NEC|Atheroembolism, site NEC
C0155757|T047|HT|446|ICD9CM|Polyarteritis nodosa and allied conditions|Polyarteritis nodosa and allied conditions
C0031036|T047|AB|446.0|ICD9CM|Polyarteritis nodosa|Polyarteritis nodosa
C0031036|T047|PT|446.0|ICD9CM|Polyarteritis nodosa|Polyarteritis nodosa
C0026691|T047|PT|446.1|ICD9CM|Acute febrile mucocutaneous lymph node syndrome [MCLS]|Acute febrile mucocutaneous lymph node syndrome [MCLS]
C0026691|T047|AB|446.1|ICD9CM|Mucocutan lymph node syn|Mucocutan lymph node syn
C0151436|T047|HT|446.2|ICD9CM|Hypersensitivity angiitis|Hypersensitivity angiitis
C0151436|T047|AB|446.20|ICD9CM|Hypersensit angiitis NOS|Hypersensit angiitis NOS
C0151436|T047|PT|446.20|ICD9CM|Hypersensitivity angiitis, unspecified|Hypersensitivity angiitis, unspecified
C0403529|T047|AB|446.21|ICD9CM|Goodpasture's syndrome|Goodpasture's syndrome
C0403529|T047|PT|446.21|ICD9CM|Goodpasture's syndrome|Goodpasture's syndrome
C0155758|T047|AB|446.29|ICD9CM|Hypersensit angiitis NEC|Hypersensit angiitis NEC
C0155758|T047|PT|446.29|ICD9CM|Other specified hypersensitivity angiitis|Other specified hypersensitivity angiitis
C0018197|T191|AB|446.3|ICD9CM|Lethal midline granuloma|Lethal midline granuloma
C0018197|T191|PT|446.3|ICD9CM|Lethal midline granuloma|Lethal midline granuloma
C3495801|T047|AB|446.4|ICD9CM|Wegener's granulomatosis|Wegener's granulomatosis
C3495801|T047|PT|446.4|ICD9CM|Wegener's granulomatosis|Wegener's granulomatosis
C0039483|T047|AB|446.5|ICD9CM|Giant cell arteritis|Giant cell arteritis
C0039483|T047|PT|446.5|ICD9CM|Giant cell arteritis|Giant cell arteritis
C2717961|T047|AB|446.6|ICD9CM|Thrombot microangiopathy|Thrombot microangiopathy
C2717961|T047|PT|446.6|ICD9CM|Thrombotic microangiopathy|Thrombotic microangiopathy
C0039263|T047|AB|446.7|ICD9CM|Takayasu's disease|Takayasu's disease
C0039263|T047|PT|446.7|ICD9CM|Takayasu's disease|Takayasu's disease
C0155759|T047|HT|447|ICD9CM|Other disorders of arteries and arterioles|Other disorders of arteries and arterioles
C1541850|T020|AB|447.0|ICD9CM|Acq arterioven fistula|Acq arterioven fistula
C1541850|T020|PT|447.0|ICD9CM|Arteriovenous fistula, acquired|Arteriovenous fistula, acquired
C0038449|T046|AB|447.1|ICD9CM|Stricture of artery|Stricture of artery
C0038449|T046|PT|447.1|ICD9CM|Stricture of artery|Stricture of artery
C0155760|T047|AB|447.2|ICD9CM|Rupture of artery|Rupture of artery
C0155760|T047|PT|447.2|ICD9CM|Rupture of artery|Rupture of artery
C0155761|T047|PT|447.3|ICD9CM|Hyperplasia of renal artery|Hyperplasia of renal artery
C0155761|T047|AB|447.3|ICD9CM|Renal artery hyperplasia|Renal artery hyperplasia
C1861783|T047|AB|447.4|ICD9CM|Celiac art compress syn|Celiac art compress syn
C1861783|T047|PT|447.4|ICD9CM|Celiac artery compression syndrome|Celiac artery compression syndrome
C0155762|T047|AB|447.5|ICD9CM|Necrosis of artery|Necrosis of artery
C0155762|T047|PT|447.5|ICD9CM|Necrosis of artery|Necrosis of artery
C0003860|T046|AB|447.6|ICD9CM|Arteritis NOS|Arteritis NOS
C0003860|T046|PT|447.6|ICD9CM|Arteritis, unspecified|Arteritis, unspecified
C0265004|T047|HT|447.7|ICD9CM|Aortic ectasia|Aortic ectasia
C2921068|T047|AB|447.70|ICD9CM|Aortic ectasia, site NOS|Aortic ectasia, site NOS
C2921068|T047|PT|447.70|ICD9CM|Aortic ectasia, unspecified site|Aortic ectasia, unspecified site
C2921069|T047|AB|447.71|ICD9CM|Thoracic aortic ectasia|Thoracic aortic ectasia
C2921069|T047|PT|447.71|ICD9CM|Thoracic aortic ectasia|Thoracic aortic ectasia
C2921070|T047|AB|447.72|ICD9CM|Abdominal aortic ectasia|Abdominal aortic ectasia
C2921070|T047|PT|447.72|ICD9CM|Abdominal aortic ectasia|Abdominal aortic ectasia
C2921071|T047|AB|447.73|ICD9CM|Thoracoabd aortc ectasia|Thoracoabd aortc ectasia
C2921071|T047|PT|447.73|ICD9CM|Thoracoabdominal aortic ectasia|Thoracoabdominal aortic ectasia
C0155763|T047|AB|447.8|ICD9CM|Arterial disease NEC|Arterial disease NEC
C0155763|T047|PT|447.8|ICD9CM|Other specified disorders of arteries and arterioles|Other specified disorders of arteries and arterioles
C0155764|T047|AB|447.9|ICD9CM|Arterial disease NOS|Arterial disease NOS
C0155764|T047|PT|447.9|ICD9CM|Unspecified disorders of arteries and arterioles|Unspecified disorders of arteries and arterioles
C0155765|T047|HT|448|ICD9CM|Disease of capillaries|Disease of capillaries
C0039445|T047|AB|448.0|ICD9CM|Heredit hemorr telangiec|Heredit hemorr telangiec
C0039445|T047|PT|448.0|ICD9CM|Hereditary hemorrhagic telangiectasia|Hereditary hemorrhagic telangiectasia
C0265027|T047|AB|448.1|ICD9CM|Nevus, non-neoplastic|Nevus, non-neoplastic
C0265027|T047|PT|448.1|ICD9CM|Nevus, non-neoplastic|Nevus, non-neoplastic
C0348651|T047|AB|448.9|ICD9CM|Capillary dis NEC/NOS|Capillary dis NEC/NOS
C0348651|T047|PT|448.9|ICD9CM|Other and unspecified capillary diseases|Other and unspecified capillary diseases
C1955786|T046|PT|449|ICD9CM|Septic arterial embolism|Septic arterial embolism
C1955786|T046|AB|449|ICD9CM|Septic arterial embolism|Septic arterial embolism
C1367972|T047|HT|451|ICD9CM|Phlebitis and thrombophlebitis|Phlebitis and thrombophlebitis
C0340270|T047|HT|451-459.99|ICD9CM|DISEASES OF VEINS AND LYMPHATICS, AND OTHER DISEASES OF CIRCULATORY SYSTEM|DISEASES OF VEINS AND LYMPHATICS, AND OTHER DISEASES OF CIRCULATORY SYSTEM
C0265057|T047|PT|451.0|ICD9CM|Phlebitis and thrombophlebitis of superficial vessels of lower extremities|Phlebitis and thrombophlebitis of superficial vessels of lower extremities
C0265057|T047|AB|451.0|ICD9CM|Superfic phlebitis-leg|Superfic phlebitis-leg
C0340711|T047|HT|451.1|ICD9CM|Phlebitis and thrombophlebitis of deep vessels of lower extremities|Phlebitis and thrombophlebitis of deep vessels of lower extremities
C0265066|T047|AB|451.11|ICD9CM|Femoral vein phlebitis|Femoral vein phlebitis
C0265066|T047|PT|451.11|ICD9CM|Phlebitis and thrombophlebitis of femoral vein (deep) (superficial)|Phlebitis and thrombophlebitis of femoral vein (deep) (superficial)
C0155770|T047|AB|451.19|ICD9CM|Deep phlebitis-leg NEC|Deep phlebitis-leg NEC
C0155770|T047|PT|451.19|ICD9CM|Phlebitis and thrombophlebitis of deep veins of lower extremities, other|Phlebitis and thrombophlebitis of deep veins of lower extremities, other
C0340712|T047|PT|451.2|ICD9CM|Phlebitis and thrombophlebitis of lower extremities, unspecified|Phlebitis and thrombophlebitis of lower extremities, unspecified
C0340712|T047|AB|451.2|ICD9CM|Thrombophlebitis leg NOS|Thrombophlebitis leg NOS
C0340692|T047|HT|451.8|ICD9CM|Phlebitis and thrombophlebitis of other sites|Phlebitis and thrombophlebitis of other sites
C0155772|T047|AB|451.81|ICD9CM|Iliac thrombophlebitis|Iliac thrombophlebitis
C0155772|T047|PT|451.81|ICD9CM|Phlebitis and thrombophlebitis of iliac vein|Phlebitis and thrombophlebitis of iliac vein
C0375311|T047|AB|451.82|ICD9CM|Phlbts sprfc vn up extrm|Phlbts sprfc vn up extrm
C0375311|T047|PT|451.82|ICD9CM|Phlebitis and thrombophlebitis of superficial veins of upper extremities|Phlebitis and thrombophlebitis of superficial veins of upper extremities
C0375312|T047|AB|451.83|ICD9CM|Phlbts deep vn up extrm|Phlbts deep vn up extrm
C0375312|T047|PT|451.83|ICD9CM|Phlebitis and thrombophlebitis of deep veins of upper extremities|Phlebitis and thrombophlebitis of deep veins of upper extremities
C0375313|T047|AB|451.84|ICD9CM|Phlbts vn NOS up extrm|Phlbts vn NOS up extrm
C0375313|T047|PT|451.84|ICD9CM|Phlebitis and thrombophlebitis of upper extremities, unspecified|Phlebitis and thrombophlebitis of upper extremities, unspecified
C0340692|T047|PT|451.89|ICD9CM|Phlebitis and thrombophlebitis of other sites|Phlebitis and thrombophlebitis of other sites
C0340692|T047|AB|451.89|ICD9CM|Thrombophlebitis NEC|Thrombophlebitis NEC
C1367972|T047|PT|451.9|ICD9CM|Phlebitis and thrombophlebitis of unspecified site|Phlebitis and thrombophlebitis of unspecified site
C1367972|T047|AB|451.9|ICD9CM|Thrombophlebitis NOS|Thrombophlebitis NOS
C0155773|T047|AB|452|ICD9CM|Portal vein thrombosis|Portal vein thrombosis
C0155773|T047|PT|452|ICD9CM|Portal vein thrombosis|Portal vein thrombosis
C0155774|T047|HT|453|ICD9CM|Other venous embolism and thrombosis|Other venous embolism and thrombosis
C0856761|T047|AB|453.0|ICD9CM|Budd-chiari syndrome|Budd-chiari syndrome
C0856761|T047|PT|453.0|ICD9CM|Budd-chiari syndrome|Budd-chiari syndrome
C0152250|T047|AB|453.1|ICD9CM|Thrombophlebitis migrans|Thrombophlebitis migrans
C0152250|T047|PT|453.1|ICD9CM|Thrombophlebitis migrans|Thrombophlebitis migrans
C2712843|T046|AB|453.2|ICD9CM|Oth inf vena cava thromb|Oth inf vena cava thromb
C2712843|T046|PT|453.2|ICD9CM|Other venous embolism and thrombosis of inferior vena cava|Other venous embolism and thrombosis of inferior vena cava
C0155776|T046|PT|453.3|ICD9CM|Other venous embolism and thrombosis of renal vein|Other venous embolism and thrombosis of renal vein
C0155776|T046|AB|453.3|ICD9CM|Renal vein thrombosis|Renal vein thrombosis
C2712859|T046|HT|453.4|ICD9CM|Acute venous embolism and thrombosis of deep vessels of lower extremity|Acute venous embolism and thrombosis of deep vessels of lower extremity
C2712629|T046|AB|453.40|ICD9CM|Ac DVT/embl low ext NOS|Ac DVT/embl low ext NOS
C2712629|T046|PT|453.40|ICD9CM|Acute venous embolism and thrombosis of unspecified deep vessels of lower extremity|Acute venous embolism and thrombosis of unspecified deep vessels of lower extremity
C2712619|T046|AB|453.41|ICD9CM|Ac DVT/emb prox low ext|Ac DVT/emb prox low ext
C2712619|T046|PT|453.41|ICD9CM|Acute venous embolism and thrombosis of deep vessels of proximal lower extremity|Acute venous embolism and thrombosis of deep vessels of proximal lower extremity
C2712631|T046|AB|453.42|ICD9CM|Ac DVT/emb distl low ext|Ac DVT/emb distl low ext
C2712631|T046|PT|453.42|ICD9CM|Acute venous embolism and thrombosis of deep vessels of distal lower extremity|Acute venous embolism and thrombosis of deep vessels of distal lower extremity
C2712872|T046|HT|453.5|ICD9CM|Chronic venous embolism and thrombosis of deep vessels of lower extremity|Chronic venous embolism and thrombosis of deep vessels of lower extremity
C2712815|T046|AB|453.50|ICD9CM|Ch DVT/embl low ext NOS|Ch DVT/embl low ext NOS
C2712815|T046|PT|453.50|ICD9CM|Chronic venous embolism and thrombosis of unspecified deep vessels of lower extremity|Chronic venous embolism and thrombosis of unspecified deep vessels of lower extremity
C2712828|T046|AB|453.51|ICD9CM|Ch DVT/embl prox low ext|Ch DVT/embl prox low ext
C2712828|T046|PT|453.51|ICD9CM|Chronic venous embolism and thrombosis of deep vessels of proximal lower extremity|Chronic venous embolism and thrombosis of deep vessels of proximal lower extremity
C2712817|T046|AB|453.52|ICD9CM|Ch DVT/embl dstl low ext|Ch DVT/embl dstl low ext
C2712817|T046|PT|453.52|ICD9CM|Chronic venous embolism and thrombosis of deep vessels of distal lower extremity|Chronic venous embolism and thrombosis of deep vessels of distal lower extremity
C2712884|T046|AB|453.6|ICD9CM|Embl suprfcl ves low ext|Embl suprfcl ves low ext
C2712884|T046|PT|453.6|ICD9CM|Venous embolism and thrombosis of superficial vessels of lower extremity|Venous embolism and thrombosis of superficial vessels of lower extremity
C2712896|T046|HT|453.7|ICD9CM|Chronic venous embolism and thrombosis of other specified vessels|Chronic venous embolism and thrombosis of other specified vessels
C2712938|T046|AB|453.71|ICD9CM|Ch emblsm suprfcl up ext|Ch emblsm suprfcl up ext
C2712938|T046|PT|453.71|ICD9CM|Chronic venous embolism and thrombosis of superficial veins of upper extremity|Chronic venous embolism and thrombosis of superficial veins of upper extremity
C2712948|T046|AB|453.72|ICD9CM|Ch DVT/embl up ext|Ch DVT/embl up ext
C2712948|T046|PT|453.72|ICD9CM|Chronic venous embolism and thrombosis of deep veins of upper extremity|Chronic venous embolism and thrombosis of deep veins of upper extremity
C2712966|T046|AB|453.73|ICD9CM|Ch emblsm up ext NOS|Ch emblsm up ext NOS
C2712966|T046|PT|453.73|ICD9CM|Chronic venous embolism and thrombosis of upper extremity, unspecified|Chronic venous embolism and thrombosis of upper extremity, unspecified
C2712953|T046|AB|453.74|ICD9CM|Ch emblsm axillary veins|Ch emblsm axillary veins
C2712953|T046|PT|453.74|ICD9CM|Chronic venous embolism and thrombosis of axillary veins|Chronic venous embolism and thrombosis of axillary veins
C2712755|T046|AB|453.75|ICD9CM|Ch emblsm subclav veins|Ch emblsm subclav veins
C2712755|T046|PT|453.75|ICD9CM|Chronic venous embolism and thrombosis of subclavian veins|Chronic venous embolism and thrombosis of subclavian veins
C2712765|T046|AB|453.76|ICD9CM|Ch embl internl jug vein|Ch embl internl jug vein
C2712765|T046|PT|453.76|ICD9CM|Chronic venous embolism and thrombosis of internal jugular veins|Chronic venous embolism and thrombosis of internal jugular veins
C2712794|T046|AB|453.77|ICD9CM|Ch embl thorac vein NEC|Ch embl thorac vein NEC
C2712794|T046|PT|453.77|ICD9CM|Chronic venous embolism and thrombosis of other thoracic veins|Chronic venous embolism and thrombosis of other thoracic veins
C2712814|T046|AB|453.79|ICD9CM|Ch emblsm veins NEC|Ch emblsm veins NEC
C2712814|T046|PT|453.79|ICD9CM|Chronic venous embolism and thrombosis of other specified veins|Chronic venous embolism and thrombosis of other specified veins
C2712996|T046|HT|453.8|ICD9CM|Acute venous embolism and thrombosis of other specified veins|Acute venous embolism and thrombosis of other specified veins
C2712822|T046|AB|453.81|ICD9CM|Ac embl suprfcl up ext|Ac embl suprfcl up ext
C2712822|T046|PT|453.81|ICD9CM|Acute venous embolism and thrombosis of superficial veins of upper extremity|Acute venous embolism and thrombosis of superficial veins of upper extremity
C2712834|T046|AB|453.82|ICD9CM|Ac DVT/embl up ext|Ac DVT/embl up ext
C2712834|T046|PT|453.82|ICD9CM|Acute venous embolism and thrombosis of deep veins of upper extremity|Acute venous embolism and thrombosis of deep veins of upper extremity
C2712845|T046|AB|453.83|ICD9CM|Ac emblsm up ext NOS|Ac emblsm up ext NOS
C2712845|T046|PT|453.83|ICD9CM|Acute venous embolism and thrombosis of upper extremity, unspecified|Acute venous embolism and thrombosis of upper extremity, unspecified
C2712855|T046|AB|453.84|ICD9CM|Ac emblsm axillary veins|Ac emblsm axillary veins
C2712855|T046|PT|453.84|ICD9CM|Acute venous embolism and thrombosis of axillary veins|Acute venous embolism and thrombosis of axillary veins
C2712847|T046|AB|453.85|ICD9CM|Ac embl subclav veins|Ac embl subclav veins
C2712847|T046|PT|453.85|ICD9CM|Acute venous embolism and thrombosis of subclavian veins|Acute venous embolism and thrombosis of subclavian veins
C2712858|T046|AB|453.86|ICD9CM|Ac embl internl jug vein|Ac embl internl jug vein
C2712858|T046|PT|453.86|ICD9CM|Acute venous embolism and thrombosis of internal jugular veins|Acute venous embolism and thrombosis of internal jugular veins
C2712704|T046|AB|453.87|ICD9CM|Ac embl thorac vein NEC|Ac embl thorac vein NEC
C2712704|T046|PT|453.87|ICD9CM|Acute venous embolism and thrombosis of other thoracic veins|Acute venous embolism and thrombosis of other thoracic veins
C2712736|T046|AB|453.89|ICD9CM|Ac embolism veins NEC|Ac embolism veins NEC
C2712736|T046|PT|453.89|ICD9CM|Acute venous embolism and thrombosis of other specified veins|Acute venous embolism and thrombosis of other specified veins
C0040038|T046|PT|453.9|ICD9CM|Other venous embolism and thrombosis of unspecified site|Other venous embolism and thrombosis of unspecified site
C0040038|T046|AB|453.9|ICD9CM|Venous thrombosis NOS|Venous thrombosis NOS
C0155778|T047|HT|454|ICD9CM|Varicose veins of lower extremities|Varicose veins of lower extremities
C0553570|T047|AB|454.0|ICD9CM|Leg varicosity w ulcer|Leg varicosity w ulcer
C0553570|T047|PT|454.0|ICD9CM|Varicose veins of lower extremities with ulcer|Varicose veins of lower extremities with ulcer
C0042347|T047|AB|454.1|ICD9CM|Leg varicosity w inflam|Leg varicosity w inflam
C0042347|T047|PT|454.1|ICD9CM|Varicose veins of lower extremities with inflammation|Varicose veins of lower extremities with inflammation
C0155779|T047|AB|454.2|ICD9CM|Varicos leg ulcer/inflam|Varicos leg ulcer/inflam
C0155779|T047|PT|454.2|ICD9CM|Varicose veins of lower extremities with ulcer and inflammation|Varicose veins of lower extremities with ulcer and inflammation
C1135217|T047|AB|454.8|ICD9CM|Varic vein leg,comp NEC|Varic vein leg,comp NEC
C1135217|T047|PT|454.8|ICD9CM|Varicose veins of lower extremities with other complications|Varicose veins of lower extremities with other complications
C1135335|T047|AB|454.9|ICD9CM|Asympt varicose veins|Asympt varicose veins
C1135335|T047|PT|454.9|ICD9CM|Asymptomatic varicose veins|Asymptomatic varicose veins
C0019112|T047|HT|455|ICD9CM|Hemorrhoids|Hemorrhoids
C0265035|T047|AB|455.0|ICD9CM|Int hemorrhoid w/o compl|Int hemorrhoid w/o compl
C0265035|T047|PT|455.0|ICD9CM|Internal hemorrhoids without mention of complication|Internal hemorrhoids without mention of complication
C0155781|T047|AB|455.1|ICD9CM|Int thrombos hemorrhoid|Int thrombos hemorrhoid
C0155781|T047|PT|455.1|ICD9CM|Internal thrombosed hemorrhoids|Internal thrombosed hemorrhoids
C0155782|T047|AB|455.2|ICD9CM|Int hemrrhoid w comp NEC|Int hemrrhoid w comp NEC
C0155782|T047|PT|455.2|ICD9CM|Internal hemorrhoids with other complication|Internal hemorrhoids with other complication
C0265041|T047|AB|455.3|ICD9CM|Ext hemorrhoid w/o compl|Ext hemorrhoid w/o compl
C0265041|T047|PT|455.3|ICD9CM|External hemorrhoids without mention of complication|External hemorrhoids without mention of complication
C0155784|T020|AB|455.4|ICD9CM|Ext thrombos hemorrhoid|Ext thrombos hemorrhoid
C0155784|T020|PT|455.4|ICD9CM|External thrombosed hemorrhoids|External thrombosed hemorrhoids
C0155785|T047|AB|455.5|ICD9CM|Ext hemrrhoid w comp NEC|Ext hemrrhoid w comp NEC
C0155785|T047|PT|455.5|ICD9CM|External hemorrhoids with other complication|External hemorrhoids with other complication
C0041844|T020|AB|455.6|ICD9CM|Hemorrhoids NOS|Hemorrhoids NOS
C0041844|T020|PT|455.6|ICD9CM|Unspecified hemorrhoids without mention of complication|Unspecified hemorrhoids without mention of complication
C0235326|T047|AB|455.7|ICD9CM|Thrombos hemorrhoids NOS|Thrombos hemorrhoids NOS
C0235326|T047|PT|455.7|ICD9CM|Unspecified thrombosed hemorrhoids|Unspecified thrombosed hemorrhoids
C0155787|T046|AB|455.8|ICD9CM|Hemrrhoid NOS w comp NEC|Hemrrhoid NOS w comp NEC
C0155787|T046|PT|455.8|ICD9CM|Unspecified hemorrhoids with other complication|Unspecified hemorrhoids with other complication
C0155788|T190|AB|455.9|ICD9CM|Residual hemorrhoid tags|Residual hemorrhoid tags
C0155788|T190|PT|455.9|ICD9CM|Residual hemorrhoidal skin tags|Residual hemorrhoidal skin tags
C0155797|T047|HT|456|ICD9CM|Varicose veins of other sites|Varicose veins of other sites
C0155789|T047|AB|456.0|ICD9CM|Esophag varices w bleed|Esophag varices w bleed
C0155789|T047|PT|456.0|ICD9CM|Esophageal varices with bleeding|Esophageal varices with bleeding
C0267092|T047|AB|456.1|ICD9CM|Esoph varices w/o bleed|Esoph varices w/o bleed
C0267092|T047|PT|456.1|ICD9CM|Esophageal varices without mention of bleeding|Esophageal varices without mention of bleeding
C0155791|T047|HT|456.2|ICD9CM|Esophageal varices in diseases classified elsewhere|Esophageal varices in diseases classified elsewhere
C0155792|T047|AB|456.20|ICD9CM|Bleed esoph var oth dis|Bleed esoph var oth dis
C0155792|T047|PT|456.20|ICD9CM|Esophageal varices in diseases classified elsewhere, with bleeding|Esophageal varices in diseases classified elsewhere, with bleeding
C0155793|T047|AB|456.21|ICD9CM|Esoph varice oth dis NOS|Esoph varice oth dis NOS
C0155793|T047|PT|456.21|ICD9CM|Esophageal varices in diseases classified elsewhere, without mention of bleeding|Esophageal varices in diseases classified elsewhere, without mention of bleeding
C0155794|T020|AB|456.3|ICD9CM|Sublingual varices|Sublingual varices
C0155794|T020|PT|456.3|ICD9CM|Sublingual varices|Sublingual varices
C0042341|T047|AB|456.4|ICD9CM|Scrotal varices|Scrotal varices
C0042341|T047|PT|456.4|ICD9CM|Scrotal varices|Scrotal varices
C0155795|T047|AB|456.5|ICD9CM|Pelvic varices|Pelvic varices
C0155795|T047|PT|456.5|ICD9CM|Pelvic varices|Pelvic varices
C0155796|T047|AB|456.6|ICD9CM|Vulval varices|Vulval varices
C0155796|T047|PT|456.6|ICD9CM|Vulval varices|Vulval varices
C0155797|T047|AB|456.8|ICD9CM|Varices of other sites|Varices of other sites
C0155797|T047|PT|456.8|ICD9CM|Varices of other sites|Varices of other sites
C0155799|T047|HT|457|ICD9CM|Noninfectious disorders of lymphatic channels|Noninfectious disorders of lymphatic channels
C0472692|T047|AB|457.0|ICD9CM|Postmastect lymphedema|Postmastect lymphedema
C0472692|T047|PT|457.0|ICD9CM|Postmastectomy lymphedema syndrome|Postmastectomy lymphedema syndrome
C0029659|T046|AB|457.1|ICD9CM|Other lymphedema|Other lymphedema
C0029659|T046|PT|457.1|ICD9CM|Other lymphedema|Other lymphedema
C0024225|T047|AB|457.2|ICD9CM|Lymphangitis|Lymphangitis
C0024225|T047|PT|457.2|ICD9CM|Lymphangitis|Lymphangitis
C0029673|T047|AB|457.8|ICD9CM|Noninfect lymph dis NEC|Noninfect lymph dis NEC
C0029673|T047|PT|457.8|ICD9CM|Other noninfectious disorders of lymphatic channels|Other noninfectious disorders of lymphatic channels
C0155799|T047|AB|457.9|ICD9CM|Noninfect lymph dis NOS|Noninfect lymph dis NOS
C0155799|T047|PT|457.9|ICD9CM|Unspecified noninfectious disorder of lymphatic channels|Unspecified noninfectious disorder of lymphatic channels
C0020649|T033|HT|458|ICD9CM|Hypotension|Hypotension
C0020651|T047|AB|458.0|ICD9CM|Orthostatic hypotension|Orthostatic hypotension
C0020651|T047|PT|458.0|ICD9CM|Orthostatic hypotension|Orthostatic hypotension
C0155800|T047|AB|458.1|ICD9CM|Chronic hypotension|Chronic hypotension
C0155800|T047|PT|458.1|ICD9CM|Chronic hypotension|Chronic hypotension
C0375314|T047|HT|458.2|ICD9CM|Iatrogenic hypotension|Iatrogenic hypotension
C1260413|T046|AB|458.21|ICD9CM|Hemododialysis hypotensn|Hemododialysis hypotensn
C1260413|T046|PT|458.21|ICD9CM|Hypotension of hemodialysis|Hypotension of hemodialysis
C1260414|T046|AB|458.29|ICD9CM|Iatrogenc hypotnsion NEC|Iatrogenc hypotnsion NEC
C1260414|T046|PT|458.29|ICD9CM|Other iatrogenic hypotension|Other iatrogenic hypotension
C0490007|T047|AB|458.8|ICD9CM|Hypotension NEC|Hypotension NEC
C0490007|T047|PT|458.8|ICD9CM|Other specified hypotension|Other specified hypotension
C0020649|T033|AB|458.9|ICD9CM|Hypotension NOS|Hypotension NOS
C0020649|T033|PT|458.9|ICD9CM|Hypotension, unspecified|Hypotension, unspecified
C0348668|T047|HT|459|ICD9CM|Other disorders of circulatory system|Other disorders of circulatory system
C0019080|T046|AB|459.0|ICD9CM|Hemorrhage NOS|Hemorrhage NOS
C0019080|T046|PT|459.0|ICD9CM|Hemorrhage, unspecified|Hemorrhage, unspecified
C0032807|T047|HT|459.1|ICD9CM|Postphlebitic syndrome|Postphlebitic syndrome
C1135218|T047|AB|459.10|ICD9CM|Postphlbtc synd w/o comp|Postphlbtc synd w/o comp
C1135218|T047|PT|459.10|ICD9CM|Postphlebetic syndrome without complications|Postphlebetic syndrome without complications
C1135219|T047|PT|459.11|ICD9CM|Postphlebetic syndrome with ulcer|Postphlebetic syndrome with ulcer
C1135219|T047|AB|459.11|ICD9CM|Postphlebtc synd w ulcer|Postphlebtc synd w ulcer
C1135220|T047|PT|459.12|ICD9CM|Postphlebetic syndrome with inflammation|Postphlebetic syndrome with inflammation
C1135220|T047|AB|459.12|ICD9CM|Postphlebtc syn w inflam|Postphlebtc syn w inflam
C1135221|T047|AB|459.13|ICD9CM|Postphl syn w ulc&inflam|Postphl syn w ulc&inflam
C1135221|T047|PT|459.13|ICD9CM|Postphlebetic syndrome with ulcer and inflammation|Postphlebetic syndrome with ulcer and inflammation
C1135222|T047|AB|459.19|ICD9CM|Postphleb synd comp NEC|Postphleb synd comp NEC
C1135222|T047|PT|459.19|ICD9CM|Postphlebetic syndrome with other complication|Postphlebetic syndrome with other complication
C0155802|T020|AB|459.2|ICD9CM|Compression of vein|Compression of vein
C0155802|T020|PT|459.2|ICD9CM|Compression of vein|Compression of vein
C1135223|T047|HT|459.3|ICD9CM|Chronic venous hypertension (idiopathic)|Chronic venous hypertension (idiopathic)
C1135224|T047|AB|459.30|ICD9CM|Chr venous hypr w/o comp|Chr venous hypr w/o comp
C1135224|T047|PT|459.30|ICD9CM|Chronic venous hypertension without complications|Chronic venous hypertension without complications
C1135225|T047|AB|459.31|ICD9CM|Chr venous hyper w ulcer|Chr venous hyper w ulcer
C1135225|T047|PT|459.31|ICD9CM|Chronic venous hypertension with ulcer|Chronic venous hypertension with ulcer
C1135226|T047|AB|459.32|ICD9CM|Chr venous hypr w inflam|Chr venous hypr w inflam
C1135226|T047|PT|459.32|ICD9CM|Chronic venous hypertension with inflammation|Chronic venous hypertension with inflammation
C1135227|T047|AB|459.33|ICD9CM|Chr ven hyp w ulc&inflam|Chr ven hyp w ulc&inflam
C1135227|T047|PT|459.33|ICD9CM|Chronic venous hypertension with ulcer and inflammation|Chronic venous hypertension with ulcer and inflammation
C1135228|T047|AB|459.39|ICD9CM|Chr venous hyp comp NEC|Chr venous hyp comp NEC
C1135228|T047|PT|459.39|ICD9CM|Chronic venous hypertension with other complication|Chronic venous hypertension with other complication
C0155803|T047|HT|459.8|ICD9CM|Other specified disorders of circulatory system|Other specified disorders of circulatory system
C0042485|T047|PT|459.81|ICD9CM|Venous (peripheral) insufficiency, unspecified|Venous (peripheral) insufficiency, unspecified
C0042485|T047|AB|459.81|ICD9CM|Venous insufficiency NOS|Venous insufficiency NOS
C0155803|T047|AB|459.89|ICD9CM|Circulatory disease NEC|Circulatory disease NEC
C0155803|T047|PT|459.89|ICD9CM|Other specified disorders of circulatory system|Other specified disorders of circulatory system
C0728936|T047|AB|459.9|ICD9CM|Circulatory disease NOS|Circulatory disease NOS
C0728936|T047|PT|459.9|ICD9CM|Unspecified circulatory system disorder|Unspecified circulatory system disorder
C0009443|T047|AB|460|ICD9CM|Acute nasopharyngitis|Acute nasopharyngitis
C0009443|T047|PT|460|ICD9CM|Acute nasopharyngitis [common cold]|Acute nasopharyngitis [common cold]
C0339901|T047|HT|460-466.99|ICD9CM|ACUTE RESPIRATORY INFECTIONS|ACUTE RESPIRATORY INFECTIONS
C0035204|T047|HT|460-519.99|ICD9CM|DISEASES OF THE RESPIRATORY SYSTEM|DISEASES OF THE RESPIRATORY SYSTEM
C0149512|T047|HT|461|ICD9CM|Acute sinusitis|Acute sinusitis
C0155804|T047|AB|461.0|ICD9CM|Ac maxillary sinusitis|Ac maxillary sinusitis
C0155804|T047|PT|461.0|ICD9CM|Acute maxillary sinusitis|Acute maxillary sinusitis
C0155805|T047|AB|461.1|ICD9CM|Ac frontal sinusitis|Ac frontal sinusitis
C0155805|T047|PT|461.1|ICD9CM|Acute frontal sinusitis|Acute frontal sinusitis
C0155806|T047|AB|461.2|ICD9CM|Ac ethmoidal sinusitis|Ac ethmoidal sinusitis
C0155806|T047|PT|461.2|ICD9CM|Acute ethmoidal sinusitis|Acute ethmoidal sinusitis
C0155807|T047|AB|461.3|ICD9CM|Ac sphenoidal sinusitis|Ac sphenoidal sinusitis
C0155807|T047|PT|461.3|ICD9CM|Acute sphenoidal sinusitis|Acute sphenoidal sinusitis
C0155808|T047|AB|461.8|ICD9CM|Other acute sinusitis|Other acute sinusitis
C0155808|T047|PT|461.8|ICD9CM|Other acute sinusitis|Other acute sinusitis
C0149512|T047|AB|461.9|ICD9CM|Acute sinusitis NOS|Acute sinusitis NOS
C0149512|T047|PT|461.9|ICD9CM|Acute sinusitis, unspecified|Acute sinusitis, unspecified
C0001344|T047|AB|462|ICD9CM|Acute pharyngitis|Acute pharyngitis
C0001344|T047|PT|462|ICD9CM|Acute pharyngitis|Acute pharyngitis
C0001361|T047|AB|463|ICD9CM|Acute tonsillitis|Acute tonsillitis
C0001361|T047|PT|463|ICD9CM|Acute tonsillitis|Acute tonsillitis
C0155811|T047|HT|464|ICD9CM|Acute laryngitis and tracheitis|Acute laryngitis and tracheitis
C0001327|T047|HT|464.0|ICD9CM|Acute laryngitis|Acute laryngitis
C0949122|T047|AB|464.00|ICD9CM|Ac laryngitis w/o obst|Ac laryngitis w/o obst
C0949122|T047|PT|464.00|ICD9CM|Acute laryngitis without mention of obstruction|Acute laryngitis without mention of obstruction
C0949123|T047|AB|464.01|ICD9CM|Ac laryngitis w obstruct|Ac laryngitis w obstruct
C0949123|T047|PT|464.01|ICD9CM|Acute laryngitis with obstruction|Acute laryngitis with obstruction
C0149513|T047|HT|464.1|ICD9CM|Acute tracheitis|Acute tracheitis
C0339877|T047|AB|464.10|ICD9CM|Ac tracheitis no obstruc|Ac tracheitis no obstruc
C0339877|T047|PT|464.10|ICD9CM|Acute tracheitis without mention of obstruction|Acute tracheitis without mention of obstruction
C0155810|T047|AB|464.11|ICD9CM|Ac tracheitis w obstruct|Ac tracheitis w obstruct
C0155810|T047|PT|464.11|ICD9CM|Acute tracheitis with obstruction|Acute tracheitis with obstruction
C0155811|T047|HT|464.2|ICD9CM|Acute laryngotracheitis|Acute laryngotracheitis
C0339876|T047|AB|464.20|ICD9CM|Ac laryngotrach no obstr|Ac laryngotrach no obstr
C0339876|T047|PT|464.20|ICD9CM|Acute laryngotracheitis without mention of obstruction|Acute laryngotracheitis without mention of obstruction
C0155813|T047|AB|464.21|ICD9CM|Ac laryngotrach w obstr|Ac laryngotrach w obstr
C0155813|T047|PT|464.21|ICD9CM|Acute laryngotracheitis with obstruction|Acute laryngotracheitis with obstruction
C0155814|T047|HT|464.3|ICD9CM|Acute epiglottitis|Acute epiglottitis
C0396041|T047|AB|464.30|ICD9CM|Ac epiglottitis no obstr|Ac epiglottitis no obstr
C0396041|T047|PT|464.30|ICD9CM|Acute epiglottitis without mention of obstruction|Acute epiglottitis without mention of obstruction
C0155815|T047|AB|464.31|ICD9CM|Ac epiglottitis w obstr|Ac epiglottitis w obstr
C0155815|T047|PT|464.31|ICD9CM|Acute epiglottitis with obstruction|Acute epiglottitis with obstruction
C0010380|T047|AB|464.4|ICD9CM|Croup|Croup
C0010380|T047|PT|464.4|ICD9CM|Croup|Croup
C0749165|T047|HT|464.5|ICD9CM|Supraglottitis, unspecified|Supraglottitis, unspecified
C2887377|T047|AB|464.50|ICD9CM|Supraglottis w/o obs NOS|Supraglottis w/o obs NOS
C2887377|T047|PT|464.50|ICD9CM|Supraglottitis unspecified, without obstruction|Supraglottitis unspecified, without obstruction
C0949126|T047|AB|464.51|ICD9CM|Supraglottis w obstr NOS|Supraglottis w obstr NOS
C0949126|T047|PT|464.51|ICD9CM|Supraglottitis unspecified, with obstruction|Supraglottitis unspecified, with obstruction
C0155816|T047|HT|465|ICD9CM|Acute upper respiratory infections of multiple or unspecified sites|Acute upper respiratory infections of multiple or unspecified sites
C0155817|T047|AB|465.0|ICD9CM|Acute laryngopharyngitis|Acute laryngopharyngitis
C0155817|T047|PT|465.0|ICD9CM|Acute laryngopharyngitis|Acute laryngopharyngitis
C0155818|T047|PT|465.8|ICD9CM|Acute upper respiratory infections of other multiple sites|Acute upper respiratory infections of other multiple sites
C0155818|T047|AB|465.8|ICD9CM|Acute uri mult sites NEC|Acute uri mult sites NEC
C0264222|T047|PT|465.9|ICD9CM|Acute upper respiratory infections of unspecified site|Acute upper respiratory infections of unspecified site
C0264222|T047|AB|465.9|ICD9CM|Acute uri NOS|Acute uri NOS
C0155820|T047|HT|466|ICD9CM|Acute bronchitis and bronchiolitis|Acute bronchitis and bronchiolitis
C0149514|T047|AB|466.0|ICD9CM|Acute bronchitis|Acute bronchitis
C0149514|T047|PT|466.0|ICD9CM|Acute bronchitis|Acute bronchitis
C0001311|T047|HT|466.1|ICD9CM|Acute bronchiolitis|Acute bronchiolitis
C0348799|T047|AB|466.11|ICD9CM|Acu broncholitis d/t RSV|Acu broncholitis d/t RSV
C0348799|T047|PT|466.11|ICD9CM|Acute bronchiolitis due to respiratory syncytial virus (RSV)|Acute bronchiolitis due to respiratory syncytial virus (RSV)
C0375319|T047|AB|466.19|ICD9CM|Acu brnchlts d/t oth org|Acu brnchlts d/t oth org
C0375319|T047|PT|466.19|ICD9CM|Acute bronchiolitis due to other infectious organisms|Acute bronchiolitis due to other infectious organisms
C0549397|T033|AB|470|ICD9CM|Deviated nasal septum|Deviated nasal septum
C0549397|T033|PT|470|ICD9CM|Deviated nasal septum|Deviated nasal septum
C0155839|T047|HT|470-478.99|ICD9CM|OTHER DISEASES OF THE UPPER RESPIRATORY TRACT|OTHER DISEASES OF THE UPPER RESPIRATORY TRACT
C0027430|T047|HT|471|ICD9CM|Nasal polyps|Nasal polyps
C0027430|T047|AB|471.0|ICD9CM|Polyp of nasal cavity|Polyp of nasal cavity
C0027430|T047|PT|471.0|ICD9CM|Polyp of nasal cavity|Polyp of nasal cavity
C0155822|T047|AB|471.1|ICD9CM|Polypoid sinus degen|Polypoid sinus degen
C0155822|T047|PT|471.1|ICD9CM|Polypoid sinus degeneration|Polypoid sinus degeneration
C0155823|T047|AB|471.8|ICD9CM|Nasal sinus polyp NEC|Nasal sinus polyp NEC
C0155823|T047|PT|471.8|ICD9CM|Other polyp of sinus|Other polyp of sinus
C0027430|T047|AB|471.9|ICD9CM|Nasal polyp NOS|Nasal polyp NOS
C0027430|T047|PT|471.9|ICD9CM|Unspecified nasal polyp|Unspecified nasal polyp
C0155824|T047|HT|472|ICD9CM|Chronic pharyngitis and nasopharyngitis|Chronic pharyngitis and nasopharyngitis
C0008711|T047|AB|472.0|ICD9CM|Chronic rhinitis|Chronic rhinitis
C0008711|T047|PT|472.0|ICD9CM|Chronic rhinitis|Chronic rhinitis
C0155825|T047|AB|472.1|ICD9CM|Chronic pharyngitis|Chronic pharyngitis
C0155825|T047|PT|472.1|ICD9CM|Chronic pharyngitis|Chronic pharyngitis
C0155826|T047|AB|472.2|ICD9CM|Chronic nasopharyngitis|Chronic nasopharyngitis
C0155826|T047|PT|472.2|ICD9CM|Chronic nasopharyngitis|Chronic nasopharyngitis
C0149516|T047|HT|473|ICD9CM|Chronic sinusitis|Chronic sinusitis
C0008698|T047|AB|473.0|ICD9CM|Chr maxillary sinusitis|Chr maxillary sinusitis
C0008698|T047|PT|473.0|ICD9CM|Chronic maxillary sinusitis|Chronic maxillary sinusitis
C0008683|T047|AB|473.1|ICD9CM|Chr frontal sinusitis|Chr frontal sinusitis
C0008683|T047|PT|473.1|ICD9CM|Chronic frontal sinusitis|Chronic frontal sinusitis
C0008681|T047|AB|473.2|ICD9CM|Chr ethmoidal sinusitis|Chr ethmoidal sinusitis
C0008681|T047|PT|473.2|ICD9CM|Chronic ethmoidal sinusitis|Chronic ethmoidal sinusitis
C0008712|T047|AB|473.3|ICD9CM|Chr sphenoidal sinusitis|Chr sphenoidal sinusitis
C0008712|T047|PT|473.3|ICD9CM|Chronic sphenoidal sinusitis|Chronic sphenoidal sinusitis
C0395986|T047|AB|473.8|ICD9CM|Chronic sinusitis NEC|Chronic sinusitis NEC
C0395986|T047|PT|473.8|ICD9CM|Other chronic sinusitis|Other chronic sinusitis
C0149516|T047|AB|473.9|ICD9CM|Chronic sinusitis NOS|Chronic sinusitis NOS
C0149516|T047|PT|473.9|ICD9CM|Unspecified sinusitis (chronic)|Unspecified sinusitis (chronic)
C0155828|T047|HT|474|ICD9CM|Chronic disease of tonsils and adenoids|Chronic disease of tonsils and adenoids
C0490040|T047|HT|474.0|ICD9CM|Chronic tonsillitis and adenoiditis|Chronic tonsillitis and adenoiditis
C0149517|T047|AB|474.00|ICD9CM|Chronic tonsillitis|Chronic tonsillitis
C0149517|T047|PT|474.00|ICD9CM|Chronic tonsillitis|Chronic tonsillitis
C0396023|T047|AB|474.01|ICD9CM|Chronic adenoiditis|Chronic adenoiditis
C0396023|T047|PT|474.01|ICD9CM|Chronic adenoiditis|Chronic adenoiditis
C0490040|T047|PT|474.02|ICD9CM|Chronic tonsillitis and adenoiditis|Chronic tonsillitis and adenoiditis
C0490040|T047|AB|474.02|ICD9CM|Chronic tonsils&adenoids|Chronic tonsils&adenoids
C0155829|T047|HT|474.1|ICD9CM|Hypertrophy of tonsils and adenoids|Hypertrophy of tonsils and adenoids
C0155829|T047|PT|474.10|ICD9CM|Hypertrophy of tonsil with adenoids|Hypertrophy of tonsil with adenoids
C0155829|T047|AB|474.10|ICD9CM|Hypertrophy T and A|Hypertrophy T and A
C0155831|T047|PT|474.11|ICD9CM|Hypertrophy of tonsils alone|Hypertrophy of tonsils alone
C0155831|T047|AB|474.11|ICD9CM|Hypertrophy tonsils|Hypertrophy tonsils
C0149825|T047|AB|474.12|ICD9CM|Hypertrophy adenoids|Hypertrophy adenoids
C0149825|T047|PT|474.12|ICD9CM|Hypertrophy of adenoids alone|Hypertrophy of adenoids alone
C0155833|T047|AB|474.2|ICD9CM|Adenoid vegetations|Adenoid vegetations
C0155833|T047|PT|474.2|ICD9CM|Adenoid vegetations|Adenoid vegetations
C0155834|T047|AB|474.8|ICD9CM|Chr T & A dis NEC|Chr T & A dis NEC
C0155834|T047|PT|474.8|ICD9CM|Other chronic disease of tonsils and adenoids|Other chronic disease of tonsils and adenoids
C0155828|T047|AB|474.9|ICD9CM|Chr T & A dis NOS|Chr T & A dis NOS
C0155828|T047|PT|474.9|ICD9CM|Unspecified chronic disease of tonsils and adenoids|Unspecified chronic disease of tonsils and adenoids
C0031157|T047|AB|475|ICD9CM|Peritonsillar abscess|Peritonsillar abscess
C0031157|T047|PT|475|ICD9CM|Peritonsillar abscess|Peritonsillar abscess
C0155835|T047|HT|476|ICD9CM|Chronic laryngitis and laryngotracheitis|Chronic laryngitis and laryngotracheitis
C0155836|T047|AB|476.0|ICD9CM|Chronic laryngitis|Chronic laryngitis
C0155836|T047|PT|476.0|ICD9CM|Chronic laryngitis|Chronic laryngitis
C0155837|T047|AB|476.1|ICD9CM|Chr laryngotracheitis|Chr laryngotracheitis
C0155837|T047|PT|476.1|ICD9CM|Chronic laryngotracheitis|Chronic laryngotracheitis
C2607914|T047|HT|477|ICD9CM|Allergic rhinitis|Allergic rhinitis
C0018621|T047|PT|477.0|ICD9CM|Allergic rhinitis due to pollen|Allergic rhinitis due to pollen
C0018621|T047|AB|477.0|ICD9CM|Rhinitis due to pollen|Rhinitis due to pollen
C0878694|T047|PT|477.1|ICD9CM|Allergic rhinitis due to food|Allergic rhinitis due to food
C0878694|T047|AB|477.1|ICD9CM|Allergic rhinitis-food|Allergic rhinitis-food
C1456066|T047|AB|477.2|ICD9CM|Allerg rhinitis-cat/dog|Allerg rhinitis-cat/dog
C1456066|T047|PT|477.2|ICD9CM|Allergic rhinitis due to animal (cat) (dog) hair and dander|Allergic rhinitis due to animal (cat) (dog) hair and dander
C2712343|T047|PT|477.8|ICD9CM|Allergic rhinitis due to other allergen|Allergic rhinitis due to other allergen
C2712343|T047|AB|477.8|ICD9CM|Allergic rhinitis NEC|Allergic rhinitis NEC
C2607914|T047|AB|477.9|ICD9CM|Allergic rhinitis NOS|Allergic rhinitis NOS
C2607914|T047|PT|477.9|ICD9CM|Allergic rhinitis, cause unspecified|Allergic rhinitis, cause unspecified
C0155839|T047|HT|478|ICD9CM|Other diseases of upper respiratory tract|Other diseases of upper respiratory tract
C0155840|T047|PT|478.0|ICD9CM|Hypertrophy of nasal turbinates|Hypertrophy of nasal turbinates
C0155840|T047|AB|478.0|ICD9CM|Hypertrph nasal turbinat|Hypertrph nasal turbinat
C0029581|T047|HT|478.1|ICD9CM|Other diseases of nasal cavity and sinuses|Other diseases of nasal cavity and sinuses
C0235963|T047|AB|478.11|ICD9CM|Nasal mucositis (ulcer)|Nasal mucositis (ulcer)
C0235963|T047|PT|478.11|ICD9CM|Nasal mucositis (ulcerative)|Nasal mucositis (ulcerative)
C0029581|T047|AB|478.19|ICD9CM|Nasal & sinus dis NEC|Nasal & sinus dis NEC
C0029581|T047|PT|478.19|ICD9CM|Other disease of nasal cavity and sinuses|Other disease of nasal cavity and sinuses
C0795699|T047|HT|478.2|ICD9CM|Other diseases of pharynx, not elsewhere classified|Other diseases of pharynx, not elsewhere classified
C0031345|T047|AB|478.20|ICD9CM|Disease of pharynx NOS|Disease of pharynx NOS
C0031345|T047|PT|478.20|ICD9CM|Unspecified disease of pharynx|Unspecified disease of pharynx
C0155841|T047|AB|478.21|ICD9CM|Cellulitis of pharynx|Cellulitis of pharynx
C0155841|T047|PT|478.21|ICD9CM|Cellulitis of pharynx or nasopharynx|Cellulitis of pharynx or nasopharynx
C0155842|T047|AB|478.22|ICD9CM|Parapharyngeal abscess|Parapharyngeal abscess
C0155842|T047|PT|478.22|ICD9CM|Parapharyngeal abscess|Parapharyngeal abscess
C0155843|T047|AB|478.24|ICD9CM|Retropharyngeal abscess|Retropharyngeal abscess
C0155843|T047|PT|478.24|ICD9CM|Retropharyngeal abscess|Retropharyngeal abscess
C0155844|T047|PT|478.25|ICD9CM|Edema of pharynx or nasopharynx|Edema of pharynx or nasopharynx
C0155844|T047|AB|478.25|ICD9CM|Edema pharynx/nasopharyx|Edema pharynx/nasopharyx
C0155845|T047|PT|478.26|ICD9CM|Cyst of pharynx or nasopharynx|Cyst of pharynx or nasopharynx
C0155845|T047|AB|478.26|ICD9CM|Cyst pharynx/nasopharynx|Cyst pharynx/nasopharynx
C0795699|T047|AB|478.29|ICD9CM|Disease of pharynx NEC|Disease of pharynx NEC
C0795699|T047|PT|478.29|ICD9CM|Other diseases of pharynx, not elsewhere classified|Other diseases of pharynx, not elsewhere classified
C0494657|T047|HT|478.3|ICD9CM|Paralysis of vocal cords or larynx|Paralysis of vocal cords or larynx
C0042928|T047|PT|478.30|ICD9CM|Paralysis of vocal cords or larynx, unspecified|Paralysis of vocal cords or larynx, unspecified
C0042928|T047|AB|478.30|ICD9CM|Vocal cord paralysis NOS|Vocal cord paralysis NOS
C0155847|T047|PT|478.31|ICD9CM|Unilateral paralysis of vocal cords or larynx, partial|Unilateral paralysis of vocal cords or larynx, partial
C0155847|T047|AB|478.31|ICD9CM|Vocal paral unilat part|Vocal paral unilat part
C0155848|T047|PT|478.32|ICD9CM|Unilateral paralysis of vocal cords or larynx, complete|Unilateral paralysis of vocal cords or larynx, complete
C0155848|T047|AB|478.32|ICD9CM|Vocal paral unilat total|Vocal paral unilat total
C0155849|T047|PT|478.33|ICD9CM|Bilateral paralysis of vocal cords or larynx, partial|Bilateral paralysis of vocal cords or larynx, partial
C0155849|T047|AB|478.33|ICD9CM|Vocal paral bilat part|Vocal paral bilat part
C0155850|T047|PT|478.34|ICD9CM|Bilateral paralysis of vocal cords or larynx, complete|Bilateral paralysis of vocal cords or larynx, complete
C0155850|T047|AB|478.34|ICD9CM|Vocal paral bilat total|Vocal paral bilat total
C0155851|T047|PT|478.4|ICD9CM|Polyp of vocal cord or larynx|Polyp of vocal cord or larynx
C0155851|T047|AB|478.4|ICD9CM|Vocal cord/larynx polyp|Vocal cord/larynx polyp
C0155852|T047|PT|478.5|ICD9CM|Other diseases of vocal cords|Other diseases of vocal cords
C0155852|T047|AB|478.5|ICD9CM|Vocal cord disease NEC|Vocal cord disease NEC
C0023052|T046|AB|478.6|ICD9CM|Edema of larynx|Edema of larynx
C0023052|T046|PT|478.6|ICD9CM|Edema of larynx|Edema of larynx
C1561612|T047|HT|478.7|ICD9CM|Other diseases of larynx, not elsewhere classified|Other diseases of larynx, not elsewhere classified
C0023051|T047|AB|478.70|ICD9CM|Disease of larynx NOS|Disease of larynx NOS
C0023051|T047|PT|478.70|ICD9CM|Unspecified disease of larynx|Unspecified disease of larynx
C0155853|T047|PT|478.71|ICD9CM|Cellulitis and perichondritis of larynx|Cellulitis and perichondritis of larynx
C0155853|T047|AB|478.71|ICD9CM|Laryngeal cellulitis|Laryngeal cellulitis
C0023075|T047|AB|478.74|ICD9CM|Stenosis of larynx|Stenosis of larynx
C0023075|T047|PT|478.74|ICD9CM|Stenosis of larynx|Stenosis of larynx
C0023066|T047|AB|478.75|ICD9CM|Laryngeal spasm|Laryngeal spasm
C0023066|T047|PT|478.75|ICD9CM|Laryngeal spasm|Laryngeal spasm
C1561612|T047|AB|478.79|ICD9CM|Disease of larynx NEC|Disease of larynx NEC
C1561612|T047|PT|478.79|ICD9CM|Other diseases of larynx, not elsewhere classified|Other diseases of larynx, not elsewhere classified
C0375321|T047|PT|478.8|ICD9CM|Upper respiratory tract hypersensitivity reaction, site unspecified|Upper respiratory tract hypersensitivity reaction, site unspecified
C0375321|T047|AB|478.8|ICD9CM|Urt hypersens react NOS|Urt hypersens react NOS
C0155839|T047|PT|478.9|ICD9CM|Other and unspecified diseases of upper respiratory tract|Other and unspecified diseases of upper respiratory tract
C0155839|T047|AB|478.9|ICD9CM|Upper resp dis NEC/NOS|Upper resp dis NEC/NOS
C0032310|T047|HT|480|ICD9CM|Viral pneumonia|Viral pneumonia
C0155870|T047|HT|480-488.99|ICD9CM|PNEUMONIA AND INFLUENZA|PNEUMONIA AND INFLUENZA
C0276156|T047|AB|480.0|ICD9CM|Adenoviral pneumonia|Adenoviral pneumonia
C0276156|T047|PT|480.0|ICD9CM|Pneumonia due to adenovirus|Pneumonia due to adenovirus
C0152413|T047|PT|480.1|ICD9CM|Pneumonia due to respiratory syncytial virus|Pneumonia due to respiratory syncytial virus
C0152413|T047|AB|480.1|ICD9CM|Resp syncyt viral pneum|Resp syncyt viral pneum
C0276333|T047|AB|480.2|ICD9CM|Parinfluenza viral pneum|Parinfluenza viral pneum
C0276333|T047|PT|480.2|ICD9CM|Pneumonia due to parainfluenza virus|Pneumonia due to parainfluenza virus
C1260415|T047|AB|480.3|ICD9CM|Pneumonia due to SARS|Pneumonia due to SARS
C1260415|T047|PT|480.3|ICD9CM|Pneumonia due to SARS-associated coronavirus|Pneumonia due to SARS-associated coronavirus
C0302377|T047|PT|480.8|ICD9CM|Pneumonia due to other virus not elsewhere classified|Pneumonia due to other virus not elsewhere classified
C0302377|T047|AB|480.8|ICD9CM|Viral pneumonia NEC|Viral pneumonia NEC
C0032310|T047|AB|480.9|ICD9CM|Viral pneumonia NOS|Viral pneumonia NOS
C0032310|T047|PT|480.9|ICD9CM|Viral pneumonia, unspecified|Viral pneumonia, unspecified
C0155862|T047|AB|481|ICD9CM|Pneumococcal pneumonia|Pneumococcal pneumonia
C0155862|T047|PT|481|ICD9CM|Pneumococcal pneumonia [Streptococcus pneumoniae pneumonia]|Pneumococcal pneumonia [Streptococcus pneumoniae pneumonia]
C0155858|T047|HT|482|ICD9CM|Other bacterial pneumonia|Other bacterial pneumonia
C0519030|T047|AB|482.0|ICD9CM|K. pneumoniae pneumonia|K. pneumoniae pneumonia
C0519030|T047|PT|482.0|ICD9CM|Pneumonia due to Klebsiella pneumoniae|Pneumonia due to Klebsiella pneumoniae
C0155860|T047|PT|482.1|ICD9CM|Pneumonia due to Pseudomonas|Pneumonia due to Pseudomonas
C0155860|T047|AB|482.1|ICD9CM|Pseudomonal pneumonia|Pseudomonal pneumonia
C0276026|T047|AB|482.2|ICD9CM|H.influenzae pneumonia|H.influenzae pneumonia
C0276026|T047|PT|482.2|ICD9CM|Pneumonia due to Hemophilus influenzae [H. influenzae]|Pneumonia due to Hemophilus influenzae [H. influenzae]
C0155862|T047|HT|482.3|ICD9CM|Pneumonia due to Streptococcus|Pneumonia due to Streptococcus
C0155862|T047|PT|482.30|ICD9CM|Pneumonia due to Streptococcus, unspecified|Pneumonia due to Streptococcus, unspecified
C0155862|T047|AB|482.30|ICD9CM|Streptococcal pneumn NOS|Streptococcal pneumn NOS
C0375324|T047|PT|482.31|ICD9CM|Pneumonia due to Streptococcus, group A|Pneumonia due to Streptococcus, group A
C0375324|T047|AB|482.31|ICD9CM|Pneumonia strptococcus a|Pneumonia strptococcus a
C0348801|T047|PT|482.32|ICD9CM|Pneumonia due to Streptococcus, group B|Pneumonia due to Streptococcus, group B
C0348801|T047|AB|482.32|ICD9CM|Pneumonia strptococcus b|Pneumonia strptococcus b
C0375326|T047|PT|482.39|ICD9CM|Pneumonia due to other Streptococcus|Pneumonia due to other Streptococcus
C0375326|T047|AB|482.39|ICD9CM|Pneumonia oth strep|Pneumonia oth strep
C0032308|T047|HT|482.4|ICD9CM|Pneumonia due to Staphylococcus|Pneumonia due to Staphylococcus
C0032308|T047|PT|482.40|ICD9CM|Pneumonia due to Staphylococcus, unspecified|Pneumonia due to Staphylococcus, unspecified
C0032308|T047|AB|482.40|ICD9CM|Staphylococcal pneu NOS|Staphylococcal pneu NOS
C2349529|T047|AB|482.41|ICD9CM|Meth sus pneum d/t Staph|Meth sus pneum d/t Staph
C2349529|T047|PT|482.41|ICD9CM|Methicillin susceptible pneumonia due to Staphylococcus aureus|Methicillin susceptible pneumonia due to Staphylococcus aureus
C1142536|T047|AB|482.42|ICD9CM|Meth res pneu d/t Staph|Meth res pneu d/t Staph
C1142536|T047|PT|482.42|ICD9CM|Methicillin resistant pneumonia due to Staphylococcus aureus|Methicillin resistant pneumonia due to Staphylococcus aureus
C0695234|T047|PT|482.49|ICD9CM|Other Staphylococcus pneumonia|Other Staphylococcus pneumonia
C0695234|T047|AB|482.49|ICD9CM|Staph pneumonia NEC|Staph pneumonia NEC
C0032286|T047|HT|482.8|ICD9CM|Pneumonia due to other specified bacteria|Pneumonia due to other specified bacteria
C0375327|T047|AB|482.81|ICD9CM|Pneumonia anaerobes|Pneumonia anaerobes
C0375327|T047|PT|482.81|ICD9CM|Pneumonia due to anaerobes|Pneumonia due to anaerobes
C0276089|T047|PT|482.82|ICD9CM|Pneumonia due to escherichia coli [E. coli]|Pneumonia due to escherichia coli [E. coli]
C0276089|T047|AB|482.82|ICD9CM|Pneumonia e coli|Pneumonia e coli
C0854248|T047|AB|482.83|ICD9CM|Pneumo oth grm-neg bact|Pneumo oth grm-neg bact
C0854248|T047|PT|482.83|ICD9CM|Pneumonia due to other gram-negative bacteria|Pneumonia due to other gram-negative bacteria
C0023241|T047|AB|482.84|ICD9CM|Legionnaires' disease|Legionnaires' disease
C0023241|T047|PT|482.84|ICD9CM|Pneumonia due to Legionnaires' disease|Pneumonia due to Legionnaires' disease
C0032286|T047|PT|482.89|ICD9CM|Pneumonia due to other specified bacteria|Pneumonia due to other specified bacteria
C0032286|T047|AB|482.89|ICD9CM|Pneumonia oth spcf bact|Pneumonia oth spcf bact
C0004626|T047|AB|482.9|ICD9CM|Bacterial pneumonia NOS|Bacterial pneumonia NOS
C0004626|T047|PT|482.9|ICD9CM|Bacterial pneumonia, unspecified|Bacterial pneumonia, unspecified
C0032287|T047|HT|483|ICD9CM|Pneumonia due to other specified organism|Pneumonia due to other specified organism
C0032302|T047|AB|483.0|ICD9CM|Pneu mycplsm pneumoniae|Pneu mycplsm pneumoniae
C0032302|T047|PT|483.0|ICD9CM|Pneumonia due to mycoplasma pneumoniae|Pneumonia due to mycoplasma pneumoniae
C0339959|T047|AB|483.1|ICD9CM|Pneumonia d/t chlamydia|Pneumonia d/t chlamydia
C0339959|T047|PT|483.1|ICD9CM|Pneumonia due to chlamydia|Pneumonia due to chlamydia
C0032287|T047|AB|483.8|ICD9CM|Pneumon oth spec orgnsm|Pneumon oth spec orgnsm
C0032287|T047|PT|483.8|ICD9CM|Pneumonia due to other specified organism|Pneumonia due to other specified organism
C0155863|T047|HT|484|ICD9CM|Pneumonia in infectious diseases classified elsewhere|Pneumonia in infectious diseases classified elsewhere
C0276253|T047|AB|484.1|ICD9CM|Pneum w cytomeg incl dis|Pneum w cytomeg incl dis
C0276253|T047|PT|484.1|ICD9CM|Pneumonia in cytomegalic inclusion disease|Pneumonia in cytomegalic inclusion disease
C0155865|T047|AB|484.3|ICD9CM|Pneumonia in whoop cough|Pneumonia in whoop cough
C0155865|T047|PT|484.3|ICD9CM|Pneumonia in whooping cough|Pneumonia in whooping cough
C0155866|T047|AB|484.5|ICD9CM|Pneumonia in anthrax|Pneumonia in anthrax
C0155866|T047|PT|484.5|ICD9CM|Pneumonia in anthrax|Pneumonia in anthrax
C0155867|T047|AB|484.6|ICD9CM|Pneum in aspergillosis|Pneum in aspergillosis
C0155867|T047|PT|484.6|ICD9CM|Pneumonia in aspergillosis|Pneumonia in aspergillosis
C0155868|T047|AB|484.7|ICD9CM|Pneum in oth sys mycoses|Pneum in oth sys mycoses
C0155868|T047|PT|484.7|ICD9CM|Pneumonia in other systemic mycoses|Pneumonia in other systemic mycoses
C0155869|T047|AB|484.8|ICD9CM|Pneum in infect dis NEC|Pneum in infect dis NEC
C0155869|T047|PT|484.8|ICD9CM|Pneumonia in other infectious diseases classified elsewhere|Pneumonia in other infectious diseases classified elsewhere
C0006285|T047|AB|485|ICD9CM|Bronchopneumonia org NOS|Bronchopneumonia org NOS
C0006285|T047|PT|485|ICD9CM|Bronchopneumonia, organism unspecified|Bronchopneumonia, organism unspecified
C0339951|T047|AB|486|ICD9CM|Pneumonia, organism NOS|Pneumonia, organism NOS
C0339951|T047|PT|486|ICD9CM|Pneumonia, organism unspecified|Pneumonia, organism unspecified
C0021400|T047|HT|487|ICD9CM|Influenza|Influenza
C0155870|T047|AB|487.0|ICD9CM|Influenza with pneumonia|Influenza with pneumonia
C0155870|T047|PT|487.0|ICD9CM|Influenza with pneumonia|Influenza with pneumonia
C0021414|T047|AB|487.1|ICD9CM|Flu w resp manifest NEC|Flu w resp manifest NEC
C0021414|T047|PT|487.1|ICD9CM|Influenza with other respiratory manifestations|Influenza with other respiratory manifestations
C0155871|T047|AB|487.8|ICD9CM|Flu w manifestation NEC|Flu w manifestation NEC
C0155871|T047|PT|487.8|ICD9CM|Influenza with other manifestations|Influenza with other manifestations
C2712970|T047|HT|488|ICD9CM|Influenza due to certain identified influenza viruses|Influenza due to certain identified influenza viruses
C2712881|T047|HT|488.0|ICD9CM|Influenza due to identified avian influenza virus|Influenza due to identified avian influenza virus
C2921085|T047|AB|488.01|ICD9CM|Flu dt iden avian w pneu|Flu dt iden avian w pneu
C2921085|T047|PT|488.01|ICD9CM|Influenza due to identified avian influenza virus with pneumonia|Influenza due to identified avian influenza virus with pneumonia
C2921090|T047|AB|488.02|ICD9CM|Flu dt avian w oth resp|Flu dt avian w oth resp
C2921090|T047|PT|488.02|ICD9CM|Influenza due to identified avian influenza virus with other respiratory manifestations|Influenza due to identified avian influenza virus with other respiratory manifestations
C2887385|T047|AB|488.09|ICD9CM|Flu dt avian manfest NEC|Flu dt avian manfest NEC
C2887385|T047|PT|488.09|ICD9CM|Influenza due to identified avian influenza virus with other manifestations|Influenza due to identified avian influenza virus with other manifestations
C3161430|T047|HT|488.1|ICD9CM|Influenza due to identified 2009 H1N1 influenza virus|Influenza due to identified 2009 H1N1 influenza virus
C3161333|T047|AB|488.11|ICD9CM|Flu dt 2009 H1N1 w pneu|Flu dt 2009 H1N1 w pneu
C3161333|T047|PT|488.11|ICD9CM|Influenza due to identified 2009 H1N1 influenza virus with pneumonia|Influenza due to identified 2009 H1N1 influenza virus with pneumonia
C3161334|T047|AB|488.12|ICD9CM|Flu-2009 H1N1 w oth resp|Flu-2009 H1N1 w oth resp
C3161334|T047|PT|488.12|ICD9CM|Influenza due to identified 2009 H1N1 influenza virus with other respiratory manifestations|Influenza due to identified 2009 H1N1 influenza virus with other respiratory manifestations
C2887395|T047|AB|488.19|ICD9CM|Flu-2009 H1N1 w oth man|Flu-2009 H1N1 w oth man
C2887395|T047|PT|488.19|ICD9CM|Influenza due to identified 2009 H1N1 influenza virus with other manifestations|Influenza due to identified 2009 H1N1 influenza virus with other manifestations
C3161252|T047|HT|488.8|ICD9CM|Influenza due to novel influenza A|Influenza due to novel influenza A
C3161093|T047|AB|488.81|ICD9CM|Flu dt nvl A vrs w pneu|Flu dt nvl A vrs w pneu
C3161093|T047|PT|488.81|ICD9CM|Influenza due to identified novel influenza A virus with pneumonia|Influenza due to identified novel influenza A virus with pneumonia
C3161094|T047|AB|488.82|ICD9CM|Flu dt nvl A w oth resp|Flu dt nvl A w oth resp
C3161094|T047|PT|488.82|ICD9CM|Influenza due to identified novel influenza A virus with other respiratory manifestations|Influenza due to identified novel influenza A virus with other respiratory manifestations
C3161095|T047|AB|488.89|ICD9CM|Flu dt novel A w oth man|Flu dt novel A w oth man
C3161095|T047|PT|488.89|ICD9CM|Influenza due to identified novel influenza A virus with other manifestations|Influenza due to identified novel influenza A virus with other manifestations
C0006277|T047|AB|490|ICD9CM|Bronchitis NOS|Bronchitis NOS
C0006277|T047|PT|490|ICD9CM|Bronchitis, not specified as acute or chronic|Bronchitis, not specified as acute or chronic
C0178278|T047|HT|490-496.99|ICD9CM|CHRONIC OBSTRUCTIVE PULMONARY DISEASE AND ALLIED CONDITIONS|CHRONIC OBSTRUCTIVE PULMONARY DISEASE AND ALLIED CONDITIONS
C0008677|T047|HT|491|ICD9CM|Chronic bronchitis|Chronic bronchitis
C0155872|T047|AB|491.0|ICD9CM|Simple chr bronchitis|Simple chr bronchitis
C0155872|T047|PT|491.0|ICD9CM|Simple chronic bronchitis|Simple chronic bronchitis
C0155873|T047|AB|491.1|ICD9CM|Mucopurul chr bronchitis|Mucopurul chr bronchitis
C0155873|T047|PT|491.1|ICD9CM|Mucopurulent chronic bronchitis|Mucopurulent chronic bronchitis
C0155874|T047|HT|491.2|ICD9CM|Obstructive chronic bronchitis|Obstructive chronic bronchitis
C0155875|T047|AB|491.20|ICD9CM|Obst chr bronc w/o exac|Obst chr bronc w/o exac
C0155875|T047|PT|491.20|ICD9CM|Obstructive chronic bronchitis without exacerbation|Obstructive chronic bronchitis without exacerbation
C4041147|T047|AB|491.21|ICD9CM|Obs chr bronc w(ac) exac|Obs chr bronc w(ac) exac
C4041147|T047|PT|491.21|ICD9CM|Obstructive chronic bronchitis with (acute) exacerbation|Obstructive chronic bronchitis with (acute) exacerbation
C1456131|T047|AB|491.22|ICD9CM|Obs chr bronc w ac bronc|Obs chr bronc w ac bronc
C1456131|T047|PT|491.22|ICD9CM|Obstructive chronic bronchitis with acute bronchitis|Obstructive chronic bronchitis with acute bronchitis
C0029544|T047|AB|491.8|ICD9CM|Chronic bronchitis NEC|Chronic bronchitis NEC
C0029544|T047|PT|491.8|ICD9CM|Other chronic bronchitis|Other chronic bronchitis
C0008677|T047|AB|491.9|ICD9CM|Chronic bronchitis NOS|Chronic bronchitis NOS
C0008677|T047|PT|491.9|ICD9CM|Unspecified chronic bronchitis|Unspecified chronic bronchitis
C0034067|T047|HT|492|ICD9CM|Emphysema|Emphysema
C0152242|T033|AB|492.0|ICD9CM|Emphysematous bleb|Emphysematous bleb
C0152242|T033|PT|492.0|ICD9CM|Emphysematous bleb|Emphysematous bleb
C0029607|T047|AB|492.8|ICD9CM|Emphysema NEC|Emphysema NEC
C0029607|T047|PT|492.8|ICD9CM|Other emphysema|Other emphysema
C0004096|T047|HT|493|ICD9CM|Asthma|Asthma
C0155877|T047|HT|493.0|ICD9CM|Extrinsic asthma|Extrinsic asthma
C0155878|T047|AB|493.00|ICD9CM|Extrinsic asthma NOS|Extrinsic asthma NOS
C0155878|T047|PT|493.00|ICD9CM|Extrinsic asthma, unspecified|Extrinsic asthma, unspecified
C0155879|T047|AB|493.01|ICD9CM|Ext asthma w status asth|Ext asthma w status asth
C0155879|T047|PT|493.01|ICD9CM|Extrinsic asthma with status asthmaticus|Extrinsic asthma with status asthmaticus
C1176339|T047|AB|493.02|ICD9CM|Ext asthma w(acute) exac|Ext asthma w(acute) exac
C1176339|T047|PT|493.02|ICD9CM|Extrinsic asthma with (acute) exacerbation|Extrinsic asthma with (acute) exacerbation
C0155880|T047|HT|493.1|ICD9CM|Intrinsic asthma|Intrinsic asthma
C0155881|T047|AB|493.10|ICD9CM|Intrinsic asthma NOS|Intrinsic asthma NOS
C0155881|T047|PT|493.10|ICD9CM|Intrinsic asthma, unspecified|Intrinsic asthma, unspecified
C0155882|T047|AB|493.11|ICD9CM|Int asthma w status asth|Int asthma w status asth
C0155882|T047|PT|493.11|ICD9CM|Intrinsic asthma with status asthmaticus|Intrinsic asthma with status asthmaticus
C1176340|T047|AB|493.12|ICD9CM|Int asthma w (ac) exac|Int asthma w (ac) exac
C1176340|T047|PT|493.12|ICD9CM|Intrinsic asthma with (acute) exacerbation|Intrinsic asthma with (acute) exacerbation
C0155883|T047|HT|493.2|ICD9CM|Chronic obstructive asthma|Chronic obstructive asthma
C0375333|T047|AB|493.20|ICD9CM|Chronic obst asthma NOS|Chronic obst asthma NOS
C0375333|T047|PT|493.20|ICD9CM|Chronic obstructive asthma, unspecified|Chronic obstructive asthma, unspecified
C0375334|T047|AB|493.21|ICD9CM|Ch ob asthma w stat asth|Ch ob asthma w stat asth
C0375334|T047|PT|493.21|ICD9CM|Chronic obstructive asthma with status asthmaticus|Chronic obstructive asthma with status asthmaticus
C1176341|T047|AB|493.22|ICD9CM|Ch obst asth w (ac) exac|Ch obst asth w (ac) exac
C1176341|T047|PT|493.22|ICD9CM|Chronic obstructive asthma with (acute) exacerbation|Chronic obstructive asthma with (acute) exacerbation
C1260416|T047|HT|493.8|ICD9CM|Other forms of asthma|Other forms of asthma
C0015263|T047|PT|493.81|ICD9CM|Exercise induced bronchospasm|Exercise induced bronchospasm
C0015263|T047|AB|493.81|ICD9CM|Exercse ind bronchospasm|Exercse ind bronchospasm
C0694548|T047|AB|493.82|ICD9CM|Cough variant asthma|Cough variant asthma
C0694548|T047|PT|493.82|ICD9CM|Cough variant asthma|Cough variant asthma
C0004096|T047|HT|493.9|ICD9CM|Asthma, unspecified|Asthma, unspecified
C0155886|T047|AB|493.90|ICD9CM|Asthma NOS|Asthma NOS
C0155886|T047|PT|493.90|ICD9CM|Asthma, unspecified type, unspecified|Asthma, unspecified type, unspecified
C0038218|T047|AB|493.91|ICD9CM|Asthma w status asthmat|Asthma w status asthmat
C0038218|T047|PT|493.91|ICD9CM|Asthma, unspecified type, with status asthmaticus|Asthma, unspecified type, with status asthmaticus
C1176342|T047|AB|493.92|ICD9CM|Asthma NOS w (ac) exac|Asthma NOS w (ac) exac
C1176342|T047|PT|493.92|ICD9CM|Asthma, unspecified type, with (acute) exacerbation|Asthma, unspecified type, with (acute) exacerbation
C0006267|T047|HT|494|ICD9CM|Bronchiectasis|Bronchiectasis
C0878695|T047|AB|494.0|ICD9CM|Bronchiectas w/o ac exac|Bronchiectas w/o ac exac
C0878695|T047|PT|494.0|ICD9CM|Bronchiectasis without acute exacerbation|Bronchiectasis without acute exacerbation
C0878696|T047|AB|494.1|ICD9CM|Bronchiectasis w ac exac|Bronchiectasis w ac exac
C0878696|T047|PT|494.1|ICD9CM|Bronchiectasis with acute exacerbation|Bronchiectasis with acute exacerbation
C0002390|T047|HT|495|ICD9CM|Extrinsic allergic alveolitis|Extrinsic allergic alveolitis
C0015634|T047|AB|495.0|ICD9CM|Farmers' lung|Farmers' lung
C0015634|T047|PT|495.0|ICD9CM|Farmers' lung|Farmers' lung
C0004681|T047|AB|495.1|ICD9CM|Bagassosis|Bagassosis
C0004681|T047|PT|495.1|ICD9CM|Bagassosis|Bagassosis
C0005592|T047|AB|495.2|ICD9CM|Bird-fanciers' lung|Bird-fanciers' lung
C0005592|T047|PT|495.2|ICD9CM|Bird-fanciers' lung|Bird-fanciers' lung
C0152108|T047|AB|495.3|ICD9CM|Suberosis|Suberosis
C0152108|T047|PT|495.3|ICD9CM|Suberosis|Suberosis
C0155888|T047|AB|495.4|ICD9CM|Malt workers' lung|Malt workers' lung
C0155888|T047|PT|495.4|ICD9CM|Malt workers' lung|Malt workers' lung
C0155889|T047|AB|495.5|ICD9CM|Mushroom workers' lung|Mushroom workers' lung
C0155889|T047|PT|495.5|ICD9CM|Mushroom workers' lung|Mushroom workers' lung
C0155890|T047|AB|495.6|ICD9CM|Mapl bark-stripprs' lung|Mapl bark-stripprs' lung
C0155890|T047|PT|495.6|ICD9CM|Maple bark-strippers' lung|Maple bark-strippers' lung
C0155891|T047|AB|495.7|ICD9CM|"ventilation" pneumonit|"ventilation" pneumonit
C0155891|T047|PT|495.7|ICD9CM|"Ventilation" pneumonitis|"Ventilation" pneumonitis
C0155892|T047|AB|495.8|ICD9CM|Allerg alveol/pneum NEC|Allerg alveol/pneum NEC
C0155892|T047|PT|495.8|ICD9CM|Other specified allergic alveolitis and pneumonitis|Other specified allergic alveolitis and pneumonitis
C0002390|T047|AB|495.9|ICD9CM|Allerg alveol/pneum NOS|Allerg alveol/pneum NOS
C0002390|T047|PT|495.9|ICD9CM|Unspecified allergic alveolitis and pneumonitis|Unspecified allergic alveolitis and pneumonitis
C0302378|T047|AB|496|ICD9CM|Chr airway obstruct NEC|Chr airway obstruct NEC
C0302378|T047|PT|496|ICD9CM|Chronic airway obstruction, not elsewhere classified|Chronic airway obstruction, not elsewhere classified
C0003165|T047|AB|500|ICD9CM|Coal workers' pneumocon|Coal workers' pneumocon
C0003165|T047|PT|500|ICD9CM|Coal workers' pneumoconiosis|Coal workers' pneumoconiosis
C0178279|T047|HT|500-508.99|ICD9CM|PNEUMOCONIOSES AND OTHER LUNG DISEASES DUE TO EXTERNAL AGENTS|PNEUMOCONIOSES AND OTHER LUNG DISEASES DUE TO EXTERNAL AGENTS
C0003949|T047|AB|501|ICD9CM|Asbestosis|Asbestosis
C0003949|T047|PT|501|ICD9CM|Asbestosis|Asbestosis
C0037116|T047|PT|502|ICD9CM|Pneumoconiosis due to other silica or silicates|Pneumoconiosis due to other silica or silicates
C0037116|T047|AB|502|ICD9CM|Silica pneumocon NEC|Silica pneumocon NEC
C0032274|T047|AB|503|ICD9CM|Inorg dust pneumocon NEC|Inorg dust pneumocon NEC
C0032274|T047|PT|503|ICD9CM|Pneumoconiosis due to other inorganic dust|Pneumoconiosis due to other inorganic dust
C0032318|T047|AB|504|ICD9CM|Dust pneumonopathy NEC|Dust pneumonopathy NEC
C0032318|T047|PT|504|ICD9CM|Pneumonopathy due to inhalation of other dust|Pneumonopathy due to inhalation of other dust
C0032273|T047|AB|505|ICD9CM|Pneumoconiosis NOS|Pneumoconiosis NOS
C0032273|T047|PT|505|ICD9CM|Pneumoconiosis, unspecified|Pneumoconiosis, unspecified
C0155893|T047|HT|506|ICD9CM|Respiratory conditions due to chemical fumes and vapors|Respiratory conditions due to chemical fumes and vapors
C0155894|T047|PT|506.0|ICD9CM|Bronchitis and pneumonitis due to fumes and vapors|Bronchitis and pneumonitis due to fumes and vapors
C0155894|T047|AB|506.0|ICD9CM|Fum/vapor bronc/pneumon|Fum/vapor bronc/pneumon
C0155895|T047|PT|506.1|ICD9CM|Acute pulmonary edema due to fumes and vapors|Acute pulmonary edema due to fumes and vapors
C0155895|T047|AB|506.1|ICD9CM|Fum/vapor ac pulm edema|Fum/vapor ac pulm edema
C0155896|T047|AB|506.2|ICD9CM|Fum/vapor up resp inflam|Fum/vapor up resp inflam
C0155896|T047|PT|506.2|ICD9CM|Upper respiratory inflammation due to fumes and vapors|Upper respiratory inflammation due to fumes and vapors
C0155897|T047|AB|506.3|ICD9CM|Fum/vap ac resp cond NEC|Fum/vap ac resp cond NEC
C0155897|T047|PT|506.3|ICD9CM|Other acute and subacute respiratory conditions due to fumes and vapors|Other acute and subacute respiratory conditions due to fumes and vapors
C0155898|T047|PT|506.4|ICD9CM|Chronic respiratory conditions due to fumes and vapors|Chronic respiratory conditions due to fumes and vapors
C0155898|T047|AB|506.4|ICD9CM|Fum/vapor chr resp cond|Fum/vapor chr resp cond
C0041881|T047|AB|506.9|ICD9CM|Fum/vapor resp cond NOS|Fum/vapor resp cond NOS
C0041881|T047|PT|506.9|ICD9CM|Unspecified respiratory conditions due to fumes and vapors|Unspecified respiratory conditions due to fumes and vapors
C0155899|T047|HT|507|ICD9CM|Pneumonitis due to solids and liquids|Pneumonitis due to solids and liquids
C0260334|T047|AB|507.0|ICD9CM|Food/vomit pneumonitis|Food/vomit pneumonitis
C0260334|T047|PT|507.0|ICD9CM|Pneumonitis due to inhalation of food or vomitus|Pneumonitis due to inhalation of food or vomitus
C0494675|T047|AB|507.1|ICD9CM|Oil/essence pneumonitis|Oil/essence pneumonitis
C0494675|T047|PT|507.1|ICD9CM|Pneumonitis due to inhalation of oils and essences|Pneumonitis due to inhalation of oils and essences
C0155900|T047|PT|507.8|ICD9CM|Pneumonitis due to other solids and liquids|Pneumonitis due to other solids and liquids
C0155900|T047|AB|507.8|ICD9CM|Solid/liq pneumonit NEC|Solid/liq pneumonit NEC
C0155901|T046|HT|508|ICD9CM|Respiratory conditions due to other and unspecified external agents|Respiratory conditions due to other and unspecified external agents
C0155902|T046|AB|508.0|ICD9CM|Ac pul manif d/t radiat|Ac pul manif d/t radiat
C0155902|T046|PT|508.0|ICD9CM|Acute pulmonary manifestations due to radiation|Acute pulmonary manifestations due to radiation
C0155903|T046|AB|508.1|ICD9CM|Chr pul manif d/t radiat|Chr pul manif d/t radiat
C0155903|T046|PT|508.1|ICD9CM|Chronic and other pulmonary manifestations due to radiation|Chronic and other pulmonary manifestations due to radiation
C3161096|T047|AB|508.2|ICD9CM|Resp cond dt smoke inhal|Resp cond dt smoke inhal
C3161096|T047|PT|508.2|ICD9CM|Respiratory conditions due to smoke inhalation|Respiratory conditions due to smoke inhalation
C0155904|T047|AB|508.8|ICD9CM|Resp cond: ext agent NEC|Resp cond: ext agent NEC
C0155904|T047|PT|508.8|ICD9CM|Respiratory conditions due to other specified external agents|Respiratory conditions due to other specified external agents
C0155905|T047|AB|508.9|ICD9CM|Resp cond: ext agent NOS|Resp cond: ext agent NOS
C0155905|T047|PT|508.9|ICD9CM|Respiratory conditions due to unspecified external agent|Respiratory conditions due to unspecified external agent
C0014009|T047|HT|510|ICD9CM|Empyema|Empyema
C0029582|T047|HT|510-519.99|ICD9CM|OTHER DISEASES OF RESPIRATORY SYSTEM|OTHER DISEASES OF RESPIRATORY SYSTEM
C0740253|T047|AB|510.0|ICD9CM|Empyema with fistula|Empyema with fistula
C0740253|T047|PT|510.0|ICD9CM|Empyema with fistula|Empyema with fistula
C0730032|T047|AB|510.9|ICD9CM|Empyema w/o fistula|Empyema w/o fistula
C0730032|T047|PT|510.9|ICD9CM|Empyema without mention of fistula|Empyema without mention of fistula
C0032231|T047|HT|511|ICD9CM|Pleurisy|Pleurisy
C0032232|T047|AB|511.0|ICD9CM|Pleurisy w/o effus or TB|Pleurisy w/o effus or TB
C0032232|T047|PT|511.0|ICD9CM|Pleurisy without mention of effusion or current tuberculosis|Pleurisy without mention of effusion or current tuberculosis
C0155906|T047|AB|511.1|ICD9CM|Bact pleur/effus not TB|Bact pleur/effus not TB
C0155906|T047|PT|511.1|ICD9CM|Pleurisy with effusion, with mention of a bacterial cause other than tuberculosis|Pleurisy with effusion, with mention of a bacterial cause other than tuberculosis
C0029799|T047|HT|511.8|ICD9CM|Other specified forms of pleural effusion, except tuberculous|Other specified forms of pleural effusion, except tuberculous
C0080032|T047|PT|511.81|ICD9CM|Malignant pleural effusion|Malignant pleural effusion
C0080032|T047|AB|511.81|ICD9CM|Malignant pleural effusn|Malignant pleural effusn
C2349532|T047|AB|511.89|ICD9CM|Effusion NEC exc tb|Effusion NEC exc tb
C2349532|T047|PT|511.89|ICD9CM|Other specified forms of effusion, except tuberculous|Other specified forms of effusion, except tuberculous
C0032227|T047|AB|511.9|ICD9CM|Pleural effusion NOS|Pleural effusion NOS
C0032227|T047|PT|511.9|ICD9CM|Unspecified pleural effusion|Unspecified pleural effusion
C3161433|T047|HT|512|ICD9CM|Pneumothorax and air leak|Pneumothorax and air leak
C0155907|T047|AB|512.0|ICD9CM|Spont tens pneumothorax|Spont tens pneumothorax
C0155907|T047|PT|512.0|ICD9CM|Spontaneous tension pneumothorax|Spontaneous tension pneumothorax
C0375336|T047|AB|512.1|ICD9CM|Iatrogenic pneumothorax|Iatrogenic pneumothorax
C0375336|T047|PT|512.1|ICD9CM|Iatrogenic pneumothorax|Iatrogenic pneumothorax
C3161097|T046|AB|512.2|ICD9CM|Postoperative air leak|Postoperative air leak
C3161097|T046|PT|512.2|ICD9CM|Postoperative air leak|Postoperative air leak
C3161434|T047|HT|512.8|ICD9CM|Other pneumothorax and air leak|Other pneumothorax and air leak
C1868193|T047|AB|512.81|ICD9CM|Prim spont pneumothorax|Prim spont pneumothorax
C1868193|T047|PT|512.81|ICD9CM|Primary spontaneous pneumothorax|Primary spontaneous pneumothorax
C3161098|T047|AB|512.82|ICD9CM|Sec spont pneumothorax|Sec spont pneumothorax
C3161098|T047|PT|512.82|ICD9CM|Secondary spontaneous pneumothorax|Secondary spontaneous pneumothorax
C0264557|T047|AB|512.83|ICD9CM|Chronic pneumothorax|Chronic pneumothorax
C0264557|T047|PT|512.83|ICD9CM|Chronic pneumothorax|Chronic pneumothorax
C3161099|T033|AB|512.84|ICD9CM|Other air leak|Other air leak
C3161099|T033|PT|512.84|ICD9CM|Other air leak|Other air leak
C0348708|T047|AB|512.89|ICD9CM|Other pneumothorax|Other pneumothorax
C0348708|T047|PT|512.89|ICD9CM|Other pneumothorax|Other pneumothorax
C0155908|T047|HT|513|ICD9CM|Abscess of lung and mediastinum|Abscess of lung and mediastinum
C0024110|T047|AB|513.0|ICD9CM|Abscess of lung|Abscess of lung
C0024110|T047|PT|513.0|ICD9CM|Abscess of lung|Abscess of lung
C0155909|T047|AB|513.1|ICD9CM|Abscess of mediastinum|Abscess of mediastinum
C0155909|T047|PT|513.1|ICD9CM|Abscess of mediastinum|Abscess of mediastinum
C0155910|T047|AB|514|ICD9CM|Pulm congest/hypostasis|Pulm congest/hypostasis
C0155910|T047|PT|514|ICD9CM|Pulmonary congestion and hypostasis|Pulmonary congestion and hypostasis
C0175999|T047|AB|515|ICD9CM|Postinflam pulm fibrosis|Postinflam pulm fibrosis
C0175999|T047|PT|515|ICD9CM|Postinflammatory pulmonary fibrosis|Postinflammatory pulmonary fibrosis
C0859814|T047|HT|516|ICD9CM|Other alveolar and parietoalveolar pneumonopathy|Other alveolar and parietoalveolar pneumonopathy
C0034050|T047|AB|516.0|ICD9CM|Pul alveolar proteinosis|Pul alveolar proteinosis
C0034050|T047|PT|516.0|ICD9CM|Pulmonary alveolar proteinosis|Pulmonary alveolar proteinosis
C0020807|T047|AB|516.1|ICD9CM|Idio pulm hemosiderosis|Idio pulm hemosiderosis
C0020807|T047|PT|516.1|ICD9CM|Idiopathic pulmonary hemosiderosis|Idiopathic pulmonary hemosiderosis
C0155912|T047|AB|516.2|ICD9CM|Pulm alveolar microlith|Pulm alveolar microlith
C0155912|T047|PT|516.2|ICD9CM|Pulmonary alveolar microlithiasis|Pulmonary alveolar microlithiasis
C2350236|T047|HT|516.3|ICD9CM|Idiopathic interstitial pneumonia|Idiopathic interstitial pneumonia
C3161100|T046|AB|516.30|ICD9CM|Idiopath inters pneu NOS|Idiopath inters pneu NOS
C3161100|T046|PT|516.30|ICD9CM|Idiopathic interstitial pneumonia, not otherwise specified|Idiopathic interstitial pneumonia, not otherwise specified
C1800706|T047|AB|516.31|ICD9CM|Idiopath pulmon fibrosis|Idiopath pulmon fibrosis
C1800706|T047|PT|516.31|ICD9CM|Idiopathic pulmonary fibrosis|Idiopathic pulmonary fibrosis
C3161102|T047|AB|516.32|ICD9CM|Idio non-spec inter pneu|Idio non-spec inter pneu
C3161102|T047|PT|516.32|ICD9CM|Idiopathic non-specific interstitial pneumonitis|Idiopathic non-specific interstitial pneumonitis
C1279945|T047|AB|516.33|ICD9CM|Acute interstitial pneum|Acute interstitial pneum
C1279945|T047|PT|516.33|ICD9CM|Acute interstitial pneumonitis|Acute interstitial pneumonitis
C0238378|T047|AB|516.34|ICD9CM|Resp brncio interst lung|Resp brncio interst lung
C0238378|T047|PT|516.34|ICD9CM|Respiratory bronchiolitis interstitial lung disease|Respiratory bronchiolitis interstitial lung disease
C3161103|T047|PT|516.35|ICD9CM|Idiopathic lymphoid interstitial pneumonia|Idiopathic lymphoid interstitial pneumonia
C3161103|T047|AB|516.35|ICD9CM|Idiopth lym interst pneu|Idiopth lym interst pneu
C0242770|T047|AB|516.36|ICD9CM|Cryptogenic organiz pneu|Cryptogenic organiz pneu
C0242770|T047|PT|516.36|ICD9CM|Cryptogenic organizing pneumonia|Cryptogenic organizing pneumonia
C0238378|T047|PT|516.37|ICD9CM|Desquamative interstitial pneumonia|Desquamative interstitial pneumonia
C0238378|T047|AB|516.37|ICD9CM|Desquamatv interst pneu|Desquamatv interst pneu
C0751674|T191|PT|516.4|ICD9CM|Lymphangioleiomyomatosis|Lymphangioleiomyomatosis
C0751674|T191|AB|516.4|ICD9CM|Lymphangioleiomyomatosis|Lymphangioleiomyomatosis
C3161104|T047|AB|516.5|ICD9CM|Adlt pul Langs cell hist|Adlt pul Langs cell hist
C3161104|T047|PT|516.5|ICD9CM|Adult pulmonary Langerhans cell histiocytosis|Adult pulmonary Langerhans cell histiocytosis
C3161253|T047|HT|516.6|ICD9CM|Interstitial lung diseases of childhood|Interstitial lung diseases of childhood
C3161105|T047|AB|516.61|ICD9CM|Neuroend cell hyprpl inf|Neuroend cell hyprpl inf
C3161105|T047|PT|516.61|ICD9CM|Neuroendocrine cell hyperplasia of infancy|Neuroendocrine cell hyperplasia of infancy
C3161106|T047|AB|516.62|ICD9CM|Pulm interstitl glycogen|Pulm interstitl glycogen
C3161106|T047|PT|516.62|ICD9CM|Pulmonary interstitial glycogenosis|Pulmonary interstitial glycogenosis
C3161107|T047|AB|516.63|ICD9CM|Surfactant mutation lung|Surfactant mutation lung
C3161107|T047|PT|516.63|ICD9CM|Surfactant mutations of the lung|Surfactant mutations of the lung
C3161108|T047|AB|516.64|ICD9CM|Alv cap dysp w vn misaln|Alv cap dysp w vn misaln
C3161108|T047|PT|516.64|ICD9CM|Alveolar capillary dysplasia with vein misalignment|Alveolar capillary dysplasia with vein misalignment
C3161109|T047|AB|516.69|ICD9CM|Oth intrst lung dis chld|Oth intrst lung dis chld
C3161109|T047|PT|516.69|ICD9CM|Other interstitial lung diseases of childhood|Other interstitial lung diseases of childhood
C0155913|T047|AB|516.8|ICD9CM|Alveol pneumonopathy NEC|Alveol pneumonopathy NEC
C0155913|T047|PT|516.8|ICD9CM|Other specified alveolar and parietoalveolar pneumonopathies|Other specified alveolar and parietoalveolar pneumonopathies
C0155914|T047|AB|516.9|ICD9CM|Alveol pneumonopathy NOS|Alveol pneumonopathy NOS
C0155914|T047|PT|516.9|ICD9CM|Unspecified alveolar and parietoalveolar pneumonopathy|Unspecified alveolar and parietoalveolar pneumonopathy
C0155915|T047|HT|517|ICD9CM|Lung involvement in conditions classified elsewhere|Lung involvement in conditions classified elsewhere
C0152450|T047|AB|517.1|ICD9CM|Rheumatic pneumonia|Rheumatic pneumonia
C0152450|T047|PT|517.1|ICD9CM|Rheumatic pneumonia|Rheumatic pneumonia
C0339904|T047|PT|517.2|ICD9CM|Lung involvement in systemic sclerosis|Lung involvement in systemic sclerosis
C0339904|T047|AB|517.2|ICD9CM|Syst sclerosis lung dis|Syst sclerosis lung dis
C0742343|T047|AB|517.3|ICD9CM|Acute chest syndrome|Acute chest syndrome
C0742343|T047|PT|517.3|ICD9CM|Acute chest syndrome|Acute chest syndrome
C0155917|T047|AB|517.8|ICD9CM|Lung involv in oth dis|Lung involv in oth dis
C0155917|T047|PT|517.8|ICD9CM|Lung involvement in other diseases classified elsewhere|Lung involvement in other diseases classified elsewhere
C0348712|T047|HT|518|ICD9CM|Other diseases of lung|Other diseases of lung
C0004144|T046|AB|518.0|ICD9CM|Pulmonary collapse|Pulmonary collapse
C0004144|T046|PT|518.0|ICD9CM|Pulmonary collapse|Pulmonary collapse
C1370824|T047|AB|518.1|ICD9CM|Interstitial emphysema|Interstitial emphysema
C1370824|T047|PT|518.1|ICD9CM|Interstitial emphysema|Interstitial emphysema
C0155918|T047|AB|518.2|ICD9CM|Compensatory emphysema|Compensatory emphysema
C0155918|T047|PT|518.2|ICD9CM|Compensatory emphysema|Compensatory emphysema
C0034068|T047|AB|518.3|ICD9CM|Pulmonary eosinophilia|Pulmonary eosinophilia
C0034068|T047|PT|518.3|ICD9CM|Pulmonary eosinophilia|Pulmonary eosinophilia
C0155919|T047|PT|518.4|ICD9CM|Acute edema of lung, unspecified|Acute edema of lung, unspecified
C0155919|T047|AB|518.4|ICD9CM|Acute lung edema NOS|Acute lung edema NOS
C0034076|T047|HT|518.5|ICD9CM|Pulmonary insufficiency following trauma and surgery|Pulmonary insufficiency following trauma and surgery
C3161110|T047|AB|518.51|ICD9CM|Ac resp flr fol trma/srg|Ac resp flr fol trma/srg
C3161110|T047|PT|518.51|ICD9CM|Acute respiratory failure following trauma and surgery|Acute respiratory failure following trauma and surgery
C3161111|T046|AB|518.52|ICD9CM|Ot pul insuf fol trm/srg|Ot pul insuf fol trm/srg
C3161111|T046|PT|518.52|ICD9CM|Other pulmonary insufficiency, not elsewhere classified, following trauma and surgery|Other pulmonary insufficiency, not elsewhere classified, following trauma and surgery
C3161112|T047|AB|518.53|ICD9CM|Ac/chr rsp flr fol tr/sg|Ac/chr rsp flr fol tr/sg
C3161112|T047|PT|518.53|ICD9CM|Acute and chronic respiratory failure following trauma and surgery|Acute and chronic respiratory failure following trauma and surgery
C0004031|T047|PT|518.6|ICD9CM|Allergic bronchopulmonary aspergillosis|Allergic bronchopulmonary aspergillosis
C0004031|T047|AB|518.6|ICD9CM|Alrgc brncpul asprglosis|Alrgc brncpul asprglosis
C0948343|T047|AB|518.7|ICD9CM|Transfsn rel ac lung inj|Transfsn rel ac lung inj
C0948343|T047|PT|518.7|ICD9CM|Transfusion related acute lung injury (TRALI)|Transfusion related acute lung injury (TRALI)
C0348712|T047|HT|518.8|ICD9CM|Other diseases of lung|Other diseases of lung
C0264490|T047|PT|518.81|ICD9CM|Acute respiratory failure|Acute respiratory failure
C0264490|T047|AB|518.81|ICD9CM|Acute respiratry failure|Acute respiratry failure
C0302379|T047|AB|518.82|ICD9CM|Other pulmonary insuff|Other pulmonary insuff
C0302379|T047|PT|518.82|ICD9CM|Other pulmonary insufficiency, not elsewhere classified|Other pulmonary insufficiency, not elsewhere classified
C0264492|T047|AB|518.83|ICD9CM|Chronic respiratory fail|Chronic respiratory fail
C0264492|T047|PT|518.83|ICD9CM|Chronic respiratory failure|Chronic respiratory failure
C0264491|T047|AB|518.84|ICD9CM|Acute & chronc resp fail|Acute & chronc resp fail
C0264491|T047|PT|518.84|ICD9CM|Acute and chronic respiratory failure|Acute and chronic respiratory failure
C0029579|T047|PT|518.89|ICD9CM|Other diseases of lung, not elsewhere classified|Other diseases of lung, not elsewhere classified
C0029579|T047|AB|518.89|ICD9CM|Other lung disease NEC|Other lung disease NEC
C0029582|T047|HT|519|ICD9CM|Other diseases of respiratory system|Other diseases of respiratory system
C0155921|T046|HT|519.0|ICD9CM|Tracheostomy complications|Tracheostomy complications
C0155921|T046|AB|519.00|ICD9CM|Tracheostomy comp NOS|Tracheostomy comp NOS
C0155921|T046|PT|519.00|ICD9CM|Tracheostomy complication, unspecified|Tracheostomy complication, unspecified
C0695236|T047|PT|519.01|ICD9CM|Infection of tracheostomy|Infection of tracheostomy
C0695236|T047|AB|519.01|ICD9CM|Tracheostomy infection|Tracheostomy infection
C0695237|T046|PT|519.02|ICD9CM|Mechanical complication of tracheostomy|Mechanical complication of tracheostomy
C0695237|T046|AB|519.02|ICD9CM|Tracheostomy - mech comp|Tracheostomy - mech comp
C0695238|T046|PT|519.09|ICD9CM|Other tracheostomy complications|Other tracheostomy complications
C0695238|T046|AB|519.09|ICD9CM|Tracheostomy comp NEC|Tracheostomy comp NEC
C0869292|T047|HT|519.1|ICD9CM|Other diseases of trachea and bronchus, not elsewhere classified|Other diseases of trachea and bronchus, not elsewhere classified
C0741804|T047|PT|519.11|ICD9CM|Acute bronchospasm|Acute bronchospasm
C0741804|T047|AB|519.11|ICD9CM|Acute bronchospasm|Acute bronchospasm
C1719483|T047|PT|519.19|ICD9CM|Other diseases of trachea and bronchus|Other diseases of trachea and bronchus
C1719483|T047|AB|519.19|ICD9CM|Trachea & bronch dis NEC|Trachea & bronch dis NEC
C0025064|T047|AB|519.2|ICD9CM|Mediastinitis|Mediastinitis
C0025064|T047|PT|519.2|ICD9CM|Mediastinitis|Mediastinitis
C0869275|T047|AB|519.3|ICD9CM|Mediastinum disease NEC|Mediastinum disease NEC
C0869275|T047|PT|519.3|ICD9CM|Other diseases of mediastinum, not elsewhere classified|Other diseases of mediastinum, not elsewhere classified
C0152097|T047|AB|519.4|ICD9CM|Disorders of diaphragm|Disorders of diaphragm
C0152097|T047|PT|519.4|ICD9CM|Disorders of diaphragm|Disorders of diaphragm
C0869452|T047|PT|519.8|ICD9CM|Other diseases of respiratory system, not elsewhere classified|Other diseases of respiratory system, not elsewhere classified
C0869452|T047|AB|519.8|ICD9CM|Resp system disease NEC|Resp system disease NEC
C0035204|T047|AB|519.9|ICD9CM|Resp system disease NOS|Resp system disease NOS
C0035204|T047|PT|519.9|ICD9CM|Unspecified disease of respiratory system|Unspecified disease of respiratory system
C0155922|T047|HT|520|ICD9CM|Disorders of tooth development and eruption|Disorders of tooth development and eruption
C0348717|T047|HT|520-529.99|ICD9CM|DISEASES OF ORAL CAVITY, SALIVARY GLANDS, AND JAWS|DISEASES OF ORAL CAVITY, SALIVARY GLANDS, AND JAWS
C0012242|T047|HT|520-579.99|ICD9CM|DISEASES OF THE DIGESTIVE SYSTEM|DISEASES OF THE DIGESTIVE SYSTEM
C0399352|T019|AB|520.0|ICD9CM|Anodontia|Anodontia
C0399352|T019|PT|520.0|ICD9CM|Anodontia|Anodontia
C0040457|T033|AB|520.1|ICD9CM|Supernumerary teeth|Supernumerary teeth
C0040457|T033|PT|520.1|ICD9CM|Supernumerary teeth|Supernumerary teeth
C0000770|T190|AB|520.2|ICD9CM|Abnormal tooth size/form|Abnormal tooth size/form
C0000770|T190|PT|520.2|ICD9CM|Abnormalities of size and form of teeth|Abnormalities of size and form of teeth
C0026618|T047|AB|520.3|ICD9CM|Mottled teeth|Mottled teeth
C0026618|T047|PT|520.3|ICD9CM|Mottled teeth|Mottled teeth
C3495540|T047|PT|520.4|ICD9CM|Disturbances of tooth formation|Disturbances of tooth formation
C3495540|T047|AB|520.4|ICD9CM|Tooth formation disturb|Tooth formation disturb
C0868848|T019|AB|520.5|ICD9CM|Heredit tooth struct NEC|Heredit tooth struct NEC
C0868848|T019|PT|520.5|ICD9CM|Hereditary disturbances in tooth structure, not elsewhere classified|Hereditary disturbances in tooth structure, not elsewhere classified
C0012767|T047|PT|520.6|ICD9CM|Disturbances in tooth eruption|Disturbances in tooth eruption
C0012767|T047|AB|520.6|ICD9CM|Tooth eruption disturb|Tooth eruption disturb
C0039437|T033|AB|520.7|ICD9CM|Teething syndrome|Teething syndrome
C0039437|T033|PT|520.7|ICD9CM|Teething syndrome|Teething syndrome
C0155924|T047|PT|520.8|ICD9CM|Other specified disorders of tooth development and eruption|Other specified disorders of tooth development and eruption
C0155924|T047|AB|520.8|ICD9CM|Tooth devel/erup dis NEC|Tooth devel/erup dis NEC
C0155922|T047|AB|520.9|ICD9CM|Tooth devel/erup dis NOS|Tooth devel/erup dis NOS
C0155922|T047|PT|520.9|ICD9CM|Unspecified disorder of tooth development and eruption|Unspecified disorder of tooth development and eruption
C0155926|T047|HT|521|ICD9CM|Diseases of hard tissues of teeth|Diseases of hard tissues of teeth
C0011334|T047|HT|521.0|ICD9CM|Dental caries|Dental caries
C0011334|T047|AB|521.00|ICD9CM|Dental caries NOS|Dental caries NOS
C0011334|T047|PT|521.00|ICD9CM|Dental caries, unspecified|Dental caries, unspecified
C0266853|T047|AB|521.01|ICD9CM|Dental caries - enamel|Dental caries - enamel
C0266853|T047|PT|521.01|ICD9CM|Dental caries limited to enamel|Dental caries limited to enamel
C0266846|T047|AB|521.02|ICD9CM|Dental caries - dentine|Dental caries - dentine
C0266846|T047|PT|521.02|ICD9CM|Dental caries extending into dentine|Dental caries extending into dentine
C0399396|T047|AB|521.03|ICD9CM|Dental caries - pulp|Dental caries - pulp
C0399396|T047|PT|521.03|ICD9CM|Dental caries extending into pulp|Dental caries extending into pulp
C0266848|T047|PT|521.04|ICD9CM|Arrested dental caries|Arrested dental caries
C0266848|T047|AB|521.04|ICD9CM|Dental caries - arrested|Dental caries - arrested
C0341004|T047|AB|521.05|ICD9CM|Odontoclasia|Odontoclasia
C0341004|T047|PT|521.05|ICD9CM|Odontoclasia|Odontoclasia
C1456144|T047|PT|521.06|ICD9CM|Dental caries pit and fissure|Dental caries pit and fissure
C1456144|T047|AB|521.06|ICD9CM|Dentl caries-pit/fissure|Dentl caries-pit/fissure
C1456145|T047|PT|521.07|ICD9CM|Dental caries of smooth surface|Dental caries of smooth surface
C1456145|T047|AB|521.07|ICD9CM|Dentl caries-smooth surf|Dentl caries-smooth surf
C0162644|T047|PT|521.08|ICD9CM|Dental caries of root surface|Dental caries of root surface
C0162644|T047|AB|521.08|ICD9CM|Dental caries-root surf|Dental caries-root surf
C0348719|T047|AB|521.09|ICD9CM|Dental caries NEC|Dental caries NEC
C0348719|T047|PT|521.09|ICD9CM|Other dental caries|Other dental caries
C1456153|T047|HT|521.1|ICD9CM|Excessive dental attrition [approximal wear] [occlusal wear]|Excessive dental attrition [approximal wear] [occlusal wear]
C1456147|T047|AB|521.10|ICD9CM|Excessive attrition NOS|Excessive attrition NOS
C1456147|T047|PT|521.10|ICD9CM|Excessive attrition, unspecified|Excessive attrition, unspecified
C1456148|T047|AB|521.11|ICD9CM|Excess attrition-enamel|Excess attrition-enamel
C1456148|T047|PT|521.11|ICD9CM|Excessive attrition, limited to enamel|Excessive attrition, limited to enamel
C1456149|T047|AB|521.12|ICD9CM|Excess attrition-dentine|Excess attrition-dentine
C1456149|T047|PT|521.12|ICD9CM|Excessive attrition, extending into dentine|Excessive attrition, extending into dentine
C1456150|T047|AB|521.13|ICD9CM|Excessive attrition-pulp|Excessive attrition-pulp
C1456150|T047|PT|521.13|ICD9CM|Excessive attrition, extending into pulp|Excessive attrition, extending into pulp
C1456151|T047|AB|521.14|ICD9CM|Excess attrition-local|Excess attrition-local
C1456151|T047|PT|521.14|ICD9CM|Excessive attrition, localized|Excessive attrition, localized
C1456152|T047|AB|521.15|ICD9CM|Excess attrition-general|Excess attrition-general
C1456152|T047|PT|521.15|ICD9CM|Excessive attrition, generalized|Excessive attrition, generalized
C0040428|T046|HT|521.2|ICD9CM|Abrasion of teeth|Abrasion of teeth
C1302752|T037|AB|521.20|ICD9CM|Abrasion NOS|Abrasion NOS
C1302752|T037|PT|521.20|ICD9CM|Abrasion, unspecified|Abrasion, unspecified
C1456155|T047|AB|521.21|ICD9CM|Abrasion-enamel|Abrasion-enamel
C1456155|T047|PT|521.21|ICD9CM|Abrasion, limited to enamel|Abrasion, limited to enamel
C1456156|T047|AB|521.22|ICD9CM|Abrasion-dentine|Abrasion-dentine
C1456156|T047|PT|521.22|ICD9CM|Abrasion, extending into dentine|Abrasion, extending into dentine
C1456157|T047|AB|521.23|ICD9CM|Abrasion-pulp|Abrasion-pulp
C1456157|T047|PT|521.23|ICD9CM|Abrasion, extending into pulp|Abrasion, extending into pulp
C1456158|T047|AB|521.24|ICD9CM|Abrasion-localized|Abrasion-localized
C1456158|T047|PT|521.24|ICD9CM|Abrasion, localized|Abrasion, localized
C1456159|T047|AB|521.25|ICD9CM|Abrasion-generalized|Abrasion-generalized
C1456159|T047|PT|521.25|ICD9CM|Abrasion, generalized|Abrasion, generalized
C0040436|T047|HT|521.3|ICD9CM|Erosion of teeth|Erosion of teeth
C1456160|T047|AB|521.30|ICD9CM|Erosion NOS|Erosion NOS
C1456160|T047|PT|521.30|ICD9CM|Erosion, unspecified|Erosion, unspecified
C1456161|T047|AB|521.31|ICD9CM|Erosion-enamel|Erosion-enamel
C1456161|T047|PT|521.31|ICD9CM|Erosion, limited to enamel|Erosion, limited to enamel
C1456162|T047|AB|521.32|ICD9CM|Erosion-dentine|Erosion-dentine
C1456162|T047|PT|521.32|ICD9CM|Erosion, extending into dentine|Erosion, extending into dentine
C1456163|T047|AB|521.33|ICD9CM|Erosion-pulp|Erosion-pulp
C1456163|T047|PT|521.33|ICD9CM|Erosion, extending into pulp|Erosion, extending into pulp
C1456164|T047|AB|521.34|ICD9CM|Erosion-localized|Erosion-localized
C1456164|T047|PT|521.34|ICD9CM|Erosion, localized|Erosion, localized
C1456165|T047|AB|521.35|ICD9CM|Erosion-generalized|Erosion-generalized
C1456165|T047|PT|521.35|ICD9CM|Erosion, generalized|Erosion, generalized
C0040451|T047|HT|521.4|ICD9CM|Pathological tooth resorption|Pathological tooth resorption
C1456166|T047|AB|521.40|ICD9CM|Path resorption NOS|Path resorption NOS
C1456166|T047|PT|521.40|ICD9CM|Pathological resorption, unspecified|Pathological resorption, unspecified
C1456167|T047|AB|521.41|ICD9CM|Path resorption-internal|Path resorption-internal
C1456167|T047|PT|521.41|ICD9CM|Pathological resorption, internal|Pathological resorption, internal
C0266878|T047|AB|521.42|ICD9CM|Path resorption-external|Path resorption-external
C0266878|T047|PT|521.42|ICD9CM|Pathological resorption, external|Pathological resorption, external
C1456169|T047|PT|521.49|ICD9CM|Other pathological resorption|Other pathological resorption
C1456169|T047|AB|521.49|ICD9CM|Path resorption NEC|Path resorption NEC
C0020441|T047|AB|521.5|ICD9CM|Hypercementosis|Hypercementosis
C0020441|T047|PT|521.5|ICD9CM|Hypercementosis|Hypercementosis
C0155930|T047|AB|521.6|ICD9CM|Ankylosis of teeth|Ankylosis of teeth
C0155930|T047|PT|521.6|ICD9CM|Ankylosis of teeth|Ankylosis of teeth
C1456170|T047|AB|521.7|ICD9CM|Intrin posteruptv color|Intrin posteruptv color
C1456170|T047|PT|521.7|ICD9CM|Intrinsic posteruptive color changes|Intrinsic posteruptive color changes
C0029770|T047|HT|521.8|ICD9CM|Other specified diseases of hard tissues of teeth|Other specified diseases of hard tissues of teeth
C0010261|T033|PT|521.81|ICD9CM|Cracked tooth|Cracked tooth
C0010261|T033|AB|521.81|ICD9CM|Cracked tooth|Cracked tooth
C0029770|T047|AB|521.89|ICD9CM|Dis hard tiss teeth NEC|Dis hard tiss teeth NEC
C0029770|T047|PT|521.89|ICD9CM|Other specific diseases of hard tissues of teeth|Other specific diseases of hard tissues of teeth
C0155926|T047|AB|521.9|ICD9CM|Hard tiss dis teeth NOS|Hard tiss dis teeth NOS
C0155926|T047|PT|521.9|ICD9CM|Unspecified disease of hard tissues of teeth|Unspecified disease of hard tissues of teeth
C0155933|T047|HT|522|ICD9CM|Diseases of pulp and periapical tissues|Diseases of pulp and periapical tissues
C0034103|T047|AB|522.0|ICD9CM|Pulpitis|Pulpitis
C0034103|T047|PT|522.0|ICD9CM|Pulpitis|Pulpitis
C0011407|T047|PT|522.1|ICD9CM|Necrosis of the pulp|Necrosis of the pulp
C0011407|T047|AB|522.1|ICD9CM|Necrosis of tooth pulp|Necrosis of tooth pulp
C0034100|T047|PT|522.2|ICD9CM|Pulp degeneration|Pulp degeneration
C0034100|T047|AB|522.2|ICD9CM|Tooth pulp degeneration|Tooth pulp degeneration
C0399408|T047|AB|522.3|ICD9CM|Abn hard tiss-tooth pulp|Abn hard tiss-tooth pulp
C0399408|T047|PT|522.3|ICD9CM|Abnormal hard tissue formation in pulp|Abnormal hard tissue formation in pulp
C0155934|T047|AB|522.4|ICD9CM|Ac apical periodontitis|Ac apical periodontitis
C0155934|T047|PT|522.4|ICD9CM|Acute apical periodontitis of pulpal origin|Acute apical periodontitis of pulpal origin
C0399424|T047|AB|522.5|ICD9CM|Periapical abscess|Periapical abscess
C0399424|T047|PT|522.5|ICD9CM|Periapical abscess without sinus|Periapical abscess without sinus
C0392492|T047|AB|522.6|ICD9CM|Chr apical periodontitis|Chr apical periodontitis
C0392492|T047|PT|522.6|ICD9CM|Chronic apical periodontitis|Chronic apical periodontitis
C0266909|T047|AB|522.7|ICD9CM|Periapical absc w sinus|Periapical absc w sinus
C0266909|T047|PT|522.7|ICD9CM|Periapical abscess with sinus|Periapical abscess with sinus
C0034543|T047|AB|522.8|ICD9CM|Radicular cyst|Radicular cyst
C0034543|T047|PT|522.8|ICD9CM|Radicular cyst|Radicular cyst
C0155935|T047|PT|522.9|ICD9CM|Other and unspecified diseases of pulp and periapical tissues|Other and unspecified diseases of pulp and periapical tissues
C0155935|T047|AB|522.9|ICD9CM|Pulp/periapical dis NEC|Pulp/periapical dis NEC
C0155936|T047|HT|523|ICD9CM|Gingival and periodontal diseases|Gingival and periodontal diseases
C0155937|T047|HT|523.0|ICD9CM|Acute gingivitis|Acute gingivitis
C1719490|T047|AB|523.00|ICD9CM|Acute gingititis, plaque|Acute gingititis, plaque
C1719490|T047|PT|523.00|ICD9CM|Acute gingivitis, plaque induced|Acute gingivitis, plaque induced
C1719491|T047|AB|523.01|ICD9CM|Ac gingivitis,nonplaque|Ac gingivitis,nonplaque
C1719491|T047|PT|523.01|ICD9CM|Acute gingivitis, non-plaque induced|Acute gingivitis, non-plaque induced
C0008684|T047|HT|523.1|ICD9CM|Chronic gingivitis|Chronic gingivitis
C1719717|T047|AB|523.10|ICD9CM|Chronc gingititis,plaque|Chronc gingititis,plaque
C1719717|T047|PT|523.10|ICD9CM|Chronic gingivitis, plaque induced|Chronic gingivitis, plaque induced
C1719492|T047|AB|523.11|ICD9CM|Chr gingivitis-nonplaque|Chr gingivitis-nonplaque
C1719492|T047|PT|523.11|ICD9CM|Chronic gingivitis, non-plaque induced|Chronic gingivitis, non-plaque induced
C0017572|T047|HT|523.2|ICD9CM|Gingival recession|Gingival recession
C0017572|T047|AB|523.20|ICD9CM|Gingival recession NOS|Gingival recession NOS
C0017572|T047|PT|523.20|ICD9CM|Gingival recession, unspecified|Gingival recession, unspecified
C1456171|T047|AB|523.21|ICD9CM|Gingival recess-minimal|Gingival recess-minimal
C1456171|T047|PT|523.21|ICD9CM|Gingival recession, minimal|Gingival recession, minimal
C1456172|T047|AB|523.22|ICD9CM|Gingival recess-moderate|Gingival recess-moderate
C1456172|T047|PT|523.22|ICD9CM|Gingival recession, moderate|Gingival recession, moderate
C1456173|T047|AB|523.23|ICD9CM|Gingival recess-severe|Gingival recess-severe
C1456173|T047|PT|523.23|ICD9CM|Gingival recession, severe|Gingival recession, severe
C0266916|T047|AB|523.24|ICD9CM|Gingival recession-local|Gingival recession-local
C0266916|T047|PT|523.24|ICD9CM|Gingival recession, localized|Gingival recession, localized
C0266915|T047|AB|523.25|ICD9CM|Gingival recess-general|Gingival recess-general
C0266915|T047|PT|523.25|ICD9CM|Gingival recession, generalized|Gingival recession, generalized
C0001342|T047|HT|523.3|ICD9CM|Aggressive and acute periodontitis|Aggressive and acute periodontitis
C1719493|T047|AB|523.30|ICD9CM|Aggres periodontitis NOS|Aggres periodontitis NOS
C1719493|T047|PT|523.30|ICD9CM|Aggressive periodontitis, unspecified|Aggressive periodontitis, unspecified
C1719494|T047|AB|523.31|ICD9CM|Aggres periodontitis,loc|Aggres periodontitis,loc
C1719494|T047|PT|523.31|ICD9CM|Aggressive periodontitis, localized|Aggressive periodontitis, localized
C1719495|T047|AB|523.32|ICD9CM|Aggres periodontitis,gen|Aggres periodontitis,gen
C1719495|T047|PT|523.32|ICD9CM|Aggressive periodontitis, generalized|Aggressive periodontitis, generalized
C0001342|T047|PT|523.33|ICD9CM|Acute periodontitis|Acute periodontitis
C0001342|T047|AB|523.33|ICD9CM|Acute periodontitis|Acute periodontitis
C0266929|T047|HT|523.4|ICD9CM|Chronic periodontitis|Chronic periodontitis
C0266929|T047|AB|523.40|ICD9CM|Chronc periodontitis NOS|Chronc periodontitis NOS
C0266929|T047|PT|523.40|ICD9CM|Chronic periodontitis, unspecified|Chronic periodontitis, unspecified
C1719497|T047|AB|523.41|ICD9CM|Chr periodontitis, local|Chr periodontitis, local
C1719497|T047|PT|523.41|ICD9CM|Chronic periodontitis, localized|Chronic periodontitis, localized
C1719498|T047|AB|523.42|ICD9CM|Chron periodontitis,gen|Chron periodontitis,gen
C1719498|T047|PT|523.42|ICD9CM|Chronic periodontitis, generalized|Chronic periodontitis, generalized
C0600298|T047|AB|523.5|ICD9CM|Periodontosis|Periodontosis
C0600298|T047|PT|523.5|ICD9CM|Periodontosis|Periodontosis
C0011346|T047|AB|523.6|ICD9CM|Accretions on teeth|Accretions on teeth
C0011346|T047|PT|523.6|ICD9CM|Accretions on teeth|Accretions on teeth
C0029821|T047|PT|523.8|ICD9CM|Other specified periodontal diseases|Other specified periodontal diseases
C0029821|T047|AB|523.8|ICD9CM|Periodontal disease NEC|Periodontal disease NEC
C0155936|T047|AB|523.9|ICD9CM|Gingiv/periodont dis NOS|Gingiv/periodont dis NOS
C0155936|T047|PT|523.9|ICD9CM|Unspecified gingival and periodontal disease|Unspecified gingival and periodontal disease
C0155938|T019|HT|524|ICD9CM|Dentofacial anomalies, including malocclusion|Dentofacial anomalies, including malocclusion
C0024508|T019|HT|524.0|ICD9CM|Major anomalies of jaw size|Major anomalies of jaw size
C0024508|T019|PT|524.00|ICD9CM|Major anomalies of jaw size, unspecified anomaly|Major anomalies of jaw size, unspecified anomaly
C0024508|T019|AB|524.00|ICD9CM|Unspcf anomaly jaw size|Unspcf anomaly jaw size
C2227090|T033|PT|524.01|ICD9CM|Major anomalies of jaw size, maxillary hyperplasia|Major anomalies of jaw size, maxillary hyperplasia
C2227090|T033|AB|524.01|ICD9CM|Maxillary hyperplasia|Maxillary hyperplasia
C0302501|T190|PT|524.02|ICD9CM|Major anomalies of jaw size, mandibular hyperplasia|Major anomalies of jaw size, mandibular hyperplasia
C0302501|T190|AB|524.02|ICD9CM|Mandibular hyperplasia|Mandibular hyperplasia
C0240310|T019|PT|524.03|ICD9CM|Major anomalies of jaw size, maxillary hypoplasia|Major anomalies of jaw size, maxillary hypoplasia
C0240310|T019|AB|524.03|ICD9CM|Maxillary hypoplasia|Maxillary hypoplasia
C4024589|T190|PT|524.04|ICD9CM|Major anomalies of jaw size, mandibular hypoplasia|Major anomalies of jaw size, mandibular hypoplasia
C4024589|T190|AB|524.04|ICD9CM|Mandibular hypoplasia|Mandibular hypoplasia
C0341029|T190|AB|524.05|ICD9CM|Macrogenia|Macrogenia
C0341029|T190|PT|524.05|ICD9CM|Major anomalies of jaw size, macrogenia|Major anomalies of jaw size, macrogenia
C0341030|T190|PT|524.06|ICD9CM|Major anomalies of jaw size, microgenia|Major anomalies of jaw size, microgenia
C0341030|T190|AB|524.06|ICD9CM|Microgenia|Microgenia
C1456175|T047|PT|524.07|ICD9CM|Excessive tuberosity of jaw|Excessive tuberosity of jaw
C1456175|T047|AB|524.07|ICD9CM|Excessive tuberosity-jaw|Excessive tuberosity-jaw
C0375340|T019|PT|524.09|ICD9CM|Major anomalies of jaw size, other specified anomaly|Major anomalies of jaw size, other specified anomaly
C0375340|T019|AB|524.09|ICD9CM|Oth spcf anmly jaw size|Oth spcf anmly jaw size
C0003110|T190|HT|524.1|ICD9CM|Anomalies of relationship of jaw to cranial base|Anomalies of relationship of jaw to cranial base
C0003110|T190|PT|524.10|ICD9CM|Anomalies of relationship of jaw to cranial base, unspecified anomaly|Anomalies of relationship of jaw to cranial base, unspecified anomaly
C0003110|T190|AB|524.10|ICD9CM|Unspcf anm jaw cranl bse|Unspcf anm jaw cranl bse
C0399519|T033|PT|524.11|ICD9CM|Anomalies of relationship of jaw to cranial base, maxillary asymmetry|Anomalies of relationship of jaw to cranial base, maxillary asymmetry
C0399519|T033|AB|524.11|ICD9CM|Maxillary asymmetry|Maxillary asymmetry
C0375343|T190|PT|524.12|ICD9CM|Anomalies of relationship of jaw to cranial base, other jaw asymmetry|Anomalies of relationship of jaw to cranial base, other jaw asymmetry
C0375343|T190|AB|524.12|ICD9CM|Other jaw asymmetry|Other jaw asymmetry
C0375344|T190|PT|524.19|ICD9CM|Anomalies of relationship of jaw to cranial base, other specified anomaly|Anomalies of relationship of jaw to cranial base, other specified anomaly
C0375344|T190|AB|524.19|ICD9CM|Spcfd anom jaw cranl bse|Spcfd anom jaw cranl bse
C0155939|T190|HT|524.2|ICD9CM|Anomalies of dental arch relationship|Anomalies of dental arch relationship
C0155939|T190|AB|524.20|ICD9CM|Anomaly dental arch NOS|Anomaly dental arch NOS
C0155939|T190|PT|524.20|ICD9CM|Unspecified anomaly of dental arch relationship|Unspecified anomaly of dental arch relationship
C0399523|T047|AB|524.21|ICD9CM|Malocc- Angle's class I|Malocc- Angle's class I
C0399523|T047|PT|524.21|ICD9CM|Malocclusion, Angle's class I|Malocclusion, Angle's class I
C3714535|T190|AB|524.22|ICD9CM|Malocc-Angle's class II|Malocc-Angle's class II
C3714535|T190|PT|524.22|ICD9CM|Malocclusion, Angle's class II|Malocclusion, Angle's class II
C0399526|T019|AB|524.23|ICD9CM|Malocc-Angle's class III|Malocc-Angle's class III
C0399526|T019|PT|524.23|ICD9CM|Malocclusion, Angle's class III|Malocclusion, Angle's class III
C1456180|T033|PT|524.24|ICD9CM|Open anterior occlusal relationship|Open anterior occlusal relationship
C1456180|T033|AB|524.24|ICD9CM|Open anterior occlusion|Open anterior occlusion
C1456181|T033|PT|524.25|ICD9CM|Open posterior occlusal relationship|Open posterior occlusal relationship
C1456181|T033|AB|524.25|ICD9CM|Open posterior occlusion|Open posterior occlusion
C1456182|T047|AB|524.26|ICD9CM|Excess horizontl overlap|Excess horizontl overlap
C1456182|T047|PT|524.26|ICD9CM|Excessive horizontal overlap|Excessive horizontal overlap
C1456183|T047|AB|524.27|ICD9CM|Reverse articulation|Reverse articulation
C1456183|T190|AB|524.27|ICD9CM|Reverse articulation|Reverse articulation
C1456183|T047|PT|524.27|ICD9CM|Reverse articulation|Reverse articulation
C1456183|T190|PT|524.27|ICD9CM|Reverse articulation|Reverse articulation
C1456186|T047|AB|524.28|ICD9CM|Anom interarch distance|Anom interarch distance
C1456186|T047|PT|524.28|ICD9CM|Anomalies of interarch distance|Anomalies of interarch distance
C1456189|T047|AB|524.29|ICD9CM|Anomaly dental arch NEC|Anomaly dental arch NEC
C1456189|T047|PT|524.29|ICD9CM|Other anomalies of dental arch relationship|Other anomalies of dental arch relationship
C1456201|T190|HT|524.3|ICD9CM|Anomalies of tooth position of fully erupted teeth|Anomalies of tooth position of fully erupted teeth
C0155940|T190|AB|524.30|ICD9CM|Tooth position anom NOS|Tooth position anom NOS
C0155940|T190|PT|524.30|ICD9CM|Unspecified anomaly of tooth position|Unspecified anomaly of tooth position
C0040433|T033|AB|524.31|ICD9CM|Crowding of teeth|Crowding of teeth
C0040433|T033|PT|524.31|ICD9CM|Crowding of teeth|Crowding of teeth
C1456191|T047|PT|524.32|ICD9CM|Excessive spacing of teeth|Excessive spacing of teeth
C1456191|T047|AB|524.32|ICD9CM|Excessive spacing-teeth|Excessive spacing-teeth
C1456192|T190|PT|524.33|ICD9CM|Horizontal displacement of teeth|Horizontal displacement of teeth
C1456192|T190|AB|524.33|ICD9CM|Horizontl displace-teeth|Horizontl displace-teeth
C1456194|T190|AB|524.34|ICD9CM|Vertical displace-teeth|Vertical displace-teeth
C1456194|T190|PT|524.34|ICD9CM|Vertical displacement of teeth|Vertical displacement of teeth
C0266071|T019|AB|524.35|ICD9CM|Rotation of teeth|Rotation of teeth
C0266071|T019|PT|524.35|ICD9CM|Rotation of tooth/teeth|Rotation of tooth/teeth
C1456197|T047|AB|524.36|ICD9CM|Insuf interocclusl-teeth|Insuf interocclusl-teeth
C1456197|T047|PT|524.36|ICD9CM|Insufficient interocclusal distance of teeth (ridge)|Insufficient interocclusal distance of teeth (ridge)
C1456198|T190|AB|524.37|ICD9CM|Exces interocclusl-teeth|Exces interocclusl-teeth
C1456198|T190|PT|524.37|ICD9CM|Excessive interocclusal distance of teeth|Excessive interocclusal distance of teeth
C1456200|T047|PT|524.39|ICD9CM|Other anomalies of tooth position|Other anomalies of tooth position
C1456200|T047|AB|524.39|ICD9CM|Tooth position anom NEC|Tooth position anom NEC
C0024636|T190|AB|524.4|ICD9CM|Malocclusion NOS|Malocclusion NOS
C0024636|T190|PT|524.4|ICD9CM|Malocclusion, unspecified|Malocclusion, unspecified
C0266932|T190|HT|524.5|ICD9CM|Dentofacial functional abnormalities|Dentofacial functional abnormalities
C0266932|T190|AB|524.50|ICD9CM|Dentofac funct abnor NOS|Dentofac funct abnor NOS
C0266932|T190|PT|524.50|ICD9CM|Dentofacial functional abnormality, unspecified|Dentofacial functional abnormality, unspecified
C0266933|T047|AB|524.51|ICD9CM|Abnormal jaw closure|Abnormal jaw closure
C0266933|T047|PT|524.51|ICD9CM|Abnormal jaw closure|Abnormal jaw closure
C0521590|T033|PT|524.52|ICD9CM|Limited mandibular range of motion|Limited mandibular range of motion
C0521590|T033|AB|524.52|ICD9CM|Limited mandibular ROM|Limited mandibular ROM
C1456203|T047|AB|524.53|ICD9CM|Dev open/close mandible|Dev open/close mandible
C1456203|T047|PT|524.53|ICD9CM|Deviation in opening and closing of the mandible|Deviation in opening and closing of the mandible
C1291056|T190|AB|524.54|ICD9CM|Insuff anterior guidance|Insuff anterior guidance
C1291056|T190|PT|524.54|ICD9CM|Insufficient anterior guidance|Insufficient anterior guidance
C1456205|T047|AB|524.55|ICD9CM|Centric occl intrcsp dis|Centric occl intrcsp dis
C1456205|T047|PT|524.55|ICD9CM|Centric occlusion maximum intercuspation discrepancy|Centric occlusion maximum intercuspation discrepancy
C2895155|T190|PT|524.56|ICD9CM|Non-working side interference|Non-working side interference
C2895155|T190|AB|524.56|ICD9CM|Nonwork side interfrnce|Nonwork side interfrnce
C1456207|T033|PT|524.57|ICD9CM|Lack of posterior occlusal support|Lack of posterior occlusal support
C1456207|T033|AB|524.57|ICD9CM|Lack post occlsl support|Lack post occlsl support
C1456208|T047|AB|524.59|ICD9CM|Dentofac funct abnor NEC|Dentofac funct abnor NEC
C1456208|T047|PT|524.59|ICD9CM|Other dentofacial functional abnormalities|Other dentofacial functional abnormalities
C0039494|T047|HT|524.6|ICD9CM|Temporomandibular joint disorders|Temporomandibular joint disorders
C0039494|T047|PT|524.60|ICD9CM|Temporomandibular joint disorders, unspecified|Temporomandibular joint disorders, unspecified
C0039494|T047|AB|524.60|ICD9CM|TMJ disorders NOS|TMJ disorders NOS
C0155942|T047|AB|524.61|ICD9CM|Adhesns/ankylosis - TMJ|Adhesns/ankylosis - TMJ
C0155942|T047|PT|524.61|ICD9CM|Temporomandibular joint disorders, adhesions and ankylosis (bony or fibrous)|Temporomandibular joint disorders, adhesions and ankylosis (bony or fibrous)
C0155943|T047|AB|524.62|ICD9CM|Arthralgia TMJ|Arthralgia TMJ
C0155943|T047|PT|524.62|ICD9CM|Temporomandibular joint disorders, arthralgia of temporomandibular joint|Temporomandibular joint disorders, arthralgia of temporomandibular joint
C0685925|T047|AB|524.63|ICD9CM|Articular disc disorder|Articular disc disorder
C0685925|T047|PT|524.63|ICD9CM|Temporomandibular joint disorders, articular disc disorder (reducing or non-reducing)|Temporomandibular joint disorders, articular disc disorder (reducing or non-reducing)
C1456213|T047|PT|524.64|ICD9CM|Temporomandibular joint sounds on opening and/or closing the jaw|Temporomandibular joint sounds on opening and/or closing the jaw
C1456213|T047|AB|524.64|ICD9CM|TMJ sounds opn/close jaw|TMJ sounds opn/close jaw
C0155945|T047|AB|524.69|ICD9CM|Other specf TMJ disordrs|Other specf TMJ disordrs
C0155945|T047|PT|524.69|ICD9CM|Other specified temporomandibular joint disorders|Other specified temporomandibular joint disorders
C0375346|T190|HT|524.7|ICD9CM|Dental alveolar anomalies|Dental alveolar anomalies
C0375346|T190|PT|524.70|ICD9CM|Dental alveolar anomalies, unspecified alveolar anomaly|Dental alveolar anomalies, unspecified alveolar anomaly
C0375346|T190|AB|524.70|ICD9CM|Unspf dent alvelr anmaly|Unspf dent alvelr anmaly
C0375347|T190|AB|524.71|ICD9CM|Alveolar maxil hyprplsia|Alveolar maxil hyprplsia
C0375347|T190|PT|524.71|ICD9CM|Alveolar maxillary hyperplasia|Alveolar maxillary hyperplasia
C0375348|T190|AB|524.72|ICD9CM|Alveolar mandib hyprplas|Alveolar mandib hyprplas
C0375348|T190|PT|524.72|ICD9CM|Alveolar mandibular hyperplasia|Alveolar mandibular hyperplasia
C0375349|T190|AB|524.73|ICD9CM|Alveolar maxil hypoplsia|Alveolar maxil hypoplsia
C0375349|T190|PT|524.73|ICD9CM|Alveolar maxillary hypoplasia|Alveolar maxillary hypoplasia
C0375350|T190|AB|524.74|ICD9CM|Alveolar mandb hypoplsia|Alveolar mandb hypoplsia
C0375350|T190|PT|524.74|ICD9CM|Alveolar mandibular hypoplasia|Alveolar mandibular hypoplasia
C1456214|T047|AB|524.75|ICD9CM|Vertical displace teeth|Vertical displace teeth
C1456214|T047|PT|524.75|ICD9CM|Vertical displacement of alveolus and teeth|Vertical displacement of alveolus and teeth
C1456216|T033|AB|524.76|ICD9CM|Occlusal plane deviation|Occlusal plane deviation
C1456216|T033|PT|524.76|ICD9CM|Occlusal plane deviation|Occlusal plane deviation
C0859118|T190|AB|524.79|ICD9CM|Oth spcf alveolar anmaly|Oth spcf alveolar anmaly
C0859118|T190|PT|524.79|ICD9CM|Other specified alveolar anomaly|Other specified alveolar anomaly
C0155946|T047|HT|524.8|ICD9CM|Other specified dentofacial anomalies|Other specified dentofacial anomalies
C1456217|T047|AB|524.81|ICD9CM|Anterior soft tiss impg|Anterior soft tiss impg
C1456217|T047|PT|524.81|ICD9CM|Anterior soft tissue impingement|Anterior soft tissue impingement
C1456218|T047|AB|524.82|ICD9CM|Posterior soft tiss impg|Posterior soft tiss impg
C1456218|T047|PT|524.82|ICD9CM|Posterior soft tissue impingement|Posterior soft tissue impingement
C0155946|T047|AB|524.89|ICD9CM|Dentofacial anomaly NEC|Dentofacial anomaly NEC
C0155946|T047|PT|524.89|ICD9CM|Other specified dentofacial anomalies|Other specified dentofacial anomalies
C0155947|T190|AB|524.9|ICD9CM|Dentofacial anomaly NOS|Dentofacial anomaly NOS
C0155947|T190|PT|524.9|ICD9CM|Unspecified dentofacial anomalies|Unspecified dentofacial anomalies
C0155948|T047|HT|525|ICD9CM|Other diseases and conditions of the teeth and supporting structures|Other diseases and conditions of the teeth and supporting structures
C0155949|T047|AB|525.0|ICD9CM|Exfoliation of teeth|Exfoliation of teeth
C0155949|T047|PT|525.0|ICD9CM|Exfoliation of teeth due to systemic causes|Exfoliation of teeth due to systemic causes
C1168590|T047|HT|525.1|ICD9CM|Loss of teeth due to trauma, extraction, or periodontal disease|Loss of teeth due to trauma, extraction, or periodontal disease
C0080233|T020|AB|525.10|ICD9CM|Acq absence of teeth NOS|Acq absence of teeth NOS
C0080233|T020|PT|525.10|ICD9CM|Acquired absence of teeth, unspecified|Acquired absence of teeth, unspecified
C0949130|T047|AB|525.11|ICD9CM|Loss of teeth d/t trauma|Loss of teeth d/t trauma
C0949130|T047|PT|525.11|ICD9CM|Loss of teeth due to trauma|Loss of teeth due to trauma
C0949131|T047|PT|525.12|ICD9CM|Loss of teeth due to periodontal disease|Loss of teeth due to periodontal disease
C0949131|T047|AB|525.12|ICD9CM|Loss teeth d/t peri dis|Loss teeth d/t peri dis
C0949132|T047|AB|525.13|ICD9CM|Loss of teeth d/t caries|Loss of teeth d/t caries
C0949132|T047|PT|525.13|ICD9CM|Loss of teeth due to caries|Loss of teeth due to caries
C0949133|T047|AB|525.19|ICD9CM|Loss of teeth NEC|Loss of teeth NEC
C0949133|T047|PT|525.19|ICD9CM|Other loss of teeth|Other loss of teeth
C0155951|T047|HT|525.2|ICD9CM|Atrophy of edentulous alveolar ridge|Atrophy of edentulous alveolar ridge
C1456219|T047|AB|525.20|ICD9CM|Atrophy alvlar ridge NOS|Atrophy alvlar ridge NOS
C1456219|T047|PT|525.20|ICD9CM|Unspecified atrophy of edentulous alveolar ridge|Unspecified atrophy of edentulous alveolar ridge
C1456221|T047|AB|525.21|ICD9CM|Atrophy mandible-minimal|Atrophy mandible-minimal
C1456221|T047|PT|525.21|ICD9CM|Minimal atrophy of the mandible|Minimal atrophy of the mandible
C1456222|T047|AB|525.22|ICD9CM|Atrophy mandible-modrate|Atrophy mandible-modrate
C1456222|T047|PT|525.22|ICD9CM|Moderate atrophy of the mandible|Moderate atrophy of the mandible
C1456223|T047|AB|525.23|ICD9CM|Atrophy mandible-severe|Atrophy mandible-severe
C1456223|T047|PT|525.23|ICD9CM|Severe atrophy of the mandible|Severe atrophy of the mandible
C1456224|T047|AB|525.24|ICD9CM|Atrophy maxilla-minimal|Atrophy maxilla-minimal
C1456224|T047|PT|525.24|ICD9CM|Minimal atrophy of the maxilla|Minimal atrophy of the maxilla
C1456225|T047|AB|525.25|ICD9CM|Atrophy maxilla-moderate|Atrophy maxilla-moderate
C1456225|T047|PT|525.25|ICD9CM|Moderate atrophy of the maxilla|Moderate atrophy of the maxilla
C1456226|T047|AB|525.26|ICD9CM|Atrophy maxilla-severe|Atrophy maxilla-severe
C1456226|T047|PT|525.26|ICD9CM|Severe atrophy of the maxilla|Severe atrophy of the maxilla
C0155952|T047|AB|525.3|ICD9CM|Retained dental root|Retained dental root
C0155952|T047|PT|525.3|ICD9CM|Retained dental root|Retained dental root
C1561613|T047|HT|525.4|ICD9CM|Complete edentulism|Complete edentulism
C1561613|T047|AB|525.40|ICD9CM|Complete edentulism NOS|Complete edentulism NOS
C1561613|T047|PT|525.40|ICD9CM|Complete edentulism, unspecified|Complete edentulism, unspecified
C1561614|T047|AB|525.41|ICD9CM|Comp edentulism,class I|Comp edentulism,class I
C1561614|T047|PT|525.41|ICD9CM|Complete edentulism, class I|Complete edentulism, class I
C1561615|T047|AB|525.42|ICD9CM|Comp edentulism,class II|Comp edentulism,class II
C1561615|T047|PT|525.42|ICD9CM|Complete edentulism, class II|Complete edentulism, class II
C1561616|T047|AB|525.43|ICD9CM|Comp edentulsm,class III|Comp edentulsm,class III
C1561616|T047|PT|525.43|ICD9CM|Complete edentulism, class III|Complete edentulism, class III
C1561617|T047|AB|525.44|ICD9CM|Comp edentulism,class IV|Comp edentulism,class IV
C1561617|T047|PT|525.44|ICD9CM|Complete edentulism, class IV|Complete edentulism, class IV
C1561619|T047|HT|525.5|ICD9CM|Partial edentulism|Partial edentulism
C1561619|T047|AB|525.50|ICD9CM|Partial edentulism NOS|Partial edentulism NOS
C1561619|T047|PT|525.50|ICD9CM|Partial edentulism, unspecified|Partial edentulism, unspecified
C1561620|T047|AB|525.51|ICD9CM|Part edentulism,class I|Part edentulism,class I
C1561620|T047|PT|525.51|ICD9CM|Partial edentulism, class I|Partial edentulism, class I
C1561621|T047|AB|525.52|ICD9CM|Part edentulism,class II|Part edentulism,class II
C1561621|T047|PT|525.52|ICD9CM|Partial edentulism, class II|Partial edentulism, class II
C1561622|T047|AB|525.53|ICD9CM|Part edentulsm,class III|Part edentulsm,class III
C1561622|T047|PT|525.53|ICD9CM|Partial edentulism, class III|Partial edentulism, class III
C1561623|T047|AB|525.54|ICD9CM|Part edentulism,class IV|Part edentulism,class IV
C1561623|T047|PT|525.54|ICD9CM|Partial edentulism, class IV|Partial edentulism, class IV
C1719519|T033|HT|525.6|ICD9CM|Unsatisfactory restoration of tooth|Unsatisfactory restoration of tooth
C1719507|T033|AB|525.60|ICD9CM|Unsat restore tooth NOS|Unsat restore tooth NOS
C1719507|T033|PT|525.60|ICD9CM|Unspecified unsatisfactory restoration of tooth|Unspecified unsatisfactory restoration of tooth
C1290744|T047|AB|525.61|ICD9CM|Open restoration margins|Open restoration margins
C1290744|T047|PT|525.61|ICD9CM|Open restoration margins|Open restoration margins
C2188200|T047|AB|525.62|ICD9CM|Overhang dental restore|Overhang dental restore
C2188200|T047|PT|525.62|ICD9CM|Unrepairable overhanging of dental restorative materials|Unrepairable overhanging of dental restorative materials
C1719512|T047|PT|525.63|ICD9CM|Fractured dental restorative material without loss of material|Fractured dental restorative material without loss of material
C1719512|T047|AB|525.63|ICD9CM|Fx dental mat w/o loss|Fx dental mat w/o loss
C1719513|T046|PT|525.64|ICD9CM|Fractured dental restorative material with loss of material|Fractured dental restorative material with loss of material
C1719513|T046|AB|525.64|ICD9CM|Fx dentl material w loss|Fx dentl material w loss
C1719514|T047|PT|525.65|ICD9CM|Contour of existing restoration of tooth biologically incompatible with oral health|Contour of existing restoration of tooth biologically incompatible with oral health
C1719514|T047|AB|525.65|ICD9CM|Contour restore tooth|Contour restore tooth
C1719719|T046|AB|525.66|ICD9CM|Allergy dental res mat|Allergy dental res mat
C1719719|T046|PT|525.66|ICD9CM|Allergy to existing dental restorative material|Allergy to existing dental restorative material
C1719517|T046|PT|525.67|ICD9CM|Poor aesthetics of existing restoration|Poor aesthetics of existing restoration
C1719517|T046|AB|525.67|ICD9CM|Poor aesthetics restore|Poor aesthetics restore
C1719518|T033|PT|525.69|ICD9CM|Other unsatisfactory restoration of existing tooth|Other unsatisfactory restoration of existing tooth
C1719518|T033|AB|525.69|ICD9CM|Unsat restore tooth NEC|Unsat restore tooth NEC
C1955812|T046|HT|525.7|ICD9CM|Endosseous dental implant failure|Endosseous dental implant failure
C2711774|T046|AB|525.71|ICD9CM|Osseo fail dental implnt|Osseo fail dental implnt
C2711774|T046|PT|525.71|ICD9CM|Osseointegration failure of dental implant|Osseointegration failure of dental implant
C1955799|T046|AB|525.72|ICD9CM|Post-osse biol fail impl|Post-osse biol fail impl
C1955799|T046|PT|525.72|ICD9CM|Post-osseointegration biological failure of dental implant|Post-osseointegration biological failure of dental implant
C1955807|T046|AB|525.73|ICD9CM|Post-osse mech fail impl|Post-osse mech fail impl
C1955807|T046|PT|525.73|ICD9CM|Post-osseointegration mechanical failure of dental implant|Post-osseointegration mechanical failure of dental implant
C1955810|T047|AB|525.79|ICD9CM|Endos dentl imp fail NEC|Endos dentl imp fail NEC
C1955810|T047|PT|525.79|ICD9CM|Other endosseous dental implant failure|Other endosseous dental implant failure
C0029790|T047|AB|525.8|ICD9CM|Dental disorder NEC|Dental disorder NEC
C0029790|T047|PT|525.8|ICD9CM|Other specified disorders of the teeth and supporting structures|Other specified disorders of the teeth and supporting structures
C1704330|T047|AB|525.9|ICD9CM|Dental disorder NOS|Dental disorder NOS
C1704330|T047|PT|525.9|ICD9CM|Unspecified disorder of the teeth and supporting structures|Unspecified disorder of the teeth and supporting structures
C0022362|T047|HT|526|ICD9CM|Diseases of the jaws|Diseases of the jaws
C2939144|T047|AB|526.0|ICD9CM|Devel odontogenic cysts|Devel odontogenic cysts
C2939144|T047|PT|526.0|ICD9CM|Developmental odontogenic cysts|Developmental odontogenic cysts
C0341039|T047|AB|526.1|ICD9CM|Fissural cysts of jaw|Fissural cysts of jaw
C0341039|T047|PT|526.1|ICD9CM|Fissural cysts of jaw|Fissural cysts of jaw
C0029569|T047|AB|526.2|ICD9CM|Cysts of jaws NEC|Cysts of jaws NEC
C0029569|T047|PT|526.2|ICD9CM|Other cysts of jaws|Other cysts of jaws
C0162375|T047|AB|526.3|ICD9CM|Cent giant cell granulom|Cent giant cell granulom
C0162375|T047|PT|526.3|ICD9CM|Central giant cell (reparative) granuloma|Central giant cell (reparative) granuloma
C0155954|T047|AB|526.4|ICD9CM|Inflammation of jaw|Inflammation of jaw
C0155954|T047|PT|526.4|ICD9CM|Inflammatory conditions of jaw|Inflammatory conditions of jaw
C0013240|T047|AB|526.5|ICD9CM|Alveolitis of jaw|Alveolitis of jaw
C0013240|T047|PT|526.5|ICD9CM|Alveolitis of jaw|Alveolitis of jaw
C1719524|T046|HT|526.6|ICD9CM|Periradicular pathology associated with previous endodontic treatment|Periradicular pathology associated with previous endodontic treatment
C1719521|T046|AB|526.61|ICD9CM|Perfor root canal space|Perfor root canal space
C1719521|T046|PT|526.61|ICD9CM|Perforation of root canal space|Perforation of root canal space
C1719522|T047|PT|526.62|ICD9CM|Endodontic overfill|Endodontic overfill
C1719522|T047|AB|526.62|ICD9CM|Endodontic overfill|Endodontic overfill
C1719523|T047|PT|526.63|ICD9CM|Endodontic underfill|Endodontic underfill
C1719523|T047|AB|526.63|ICD9CM|Endodontic underfill|Endodontic underfill
C1719713|T046|PT|526.69|ICD9CM|Other periradicular pathology associated with previous endodontic treatment|Other periradicular pathology associated with previous endodontic treatment
C1719713|T046|AB|526.69|ICD9CM|Periradicular path NEC|Periradicular path NEC
C0029772|T047|HT|526.8|ICD9CM|Other specified diseases of the jaws|Other specified diseases of the jaws
C0155955|T047|AB|526.81|ICD9CM|Exostosis of jaw|Exostosis of jaw
C0155955|T047|PT|526.81|ICD9CM|Exostosis of jaw|Exostosis of jaw
C0029772|T047|AB|526.89|ICD9CM|Jaw disease NEC|Jaw disease NEC
C0029772|T047|PT|526.89|ICD9CM|Other specified diseases of the jaws|Other specified diseases of the jaws
C0022362|T047|AB|526.9|ICD9CM|Jaw disease NOS|Jaw disease NOS
C0022362|T047|PT|526.9|ICD9CM|Unspecified disease of the jaws|Unspecified disease of the jaws
C0036093|T047|HT|527|ICD9CM|Diseases of the salivary glands|Diseases of the salivary glands
C0155956|T020|PT|527.0|ICD9CM|Atrophy of salivary gland|Atrophy of salivary gland
C0155956|T020|AB|527.0|ICD9CM|Salivary gland atrophy|Salivary gland atrophy
C0020569|T046|PT|527.1|ICD9CM|Hypertrophy of salivary gland|Hypertrophy of salivary gland
C0020569|T046|AB|527.1|ICD9CM|Salivary glnd hyprtrophy|Salivary glnd hyprtrophy
C0037023|T047|AB|527.2|ICD9CM|Sialoadenitis|Sialoadenitis
C0037023|T047|PT|527.2|ICD9CM|Sialoadenitis|Sialoadenitis
C0155957|T047|PT|527.3|ICD9CM|Abscess of salivary gland|Abscess of salivary gland
C0155957|T047|AB|527.3|ICD9CM|Salivary gland abscess|Salivary gland abscess
C0036094|T190|PT|527.4|ICD9CM|Fistula of salivary gland|Fistula of salivary gland
C0036094|T190|AB|527.4|ICD9CM|Salivary gland fistula|Salivary gland fistula
C0036091|T047|AB|527.5|ICD9CM|Sialolithiasis|Sialolithiasis
C0036091|T047|PT|527.5|ICD9CM|Sialolithiasis|Sialolithiasis
C0026686|T047|PT|527.6|ICD9CM|Mucocele of salivary gland|Mucocele of salivary gland
C0026686|T047|AB|527.6|ICD9CM|Salivary gland mucocele|Salivary gland mucocele
C0012765|T046|PT|527.7|ICD9CM|Disturbance of salivary secretion|Disturbance of salivary secretion
C0012765|T046|AB|527.7|ICD9CM|Salivary secretion dis|Salivary secretion dis
C0029773|T047|PT|527.8|ICD9CM|Other specified diseases of the salivary glands|Other specified diseases of the salivary glands
C0029773|T047|AB|527.8|ICD9CM|Salivary gland dis NEC|Salivary gland dis NEC
C0036093|T047|AB|527.9|ICD9CM|Salivary gland dis NOS|Salivary gland dis NOS
C0036093|T047|PT|527.9|ICD9CM|Unspecified disease of the salivary glands|Unspecified disease of the salivary glands
C0155958|T047|HT|528|ICD9CM|Diseases of the oral soft tissues, excluding lesions specific for gingiva and tongue|Diseases of the oral soft tissues, excluding lesions specific for gingiva and tongue
C1719528|T047|HT|528.0|ICD9CM|Stomatitis and mucositis (ulcerative)|Stomatitis and mucositis (ulcerative)
C1719714|T047|PT|528.00|ICD9CM|Stomatitis and mucositis, unspecified|Stomatitis and mucositis, unspecified
C1719714|T047|AB|528.00|ICD9CM|Stomatitis/mucositis NOS|Stomatitis/mucositis NOS
C1719526|T047|PT|528.01|ICD9CM|Mucositis (ulcerative) due to antineoplastic therapy|Mucositis (ulcerative) due to antineoplastic therapy
C1719526|T047|AB|528.01|ICD9CM|Mucosits d/t antineo rx|Mucosits d/t antineo rx
C1719527|T047|PT|528.02|ICD9CM|Mucositis (ulcerative) due to other drugs|Mucositis (ulcerative) due to other drugs
C1719527|T047|AB|528.02|ICD9CM|Mucositis d/t drugs NEC|Mucositis d/t drugs NEC
C1719528|T047|PT|528.09|ICD9CM|Other stomatitis and mucositis (ulcerative)|Other stomatitis and mucositis (ulcerative)
C1719528|T047|AB|528.09|ICD9CM|Stomatits & mucosits NEC|Stomatits & mucosits NEC
C0028271|T047|AB|528.1|ICD9CM|Cancrum oris|Cancrum oris
C0028271|T047|PT|528.1|ICD9CM|Cancrum oris|Cancrum oris
C0038363|T047|AB|528.2|ICD9CM|Oral aphthae|Oral aphthae
C0038363|T047|PT|528.2|ICD9CM|Oral aphthae|Oral aphthae
C0007643|T047|PT|528.3|ICD9CM|Cellulitis and abscess of oral soft tissues|Cellulitis and abscess of oral soft tissues
C0007643|T047|AB|528.3|ICD9CM|Cellulitis/abscess mouth|Cellulitis/abscess mouth
C0155959|T047|PT|528.4|ICD9CM|Cysts of oral soft tissues|Cysts of oral soft tissues
C0155959|T047|AB|528.4|ICD9CM|Oral soft tissue cyst|Oral soft tissue cyst
C0023760|T047|AB|528.5|ICD9CM|Diseases of lips|Diseases of lips
C0023760|T047|PT|528.5|ICD9CM|Diseases of lips|Diseases of lips
C1112530|T047|PT|528.6|ICD9CM|Leukoplakia of oral mucosa, including tongue|Leukoplakia of oral mucosa, including tongue
C1112530|T047|AB|528.6|ICD9CM|Leukoplakia oral mucosa|Leukoplakia oral mucosa
C0155961|T047|HT|528.7|ICD9CM|Other disturbances of oral epithelium, including tongue|Other disturbances of oral epithelium, including tongue
C1456227|T047|AB|528.71|ICD9CM|Keratin ridge mucosa-min|Keratin ridge mucosa-min
C1456227|T047|PT|528.71|ICD9CM|Minimal keratinized residual ridge mucosa|Minimal keratinized residual ridge mucosa
C1456228|T047|PT|528.72|ICD9CM|Excessive keratinized residual ridge mucosa|Excessive keratinized residual ridge mucosa
C1456228|T047|AB|528.72|ICD9CM|Keratin ridge muc-excess|Keratin ridge muc-excess
C0155961|T047|AB|528.79|ICD9CM|Dist oral epithelium NEC|Dist oral epithelium NEC
C0155961|T047|PT|528.79|ICD9CM|Other disturbances of oral epithelium, including tongue|Other disturbances of oral epithelium, including tongue
C0029171|T047|AB|528.8|ICD9CM|Oral submucosal fibrosis|Oral submucosal fibrosis
C0029171|T047|PT|528.8|ICD9CM|Oral submucosal fibrosis, including of tongue|Oral submucosal fibrosis, including of tongue
C0029498|T047|AB|528.9|ICD9CM|Oral soft tissue dis NEC|Oral soft tissue dis NEC
C0029498|T047|PT|528.9|ICD9CM|Other and unspecified diseases of the oral soft tissues|Other and unspecified diseases of the oral soft tissues
C0155962|T047|HT|529|ICD9CM|Diseases and other conditions of the tongue|Diseases and other conditions of the tongue
C0017675|T047|AB|529.0|ICD9CM|Glossitis|Glossitis
C0017675|T047|PT|529.0|ICD9CM|Glossitis|Glossitis
C0017677|T047|AB|529.1|ICD9CM|Geographic tongue|Geographic tongue
C0017677|T047|PT|529.1|ICD9CM|Geographic tongue|Geographic tongue
C0155963|T019|AB|529.2|ICD9CM|Med rhomboid glossitis|Med rhomboid glossitis
C0155963|T019|PT|529.2|ICD9CM|Median rhomboid glossitis|Median rhomboid glossitis
C0392494|T047|AB|529.3|ICD9CM|Hypertroph tongue papill|Hypertroph tongue papill
C0392494|T047|PT|529.3|ICD9CM|Hypertrophy of tongue papillae|Hypertrophy of tongue papillae
C0155964|T047|PT|529.4|ICD9CM|Atrophy of tongue papillae|Atrophy of tongue papillae
C0155964|T047|AB|529.4|ICD9CM|Atrophy tongue papillae|Atrophy tongue papillae
C0040412|T047|AB|529.5|ICD9CM|Plicated tongue|Plicated tongue
C0040412|T047|PT|529.5|ICD9CM|Plicated tongue|Plicated tongue
C0017672|T184|AB|529.6|ICD9CM|Glossodynia|Glossodynia
C0017672|T184|PT|529.6|ICD9CM|Glossodynia|Glossodynia
C0155965|T047|PT|529.8|ICD9CM|Other specified conditions of the tongue|Other specified conditions of the tongue
C0155965|T047|AB|529.8|ICD9CM|Tongue disorder NEC|Tongue disorder NEC
C0040409|T047|AB|529.9|ICD9CM|Tongue disorder NOS|Tongue disorder NOS
C0040409|T047|PT|529.9|ICD9CM|Unspecified condition of the tongue|Unspecified condition of the tongue
C0014852|T047|HT|530|ICD9CM|Diseases of esophagus|Diseases of esophagus
C0178281|T047|HT|530-539.99|ICD9CM|DISEASES OF ESOPHAGUS, STOMACH, AND DUODENUM|DISEASES OF ESOPHAGUS, STOMACH, AND DUODENUM
C0014848|T047|AB|530.0|ICD9CM|Achalasia & cardiospasm|Achalasia & cardiospasm
C0014848|T047|PT|530.0|ICD9CM|Achalasia and cardiospasm|Achalasia and cardiospasm
C0014868|T047|HT|530.1|ICD9CM|Esophagitis|Esophagitis
C0014868|T047|AB|530.10|ICD9CM|Esophagitis, unspecified|Esophagitis, unspecified
C0014868|T047|PT|530.10|ICD9CM|Esophagitis, unspecified|Esophagitis, unspecified
C0014869|T047|AB|530.11|ICD9CM|Reflux esophagitis|Reflux esophagitis
C0014869|T047|PT|530.11|ICD9CM|Reflux esophagitis|Reflux esophagitis
C0149882|T047|AB|530.12|ICD9CM|Acute esophagitis|Acute esophagitis
C0149882|T047|PT|530.12|ICD9CM|Acute esophagitis|Acute esophagitis
C0341106|T047|PT|530.13|ICD9CM|Eosinophilic esophagitis|Eosinophilic esophagitis
C0341106|T047|AB|530.13|ICD9CM|Eosinophilic esophagitis|Eosinophilic esophagitis
C0375352|T047|AB|530.19|ICD9CM|Other esophagitis|Other esophagitis
C0375352|T047|PT|530.19|ICD9CM|Other esophagitis|Other esophagitis
C0151970|T047|HT|530.2|ICD9CM|Ulcer of esophagus|Ulcer of esophagus
C1260417|T047|AB|530.20|ICD9CM|Ulc esophagus w/o bleed|Ulc esophagus w/o bleed
C1260417|T047|PT|530.20|ICD9CM|Ulcer of esophagus without bleeding|Ulcer of esophagus without bleeding
C0236127|T047|AB|530.21|ICD9CM|Ulcer esophagus w bleed|Ulcer esophagus w bleed
C0236127|T047|PT|530.21|ICD9CM|Ulcer of esophagus with bleeding|Ulcer of esophagus with bleeding
C4551650|T047|AB|530.3|ICD9CM|Esophageal stricture|Esophageal stricture
C4551650|T047|PT|530.3|ICD9CM|Stricture and stenosis of esophagus|Stricture and stenosis of esophagus
C0014860|T046|AB|530.4|ICD9CM|Perforation of esophagus|Perforation of esophagus
C0014860|T046|PT|530.4|ICD9CM|Perforation of esophagus|Perforation of esophagus
C0014858|T047|AB|530.5|ICD9CM|Dyskinesia of esophagus|Dyskinesia of esophagus
C0014858|T047|PT|530.5|ICD9CM|Dyskinesia of esophagus|Dyskinesia of esophagus
C0155966|T020|AB|530.6|ICD9CM|Acq esophag diverticulum|Acq esophag diverticulum
C0155966|T020|PT|530.6|ICD9CM|Diverticulum of esophagus, acquired|Diverticulum of esophagus, acquired
C0024633|T047|PT|530.7|ICD9CM|Gastroesophageal laceration-hemorrhage syndrome|Gastroesophageal laceration-hemorrhage syndrome
C0024633|T047|AB|530.7|ICD9CM|Mallory-weiss syndrome|Mallory-weiss syndrome
C0348727|T047|HT|530.8|ICD9CM|Other specified disorders of esophagus|Other specified disorders of esophagus
C0017168|T047|AB|530.81|ICD9CM|Esophageal reflux|Esophageal reflux
C0017168|T047|PT|530.81|ICD9CM|Esophageal reflux|Esophageal reflux
C0239293|T046|AB|530.82|ICD9CM|Esophageal hemorrhage|Esophageal hemorrhage
C0239293|T046|PT|530.82|ICD9CM|Esophageal hemorrhage|Esophageal hemorrhage
C0267095|T191|AB|530.83|ICD9CM|Esophageal leukoplakia|Esophageal leukoplakia
C0267095|T191|PT|530.83|ICD9CM|Esophageal leukoplakia|Esophageal leukoplakia
C0040588|T190|PT|530.84|ICD9CM|Tracheoesophageal fistula|Tracheoesophageal fistula
C0040588|T190|AB|530.84|ICD9CM|Tracheoesophageal fstula|Tracheoesophageal fstula
C0004763|T047|AB|530.85|ICD9CM|Barrett's esophagus|Barrett's esophagus
C0004763|T047|PT|530.85|ICD9CM|Barrett's esophagus|Barrett's esophagus
C1456233|T046|AB|530.86|ICD9CM|Esophagostomy infection|Esophagostomy infection
C1456233|T046|PT|530.86|ICD9CM|Infection of esophagostomy|Infection of esophagostomy
C1456234|T046|AB|530.87|ICD9CM|Mech comp esophagostomy|Mech comp esophagostomy
C1456234|T046|PT|530.87|ICD9CM|Mechanical complication of esophagostomy|Mechanical complication of esophagostomy
C0348727|T047|AB|530.89|ICD9CM|Other dsrders esophagus|Other dsrders esophagus
C0348727|T047|PT|530.89|ICD9CM|Other specified disorders of esophagus|Other specified disorders of esophagus
C0014852|T047|AB|530.9|ICD9CM|Esophageal disorder NOS|Esophageal disorder NOS
C0014852|T047|PT|530.9|ICD9CM|Unspecified disorder of esophagus|Unspecified disorder of esophagus
C0038358|T047|HT|531|ICD9CM|Gastric ulcer|Gastric ulcer
C0155967|T047|HT|531.0|ICD9CM|Acute gastric ulcer with hemorrhage|Acute gastric ulcer with hemorrhage
C0155968|T047|AB|531.00|ICD9CM|Ac stomach ulcer w hem|Ac stomach ulcer w hem
C0155968|T047|PT|531.00|ICD9CM|Acute gastric ulcer with hemorrhage, without mention of obstruction|Acute gastric ulcer with hemorrhage, without mention of obstruction
C0155969|T047|AB|531.01|ICD9CM|Ac stomac ulc w hem-obst|Ac stomac ulc w hem-obst
C0155969|T047|PT|531.01|ICD9CM|Acute gastric ulcer with hemorrhage, with obstruction|Acute gastric ulcer with hemorrhage, with obstruction
C0155970|T047|HT|531.1|ICD9CM|Acute gastric ulcer with perforation|Acute gastric ulcer with perforation
C0155971|T047|AB|531.10|ICD9CM|Ac stomach ulcer w perf|Ac stomach ulcer w perf
C0155971|T047|PT|531.10|ICD9CM|Acute gastric ulcer with perforation, without mention of obstruction|Acute gastric ulcer with perforation, without mention of obstruction
C0155972|T047|AB|531.11|ICD9CM|Ac stom ulc w perf-obst|Ac stom ulc w perf-obst
C0155972|T047|PT|531.11|ICD9CM|Acute gastric ulcer with perforation, with obstruction|Acute gastric ulcer with perforation, with obstruction
C0155973|T047|HT|531.2|ICD9CM|Acute gastric ulcer with hemorrhage and perforation|Acute gastric ulcer with hemorrhage and perforation
C0267123|T047|AB|531.20|ICD9CM|Ac stomac ulc w hem/perf|Ac stomac ulc w hem/perf
C0267123|T047|PT|531.20|ICD9CM|Acute gastric ulcer with hemorrhage and perforation, without mention of obstruction|Acute gastric ulcer with hemorrhage and perforation, without mention of obstruction
C0155975|T047|AB|531.21|ICD9CM|Ac stom ulc hem/perf-obs|Ac stom ulc hem/perf-obs
C0155975|T047|PT|531.21|ICD9CM|Acute gastric ulcer with hemorrhage and perforation, with obstruction|Acute gastric ulcer with hemorrhage and perforation, with obstruction
C0267124|T047|HT|531.3|ICD9CM|Acute gastric ulcer without mention of hemorrhage or perforation|Acute gastric ulcer without mention of hemorrhage or perforation
C0267125|T047|PT|531.30|ICD9CM|Acute gastric ulcer without mention of hemorrhage or perforation, without mention of obstruction|Acute gastric ulcer without mention of hemorrhage or perforation, without mention of obstruction
C0267125|T047|AB|531.30|ICD9CM|Acute stomach ulcer NOS|Acute stomach ulcer NOS
C0155978|T047|AB|531.31|ICD9CM|Ac stomach ulc NOS-obstr|Ac stomach ulc NOS-obstr
C0155978|T047|PT|531.31|ICD9CM|Acute gastric ulcer without mention of hemorrhage or perforation, with obstruction|Acute gastric ulcer without mention of hemorrhage or perforation, with obstruction
C0155979|T047|HT|531.4|ICD9CM|Chronic or unspecified gastric ulcer with hemorrhage|Chronic or unspecified gastric ulcer with hemorrhage
C0155980|T047|AB|531.40|ICD9CM|Chr stomach ulc w hem|Chr stomach ulc w hem
C0155980|T047|PT|531.40|ICD9CM|Chronic or unspecified gastric ulcer with hemorrhage, without mention of obstruction|Chronic or unspecified gastric ulcer with hemorrhage, without mention of obstruction
C0155981|T047|AB|531.41|ICD9CM|Chr stom ulc w hem-obstr|Chr stom ulc w hem-obstr
C0155981|T047|PT|531.41|ICD9CM|Chronic or unspecified gastric ulcer with hemorrhage, with obstruction|Chronic or unspecified gastric ulcer with hemorrhage, with obstruction
C0155982|T047|HT|531.5|ICD9CM|Chronic or unspecified gastric ulcer with perforation|Chronic or unspecified gastric ulcer with perforation
C0155983|T047|AB|531.50|ICD9CM|Chr stomach ulcer w perf|Chr stomach ulcer w perf
C0155983|T047|PT|531.50|ICD9CM|Chronic or unspecified gastric ulcer with perforation, without mention of obstruction|Chronic or unspecified gastric ulcer with perforation, without mention of obstruction
C0155984|T047|AB|531.51|ICD9CM|Chr stom ulc w perf-obst|Chr stom ulc w perf-obst
C0155984|T047|PT|531.51|ICD9CM|Chronic or unspecified gastric ulcer with perforation, with obstruction|Chronic or unspecified gastric ulcer with perforation, with obstruction
C0494723|T047|HT|531.6|ICD9CM|Chronic or unspecified gastric ulcer with hemorrhage and perforation|Chronic or unspecified gastric ulcer with hemorrhage and perforation
C0155986|T047|AB|531.60|ICD9CM|Chr stomach ulc hem/perf|Chr stomach ulc hem/perf
C0155986|T047|PT|531.60|ICD9CM|Chronic or unspecified gastric ulcer with hemorrhage and perforation, without mention of obstruction|Chronic or unspecified gastric ulcer with hemorrhage and perforation, without mention of obstruction
C0155987|T047|AB|531.61|ICD9CM|Chr stom ulc hem/perf-ob|Chr stom ulc hem/perf-ob
C0155987|T047|PT|531.61|ICD9CM|Chronic or unspecified gastric ulcer with hemorrhage and perforation, with obstruction|Chronic or unspecified gastric ulcer with hemorrhage and perforation, with obstruction
C0267136|T047|HT|531.7|ICD9CM|Chronic gastric ulcer without mention of hemorrhage or perforation|Chronic gastric ulcer without mention of hemorrhage or perforation
C0155989|T047|AB|531.70|ICD9CM|Chr stomach ulcer NOS|Chr stomach ulcer NOS
C0155989|T047|PT|531.70|ICD9CM|Chronic gastric ulcer without mention of hemorrhage or perforation, without mention of obstruction|Chronic gastric ulcer without mention of hemorrhage or perforation, without mention of obstruction
C0267138|T047|AB|531.71|ICD9CM|Chr stomach ulc NOS-obst|Chr stomach ulc NOS-obst
C0267138|T047|PT|531.71|ICD9CM|Chronic gastric ulcer without mention of hemorrhage or perforation, with obstruction|Chronic gastric ulcer without mention of hemorrhage or perforation, with obstruction
C0400806|T047|HT|531.9|ICD9CM|Gastric ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation|Gastric ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation
C0400806|T047|AB|531.90|ICD9CM|Stomach ulcer NOS|Stomach ulcer NOS
C0155991|T047|AB|531.91|ICD9CM|Stomach ulcer NOS-obstr|Stomach ulcer NOS-obstr
C0013295|T047|HT|532|ICD9CM|Duodenal ulcer|Duodenal ulcer
C0155992|T047|HT|532.0|ICD9CM|Acute duodenal ulcer with hemorrhage|Acute duodenal ulcer with hemorrhage
C0155993|T047|AB|532.00|ICD9CM|Ac duodenal ulcer w hem|Ac duodenal ulcer w hem
C0155993|T047|PT|532.00|ICD9CM|Acute duodenal ulcer with hemorrhage, without mention of obstruction|Acute duodenal ulcer with hemorrhage, without mention of obstruction
C0155994|T047|AB|532.01|ICD9CM|Ac duoden ulc w hem-obst|Ac duoden ulc w hem-obst
C0155994|T047|PT|532.01|ICD9CM|Acute duodenal ulcer with hemorrhage, with obstruction|Acute duodenal ulcer with hemorrhage, with obstruction
C0155995|T047|HT|532.1|ICD9CM|Acute duodenal ulcer with perforation|Acute duodenal ulcer with perforation
C0267262|T047|AB|532.10|ICD9CM|Ac duodenal ulcer w perf|Ac duodenal ulcer w perf
C0267262|T047|PT|532.10|ICD9CM|Acute duodenal ulcer with perforation, without mention of obstruction|Acute duodenal ulcer with perforation, without mention of obstruction
C0155997|T047|AB|532.11|ICD9CM|Ac duoden ulc perf-obstr|Ac duoden ulc perf-obstr
C0155997|T047|PT|532.11|ICD9CM|Acute duodenal ulcer with perforation, with obstruction|Acute duodenal ulcer with perforation, with obstruction
C0155998|T047|HT|532.2|ICD9CM|Acute duodenal ulcer with hemorrhage and perforation|Acute duodenal ulcer with hemorrhage and perforation
C0155999|T047|AB|532.20|ICD9CM|Ac duoden ulc w hem/perf|Ac duoden ulc w hem/perf
C0155999|T047|PT|532.20|ICD9CM|Acute duodenal ulcer with hemorrhage and perforation, without mention of obstruction|Acute duodenal ulcer with hemorrhage and perforation, without mention of obstruction
C0156000|T047|AB|532.21|ICD9CM|Ac duod ulc hem/perf-obs|Ac duod ulc hem/perf-obs
C0156000|T047|PT|532.21|ICD9CM|Acute duodenal ulcer with hemorrhage and perforation, with obstruction|Acute duodenal ulcer with hemorrhage and perforation, with obstruction
C0156001|T047|HT|532.3|ICD9CM|Acute duodenal ulcer without mention of hemorrhage or perforation|Acute duodenal ulcer without mention of hemorrhage or perforation
C0156002|T047|AB|532.30|ICD9CM|Acute duodenal ulcer NOS|Acute duodenal ulcer NOS
C0156002|T047|PT|532.30|ICD9CM|Acute duodenal ulcer without mention of hemorrhage or perforation, without mention of obstruction|Acute duodenal ulcer without mention of hemorrhage or perforation, without mention of obstruction
C0156003|T047|AB|532.31|ICD9CM|Ac duodenal ulc NOS-obst|Ac duodenal ulc NOS-obst
C0156003|T047|PT|532.31|ICD9CM|Acute duodenal ulcer without mention of hemorrhage or perforation, with obstruction|Acute duodenal ulcer without mention of hemorrhage or perforation, with obstruction
C0156004|T047|HT|532.4|ICD9CM|Chronic or unspecified duodenal ulcer with hemorrhage|Chronic or unspecified duodenal ulcer with hemorrhage
C0156005|T047|AB|532.40|ICD9CM|Chr duoden ulcer w hem|Chr duoden ulcer w hem
C0156005|T047|PT|532.40|ICD9CM|Chronic or unspecified duodenal ulcer with hemorrhage, without mention of obstruction|Chronic or unspecified duodenal ulcer with hemorrhage, without mention of obstruction
C0156006|T047|AB|532.41|ICD9CM|Chr duoden ulc hem-obstr|Chr duoden ulc hem-obstr
C0156006|T047|PT|532.41|ICD9CM|Chronic or unspecified duodenal ulcer with hemorrhage, with obstruction|Chronic or unspecified duodenal ulcer with hemorrhage, with obstruction
C0391983|T047|HT|532.5|ICD9CM|Chronic or unspecified duodenal ulcer with perforation|Chronic or unspecified duodenal ulcer with perforation
C0156008|T047|AB|532.50|ICD9CM|Chr duoden ulcer w perf|Chr duoden ulcer w perf
C0156008|T047|PT|532.50|ICD9CM|Chronic or unspecified duodenal ulcer with perforation, without mention of obstruction|Chronic or unspecified duodenal ulcer with perforation, without mention of obstruction
C0156009|T047|AB|532.51|ICD9CM|Chr duoden ulc perf-obst|Chr duoden ulc perf-obst
C0156009|T047|PT|532.51|ICD9CM|Chronic or unspecified duodenal ulcer with perforation, with obstruction|Chronic or unspecified duodenal ulcer with perforation, with obstruction
C0494726|T047|HT|532.6|ICD9CM|Chronic or unspecified duodenal ulcer with hemorrhage and perforation|Chronic or unspecified duodenal ulcer with hemorrhage and perforation
C0156011|T047|AB|532.60|ICD9CM|Chr duoden ulc hem/perf|Chr duoden ulc hem/perf
C0156012|T047|AB|532.61|ICD9CM|Chr duod ulc hem/perf-ob|Chr duod ulc hem/perf-ob
C0156012|T047|PT|532.61|ICD9CM|Chronic or unspecified duodenal ulcer with hemorrhage and perforation, with obstruction|Chronic or unspecified duodenal ulcer with hemorrhage and perforation, with obstruction
C0267282|T047|HT|532.7|ICD9CM|Chronic duodenal ulcer without mention of hemorrhage or perforation|Chronic duodenal ulcer without mention of hemorrhage or perforation
C0156014|T047|AB|532.70|ICD9CM|Chr duodenal ulcer NOS|Chr duodenal ulcer NOS
C0156014|T047|PT|532.70|ICD9CM|Chronic duodenal ulcer without mention of hemorrhage or perforation, without mention of obstruction|Chronic duodenal ulcer without mention of hemorrhage or perforation, without mention of obstruction
C0156015|T047|AB|532.71|ICD9CM|Chr duoden ulc NOS-obstr|Chr duoden ulc NOS-obstr
C0156015|T047|PT|532.71|ICD9CM|Chronic duodenal ulcer without mention of hemorrhage or perforation, with obstruction|Chronic duodenal ulcer without mention of hemorrhage or perforation, with obstruction
C0391984|T047|HT|532.9|ICD9CM|Duodenal ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation|Duodenal ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation
C0489962|T047|AB|532.90|ICD9CM|Duodenal ulcer NOS|Duodenal ulcer NOS
C0156016|T047|AB|532.91|ICD9CM|Duodenal ulcer NOS-obstr|Duodenal ulcer NOS-obstr
C0030920|T047|HT|533|ICD9CM|Peptic ulcer, site unspecified|Peptic ulcer, site unspecified
C0267288|T047|HT|533.0|ICD9CM|Acute peptic ulcer of unspecified site with hemorrhage|Acute peptic ulcer of unspecified site with hemorrhage
C0267288|T047|AB|533.00|ICD9CM|Ac peptic ulcer w hemorr|Ac peptic ulcer w hemorr
C0267288|T047|PT|533.00|ICD9CM|Acute peptic ulcer of unspecified site with hemorrhage, without mention of obstruction|Acute peptic ulcer of unspecified site with hemorrhage, without mention of obstruction
C0156019|T047|AB|533.01|ICD9CM|Ac peptic ulc w hem-obst|Ac peptic ulc w hem-obst
C0156019|T047|PT|533.01|ICD9CM|Acute peptic ulcer of unspecified site with hemorrhage, with obstruction|Acute peptic ulcer of unspecified site with hemorrhage, with obstruction
C0267291|T047|HT|533.1|ICD9CM|Acute peptic ulcer of unspecified site with perforation|Acute peptic ulcer of unspecified site with perforation
C1442967|T047|AB|533.10|ICD9CM|Ac peptic ulcer w perfor|Ac peptic ulcer w perfor
C1442967|T047|PT|533.10|ICD9CM|Acute peptic ulcer of unspecified site with perforation, without mention of obstruction|Acute peptic ulcer of unspecified site with perforation, without mention of obstruction
C0156022|T047|AB|533.11|ICD9CM|Ac peptic ulc w perf-obs|Ac peptic ulc w perf-obs
C0156022|T047|PT|533.11|ICD9CM|Acute peptic ulcer of unspecified site with perforation, with obstruction|Acute peptic ulcer of unspecified site with perforation, with obstruction
C0267294|T047|HT|533.2|ICD9CM|Acute peptic ulcer of unspecified site with hemorrhage and perforation|Acute peptic ulcer of unspecified site with hemorrhage and perforation
C0156024|T047|AB|533.20|ICD9CM|Ac peptic ulc w hem/perf|Ac peptic ulc w hem/perf
C0156025|T047|AB|533.21|ICD9CM|Ac pept ulc hem/perf-obs|Ac pept ulc hem/perf-obs
C0156025|T047|PT|533.21|ICD9CM|Acute peptic ulcer of unspecified site with hemorrhage and perforation, with obstruction|Acute peptic ulcer of unspecified site with hemorrhage and perforation, with obstruction
C0392499|T047|HT|533.3|ICD9CM|Acute peptic ulcer of unspecified site without mention of hemorrhage and perforation|Acute peptic ulcer of unspecified site without mention of hemorrhage and perforation
C0267298|T047|AB|533.30|ICD9CM|Acute peptic ulcer NOS|Acute peptic ulcer NOS
C0156024|T047|AB|533.31|ICD9CM|Ac peptic ulcer NOS-obst|Ac peptic ulcer NOS-obst
C0494730|T047|HT|533.4|ICD9CM|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage
C0156029|T047|AB|533.40|ICD9CM|Chr peptic ulcer w hem|Chr peptic ulcer w hem
C0156030|T047|AB|533.41|ICD9CM|Chr peptic ulc w hem-obs|Chr peptic ulc w hem-obs
C0156030|T047|PT|533.41|ICD9CM|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage, with obstruction|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage, with obstruction
C0494731|T047|HT|533.5|ICD9CM|Chronic or unspecified peptic ulcer of unspecified site with perforation|Chronic or unspecified peptic ulcer of unspecified site with perforation
C0156032|T047|AB|533.50|ICD9CM|Chr peptic ulcer w perf|Chr peptic ulcer w perf
C0156033|T047|AB|533.51|ICD9CM|Chr peptic ulc perf-obst|Chr peptic ulc perf-obst
C0156033|T047|PT|533.51|ICD9CM|Chronic or unspecified peptic ulcer of unspecified site with perforation, with obstruction|Chronic or unspecified peptic ulcer of unspecified site with perforation, with obstruction
C0494732|T047|HT|533.6|ICD9CM|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage and perforation|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage and perforation
C0156035|T047|AB|533.60|ICD9CM|Chr pept ulc w hem/perf|Chr pept ulc w hem/perf
C0156036|T047|AB|533.61|ICD9CM|Chr pept ulc hem/perf-ob|Chr pept ulc hem/perf-ob
C1279396|T047|HT|533.7|ICD9CM|Chronic peptic ulcer of unspecified site without mention of hemorrhage or perforation|Chronic peptic ulcer of unspecified site without mention of hemorrhage or perforation
C1961834|T047|AB|533.70|ICD9CM|Chronic peptic ulcer NOS|Chronic peptic ulcer NOS
C0156039|T047|AB|533.71|ICD9CM|Chr peptic ulcer NOS-obs|Chr peptic ulcer NOS-obs
C0030924|T020|AB|533.90|ICD9CM|Peptic ulcer NOS|Peptic ulcer NOS
C0156040|T047|AB|533.91|ICD9CM|Peptic ulcer NOS-obstruc|Peptic ulcer NOS-obstruc
C1384631|T020|HT|534|ICD9CM|Gastrojejunal ulcer|Gastrojejunal ulcer
C0156042|T047|HT|534.0|ICD9CM|Acute gastrojejunal ulcer with hemorrhage|Acute gastrojejunal ulcer with hemorrhage
C0156043|T047|AB|534.00|ICD9CM|Ac marginal ulcer w hem|Ac marginal ulcer w hem
C0156043|T047|PT|534.00|ICD9CM|Acute gastrojejunal ulcer with hemorrhage, without mention of obstruction|Acute gastrojejunal ulcer with hemorrhage, without mention of obstruction
C0156044|T047|AB|534.01|ICD9CM|Ac margin ulc w hem-obst|Ac margin ulc w hem-obst
C0156044|T047|PT|534.01|ICD9CM|Acute gastrojejunal ulcer, with hemorrhage, with obstruction|Acute gastrojejunal ulcer, with hemorrhage, with obstruction
C0156045|T047|HT|534.1|ICD9CM|Acute gastrojejunal ulcer with perforation|Acute gastrojejunal ulcer with perforation
C0156046|T047|AB|534.10|ICD9CM|Ac marginal ulcer w perf|Ac marginal ulcer w perf
C0156046|T047|PT|534.10|ICD9CM|Acute gastrojejunal ulcer with perforation, without mention of obstruction|Acute gastrojejunal ulcer with perforation, without mention of obstruction
C0156047|T047|AB|534.11|ICD9CM|Ac margin ulc w perf-obs|Ac margin ulc w perf-obs
C0156047|T047|PT|534.11|ICD9CM|Acute gastrojejunal ulcer with perforation, with obstruction|Acute gastrojejunal ulcer with perforation, with obstruction
C0156048|T047|HT|534.2|ICD9CM|Acute gastrojejunal ulcer with hemorrhage and perforation|Acute gastrojejunal ulcer with hemorrhage and perforation
C0156049|T047|AB|534.20|ICD9CM|Ac margin ulc w hem/perf|Ac margin ulc w hem/perf
C0156049|T047|PT|534.20|ICD9CM|Acute gastrojejunal ulcer with hemorrhage and perforation, without mention of obstruction|Acute gastrojejunal ulcer with hemorrhage and perforation, without mention of obstruction
C0156050|T047|AB|534.21|ICD9CM|Ac marg ulc hem/perf-obs|Ac marg ulc hem/perf-obs
C0156050|T047|PT|534.21|ICD9CM|Acute gastrojejunal ulcer with hemorrhage and perforation, with obstruction|Acute gastrojejunal ulcer with hemorrhage and perforation, with obstruction
C0392501|T020|HT|534.3|ICD9CM|Acute gastrojejunal ulcer without mention of hemorrhage or perforation|Acute gastrojejunal ulcer without mention of hemorrhage or perforation
C0267326|T020|AB|534.30|ICD9CM|Ac marginal ulcer NOS|Ac marginal ulcer NOS
C0156053|T047|AB|534.31|ICD9CM|Ac marginal ulc NOS-obst|Ac marginal ulc NOS-obst
C0156053|T047|PT|534.31|ICD9CM|Acute gastrojejunal ulcer without mention of hemorrhage or perforation, with obstruction|Acute gastrojejunal ulcer without mention of hemorrhage or perforation, with obstruction
C0156054|T047|HT|534.4|ICD9CM|Chronic or unspecified gastrojejunal ulcer with hemorrhage|Chronic or unspecified gastrojejunal ulcer with hemorrhage
C0156055|T047|AB|534.40|ICD9CM|Chr marginal ulcer w hem|Chr marginal ulcer w hem
C0156055|T047|PT|534.40|ICD9CM|Chronic or unspecified gastrojejunal ulcer with hemorrhage, without mention of obstruction|Chronic or unspecified gastrojejunal ulcer with hemorrhage, without mention of obstruction
C0156056|T047|AB|534.41|ICD9CM|Chr margin ulc w hem-obs|Chr margin ulc w hem-obs
C0156056|T047|PT|534.41|ICD9CM|Chronic or unspecified gastrojejunal ulcer, with hemorrhage, with obstruction|Chronic or unspecified gastrojejunal ulcer, with hemorrhage, with obstruction
C0156057|T047|HT|534.5|ICD9CM|Chronic or unspecified gastrojejunal ulcer with perforation|Chronic or unspecified gastrojejunal ulcer with perforation
C0156058|T047|AB|534.50|ICD9CM|Chr marginal ulc w perf|Chr marginal ulc w perf
C0156058|T047|PT|534.50|ICD9CM|Chronic or unspecified gastrojejunal ulcer with perforation, without mention of obstruction|Chronic or unspecified gastrojejunal ulcer with perforation, without mention of obstruction
C0156059|T047|AB|534.51|ICD9CM|Chr margin ulc perf-obst|Chr margin ulc perf-obst
C0156059|T047|PT|534.51|ICD9CM|Chronic or unspecified gastrojejunal ulcer with perforation, with obstruction|Chronic or unspecified gastrojejunal ulcer with perforation, with obstruction
C0494735|T047|HT|534.6|ICD9CM|Chronic or unspecified gastrojejunal ulcer with hemorrhage and perforation|Chronic or unspecified gastrojejunal ulcer with hemorrhage and perforation
C0156061|T047|AB|534.60|ICD9CM|Chr margin ulc hem/perf|Chr margin ulc hem/perf
C0156062|T047|AB|534.61|ICD9CM|Chr marg ulc hem/perf-ob|Chr marg ulc hem/perf-ob
C0156062|T047|PT|534.61|ICD9CM|Chronic or unspecified gastrojejunal ulcer with hemorrhage and perforation, with obstruction|Chronic or unspecified gastrojejunal ulcer with hemorrhage and perforation, with obstruction
C0392502|T020|HT|534.7|ICD9CM|Chronic gastrojejunal ulcer without mention of hemorrhage or perforation|Chronic gastrojejunal ulcer without mention of hemorrhage or perforation
C0267347|T020|AB|534.70|ICD9CM|Chr marginal ulcer NOS|Chr marginal ulcer NOS
C0156065|T047|AB|534.71|ICD9CM|Chr marginal ulc NOS-obs|Chr marginal ulc NOS-obs
C0156065|T047|PT|534.71|ICD9CM|Chronic gastrojejunal ulcer without mention of hemorrhage or perforation, with obstruction|Chronic gastrojejunal ulcer without mention of hemorrhage or perforation, with obstruction
C0494736|T047|HT|534.9|ICD9CM|Gastrojejunal ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation|Gastrojejunal ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation
C0156067|T047|AB|534.90|ICD9CM|Gastrojejunal ulcer NOS|Gastrojejunal ulcer NOS
C0156068|T047|AB|534.91|ICD9CM|Gastrojejun ulc NOS-obst|Gastrojejun ulc NOS-obst
C0267166|T047|HT|535|ICD9CM|Gastritis and duodenitis|Gastritis and duodenitis
C0149518|T047|HT|535.0|ICD9CM|Acute gastritis|Acute gastritis
C0156070|T047|PT|535.00|ICD9CM|Acute gastritis, without mention of hemorrhage|Acute gastritis, without mention of hemorrhage
C0156070|T047|AB|535.00|ICD9CM|Acute gastrtis w/o hmrhg|Acute gastrtis w/o hmrhg
C2243087|T047|AB|535.01|ICD9CM|Acute gastritis w hmrhg|Acute gastritis w hmrhg
C2243087|T047|PT|535.01|ICD9CM|Acute gastritis, with hemorrhage|Acute gastritis, with hemorrhage
C0017154|T047|HT|535.1|ICD9CM|Atrophic gastritis|Atrophic gastritis
C0156072|T047|PT|535.10|ICD9CM|Atrophic gastritis, without mention of hemorrhage|Atrophic gastritis, without mention of hemorrhage
C0156072|T047|AB|535.10|ICD9CM|Atrph gastrtis w/o hmrhg|Atrph gastrtis w/o hmrhg
C0156073|T047|PT|535.11|ICD9CM|Atrophic gastritis, with hemorrhage|Atrophic gastritis, with hemorrhage
C0156073|T047|AB|535.11|ICD9CM|Atrph gastritis w hmrhg|Atrph gastritis w hmrhg
C0017155|T047|HT|535.2|ICD9CM|Gastric mucosal hypertrophy|Gastric mucosal hypertrophy
C0156074|T047|PT|535.20|ICD9CM|Gastric mucosal hypertrophy, without mention of hemorrhage|Gastric mucosal hypertrophy, without mention of hemorrhage
C0156074|T047|AB|535.20|ICD9CM|Gstr mcsl hyprt w/o hmrg|Gstr mcsl hyprt w/o hmrg
C0156075|T047|PT|535.21|ICD9CM|Gastric mucosal hypertrophy, with hemorrhage|Gastric mucosal hypertrophy, with hemorrhage
C0156075|T047|AB|535.21|ICD9CM|Gstr mcsl hyprt w hmrg|Gstr mcsl hyprt w hmrg
C0156076|T047|HT|535.3|ICD9CM|Alcoholic gastritis|Alcoholic gastritis
C0156077|T047|AB|535.30|ICD9CM|Alchl gastrtis w/o hmrhg|Alchl gastrtis w/o hmrhg
C0156077|T047|PT|535.30|ICD9CM|Alcoholic gastritis, without mention of hemorrhage|Alcoholic gastritis, without mention of hemorrhage
C0156078|T047|AB|535.31|ICD9CM|Alchl gstritis w hmrhg|Alchl gstritis w hmrhg
C0156078|T047|PT|535.31|ICD9CM|Alcoholic gastritis, with hemorrhage|Alcoholic gastritis, with hemorrhage
C0029800|T047|HT|535.4|ICD9CM|Other specified gastritis|Other specified gastritis
C0156079|T047|AB|535.40|ICD9CM|Oth spf gstrt w/o hmrhg|Oth spf gstrt w/o hmrhg
C0156079|T047|PT|535.40|ICD9CM|Other specified gastritis, without mention of hemorrhage|Other specified gastritis, without mention of hemorrhage
C0156080|T047|AB|535.41|ICD9CM|Oth spf gastrt w hmrhg|Oth spf gastrt w hmrhg
C0156080|T047|PT|535.41|ICD9CM|Other specified gastritis, with hemorrhage|Other specified gastritis, with hemorrhage
C0041841|T047|HT|535.5|ICD9CM|Unspecified gastritis and gastroduodenitis|Unspecified gastritis and gastroduodenitis
C0156081|T047|AB|535.50|ICD9CM|Gstr/ddnts NOS w/o hmrhg|Gstr/ddnts NOS w/o hmrhg
C0156081|T047|PT|535.50|ICD9CM|Unspecified gastritis and gastroduodenitis, without mention of hemorrhage|Unspecified gastritis and gastroduodenitis, without mention of hemorrhage
C0156082|T047|AB|535.51|ICD9CM|Gstr/ddnts NOS w hmrhg|Gstr/ddnts NOS w hmrhg
C0156082|T047|PT|535.51|ICD9CM|Unspecified gastritis and gastroduodenitis, with hemorrhage|Unspecified gastritis and gastroduodenitis, with hemorrhage
C0013298|T047|HT|535.6|ICD9CM|Duodenitis|Duodenitis
C0156083|T047|AB|535.60|ICD9CM|Duodenitis w/o hmrhg|Duodenitis w/o hmrhg
C0156083|T047|PT|535.60|ICD9CM|Duodenitis, without mention of hemorrhage|Duodenitis, without mention of hemorrhage
C0341245|T047|AB|535.61|ICD9CM|Duodenitis w hmrhg|Duodenitis w hmrhg
C0341245|T047|PT|535.61|ICD9CM|Duodenitis, with hemorrhage|Duodenitis, with hemorrhage
C0267154|T047|HT|535.7|ICD9CM|Eosinophilic gastritis|Eosinophilic gastritis
C2349565|T047|AB|535.70|ICD9CM|Eosinophil gastrt wo hem|Eosinophil gastrt wo hem
C2349565|T047|PT|535.70|ICD9CM|Eosinophilic gastritis, without mention of hemorrhage|Eosinophilic gastritis, without mention of hemorrhage
C2349566|T047|AB|535.71|ICD9CM|Eosinophilc gastrt w hem|Eosinophilc gastrt w hem
C2349566|T047|PT|535.71|ICD9CM|Eosinophilic gastritis, with hemorrhage|Eosinophilic gastritis, with hemorrhage
C0156084|T047|HT|536|ICD9CM|Disorders of function of stomach|Disorders of function of stomach
C0001075|T046|AB|536.0|ICD9CM|Achlorhydria|Achlorhydria
C0001075|T046|PT|536.0|ICD9CM|Achlorhydria|Achlorhydria
C0149823|T033|AB|536.1|ICD9CM|Ac dilation of stomach|Ac dilation of stomach
C0149823|T033|PT|536.1|ICD9CM|Acute dilatation of stomach|Acute dilatation of stomach
C0152165|T184|AB|536.2|ICD9CM|Persistent vomiting|Persistent vomiting
C0152165|T184|PT|536.2|ICD9CM|Persistent vomiting|Persistent vomiting
C0152020|T047|AB|536.3|ICD9CM|Gastroparesis|Gastroparesis
C0152020|T047|PT|536.3|ICD9CM|Gastroparesis|Gastroparesis
C0587245|T046|HT|536.4|ICD9CM|Gastrostomy complications|Gastrostomy complications
C0587245|T046|AB|536.40|ICD9CM|Gastrostomy comp NOS|Gastrostomy comp NOS
C0587245|T046|PT|536.40|ICD9CM|Gastrostomy complication, unspecified|Gastrostomy complication, unspecified
C0695239|T047|AB|536.41|ICD9CM|Gastrostomy infection|Gastrostomy infection
C0695239|T047|PT|536.41|ICD9CM|Infection of gastrostomy|Infection of gastrostomy
C0695240|T046|AB|536.42|ICD9CM|Gastrostomy comp - mech|Gastrostomy comp - mech
C0695240|T046|PT|536.42|ICD9CM|Mechanical complication of gastrostomy|Mechanical complication of gastrostomy
C0695241|T046|AB|536.49|ICD9CM|Gastrostomy comp NEC|Gastrostomy comp NEC
C0695241|T046|PT|536.49|ICD9CM|Other gastrostomy complications|Other gastrostomy complications
C0013396|T047|PT|536.8|ICD9CM|Dyspepsia and other specified disorders of function of stomach|Dyspepsia and other specified disorders of function of stomach
C0013396|T047|AB|536.8|ICD9CM|Stomach function dis NEC|Stomach function dis NEC
C0156084|T047|AB|536.9|ICD9CM|Stomach function dis NOS|Stomach function dis NOS
C0156084|T047|PT|536.9|ICD9CM|Unspecified functional disorder of stomach|Unspecified functional disorder of stomach
C0156086|T047|HT|537|ICD9CM|Other disorders of stomach and duodenum|Other disorders of stomach and duodenum
C0700588|T020|AB|537.0|ICD9CM|Acq pyloric stenosis|Acq pyloric stenosis
C0700588|T020|PT|537.0|ICD9CM|Acquired hypertrophic pyloric stenosis|Acquired hypertrophic pyloric stenosis
C0038355|T190|AB|537.1|ICD9CM|Gastric diverticulum|Gastric diverticulum
C0038355|T190|PT|537.1|ICD9CM|Gastric diverticulum|Gastric diverticulum
C0156087|T047|AB|537.2|ICD9CM|Chronic duodenal ileus|Chronic duodenal ileus
C0156087|T047|PT|537.2|ICD9CM|Chronic duodenal ileus|Chronic duodenal ileus
C0029679|T047|AB|537.3|ICD9CM|Duodenal obstruction NEC|Duodenal obstruction NEC
C0029679|T047|PT|537.3|ICD9CM|Other obstruction of duodenum|Other obstruction of duodenum
C0267180|T190|PT|537.4|ICD9CM|Fistula of stomach or duodenum|Fistula of stomach or duodenum
C0267180|T190|AB|537.4|ICD9CM|Gastric/duodenal fistula|Gastric/duodenal fistula
C0156088|T190|AB|537.5|ICD9CM|Gastroptosis|Gastroptosis
C0156088|T190|PT|537.5|ICD9CM|Gastroptosis|Gastroptosis
C0267183|T047|PT|537.6|ICD9CM|Hourglass stricture or stenosis of stomach|Hourglass stricture or stenosis of stomach
C0267183|T047|AB|537.6|ICD9CM|Hourglass stricture stom|Hourglass stricture stom
C0348731|T047|HT|537.8|ICD9CM|Other specified disorders of stomach and duodenum|Other specified disorders of stomach and duodenum
C0152163|T047|AB|537.81|ICD9CM|Pylorospasm|Pylorospasm
C0152163|T047|PT|537.81|ICD9CM|Pylorospasm|Pylorospasm
C0156090|T047|AB|537.82|ICD9CM|Angio stm/dudn w/o hmrhg|Angio stm/dudn w/o hmrhg
C0156090|T047|PT|537.82|ICD9CM|Angiodysplasia of stomach and duodenum without mention of hemorrhage|Angiodysplasia of stomach and duodenum without mention of hemorrhage
C0156091|T047|AB|537.83|ICD9CM|Angio stm/dudn w hmrhg|Angio stm/dudn w hmrhg
C0156091|T047|PT|537.83|ICD9CM|Angiodysplasia of stomach and duodenum with hemorrhage|Angiodysplasia of stomach and duodenum with hemorrhage
C1135229|T047|AB|537.84|ICD9CM|Dieulafoy les,stom&duod|Dieulafoy les,stom&duod
C1135229|T047|PT|537.84|ICD9CM|Dieulafoy lesion (hemorrhagic) of stomach and duodenum|Dieulafoy lesion (hemorrhagic) of stomach and duodenum
C0348731|T047|AB|537.89|ICD9CM|Gastroduodenal dis NEC|Gastroduodenal dis NEC
C0348731|T047|PT|537.89|ICD9CM|Other specified disorders of stomach and duodenum|Other specified disorders of stomach and duodenum
C0494741|T047|AB|537.9|ICD9CM|Gastroduodenal dis NOS|Gastroduodenal dis NOS
C0494741|T047|PT|537.9|ICD9CM|Unspecified disorder of stomach and duodenum|Unspecified disorder of stomach and duodenum
C3874327|T047|PT|538|ICD9CM|Gastrointestinal mucositis (ulcerative)|Gastrointestinal mucositis (ulcerative)
C3874327|T047|AB|538|ICD9CM|GI mucositis (ulceratve)|GI mucositis (ulceratve)
C3161254|T046|HT|539|ICD9CM|Complications of bariatric procedures|Complications of bariatric procedures
C3161255|T046|HT|539.0|ICD9CM|Complications of gastric band procedure|Complications of gastric band procedure
C3161113|T046|AB|539.01|ICD9CM|Inf d/t gastrc band proc|Inf d/t gastrc band proc
C3161113|T046|PT|539.01|ICD9CM|Infection due to gastric band procedure|Infection due to gastric band procedure
C3161114|T046|AB|539.09|ICD9CM|Oth cmp gastrc band proc|Oth cmp gastrc band proc
C3161114|T046|PT|539.09|ICD9CM|Other complications of gastric band procedure|Other complications of gastric band procedure
C3161256|T046|HT|539.8|ICD9CM|Complications of other bariatric procedure|Complications of other bariatric procedure
C3161115|T046|AB|539.81|ICD9CM|Inf d/t ot bariatrc proc|Inf d/t ot bariatrc proc
C3161115|T046|PT|539.81|ICD9CM|Infection due to other bariatric procedure|Infection due to other bariatric procedure
C3161116|T046|AB|539.89|ICD9CM|Ot comp ot bariatrc proc|Ot comp ot bariatrc proc
C3161116|T046|PT|539.89|ICD9CM|Other complications of other bariatric procedure|Other complications of other bariatric procedure
C0085693|T047|HT|540|ICD9CM|Acute appendicitis|Acute appendicitis
C0003615|T047|HT|540-543.99|ICD9CM|APPENDICITIS|APPENDICITIS
C0156092|T047|AB|540.0|ICD9CM|Ac append w peritonitis|Ac append w peritonitis
C0156092|T047|PT|540.0|ICD9CM|Acute appendicitis with generalized peritonitis|Acute appendicitis with generalized peritonitis
C0156093|T047|AB|540.1|ICD9CM|Abscess of appendix|Abscess of appendix
C0156093|T047|PT|540.1|ICD9CM|Acute appendicitis with peritoneal abscess|Acute appendicitis with peritoneal abscess
C0156094|T047|AB|540.9|ICD9CM|Acute appendicitis NOS|Acute appendicitis NOS
C0156094|T047|PT|540.9|ICD9CM|Acute appendicitis without mention of peritonitis|Acute appendicitis without mention of peritonitis
C0003615|T047|AB|541|ICD9CM|Appendicitis NOS|Appendicitis NOS
C0003615|T047|PT|541|ICD9CM|Appendicitis, unqualified|Appendicitis, unqualified
C0156095|T047|AB|542|ICD9CM|Other appendicitis|Other appendicitis
C0156095|T047|PT|542|ICD9CM|Other appendicitis|Other appendicitis
C0156098|T047|HT|543|ICD9CM|Other diseases of appendix|Other diseases of appendix
C1384587|T046|AB|543.0|ICD9CM|Hyperplasia of appendix|Hyperplasia of appendix
C1384587|T046|PT|543.0|ICD9CM|Hyperplasia of appendix (lymphoid)|Hyperplasia of appendix (lymphoid)
C0156098|T047|AB|543.9|ICD9CM|Diseases of appendix NEC|Diseases of appendix NEC
C0156098|T047|PT|543.9|ICD9CM|Other and unspecified diseases of appendix|Other and unspecified diseases of appendix
C0019294|T190|HT|550|ICD9CM|Inguinal hernia|Inguinal hernia
C0178282|T190|HT|550-553.99|ICD9CM|HERNIA OF ABDOMINAL CAVITY|HERNIA OF ABDOMINAL CAVITY
C0156099|T047|HT|550.0|ICD9CM|Inguinal hernia, with gangrene|Inguinal hernia, with gangrene
C0156100|T020|PT|550.00|ICD9CM|Inguinal hernia, with gangrene, unilateral or unspecified (not specified as recurrent)|Inguinal hernia, with gangrene, unilateral or unspecified (not specified as recurrent)
C0156100|T020|AB|550.00|ICD9CM|Unilat ing hernia w gang|Unilat ing hernia w gang
C0156101|T020|PT|550.01|ICD9CM|Inguinal hernia, with gangrene, unilateral or unspecified, recurrent|Inguinal hernia, with gangrene, unilateral or unspecified, recurrent
C0156101|T020|AB|550.01|ICD9CM|Recur unil ing hern-gang|Recur unil ing hern-gang
C0375354|T020|AB|550.02|ICD9CM|Bilat ing hernia w gang|Bilat ing hernia w gang
C0375354|T020|PT|550.02|ICD9CM|Inguinal hernia, with gangrene, bilateral (not specified as recurrent)|Inguinal hernia, with gangrene, bilateral (not specified as recurrent)
C0156103|T047|PT|550.03|ICD9CM|Inguinal hernia, with gangrene, bilateral, recurrent|Inguinal hernia, with gangrene, bilateral, recurrent
C0156103|T047|AB|550.03|ICD9CM|Recur bil ing hern-gang|Recur bil ing hern-gang
C0156104|T020|HT|550.1|ICD9CM|Inguinal hernia, with obstruction, without mention of gangrene|Inguinal hernia, with obstruction, without mention of gangrene
C0554123|T020|AB|550.10|ICD9CM|Unilat ing hernia w obst|Unilat ing hernia w obst
C0156106|T020|PT|550.11|ICD9CM|Inguinal hernia, with obstruction, without mention of gangrene, unilateral or unspecified,recurrent|Inguinal hernia, with obstruction, without mention of gangrene, unilateral or unspecified,recurrent
C0156106|T020|AB|550.11|ICD9CM|Recur unil ing hern-obst|Recur unil ing hern-obst
C0401080|T020|AB|550.12|ICD9CM|Bilat ing hernia w obst|Bilat ing hernia w obst
C0554121|T020|PT|550.13|ICD9CM|Inguinal hernia, with obstruction, without mention of gangrene, bilateral, recurrent|Inguinal hernia, with obstruction, without mention of gangrene, bilateral, recurrent
C0554121|T020|AB|550.13|ICD9CM|Recur bil ing hern-obstr|Recur bil ing hern-obstr
C0021447|T190|HT|550.9|ICD9CM|Inguinal hernia, without mention of obstruction or gangrene|Inguinal hernia, without mention of obstruction or gangrene
C0156109|T020|AB|550.90|ICD9CM|Unilat inguinal hernia|Unilat inguinal hernia
C0156110|T020|PT|550.91|ICD9CM|Inguinal hernia, without mention of obstruction or gangrene, unilateral or unspecified, recurrent|Inguinal hernia, without mention of obstruction or gangrene, unilateral or unspecified, recurrent
C0156110|T020|AB|550.91|ICD9CM|Recur unilat inguin hern|Recur unilat inguin hern
C0156111|T020|AB|550.92|ICD9CM|Bilat inguinal hernia|Bilat inguinal hernia
C0156111|T020|PT|550.92|ICD9CM|Inguinal hernia, without mention of obstruction or gangrene, bilateral (not specified as recurrent)|Inguinal hernia, without mention of obstruction or gangrene, bilateral (not specified as recurrent)
C0156112|T020|PT|550.93|ICD9CM|Inguinal hernia, without mention of obstruction or gangrene, bilateral, recurrent|Inguinal hernia, without mention of obstruction or gangrene, bilateral, recurrent
C0156112|T020|AB|550.93|ICD9CM|Recur bilat inguin hern|Recur bilat inguin hern
C0156113|T020|HT|551|ICD9CM|Other hernia of abdominal cavity, with gangrene|Other hernia of abdominal cavity, with gangrene
C0156114|T047|HT|551.0|ICD9CM|Femoral hernia with gangrene|Femoral hernia with gangrene
C0156115|T020|PT|551.00|ICD9CM|Femoral hernia with gangrene, unilateral or unspecified (not specified as recurrent)|Femoral hernia with gangrene, unilateral or unspecified (not specified as recurrent)
C0156115|T020|AB|551.00|ICD9CM|Unil femoral hern w gang|Unil femoral hern w gang
C0156116|T020|PT|551.01|ICD9CM|Femoral hernia with gangrene, unilateral or unspecified, recurrent|Femoral hernia with gangrene, unilateral or unspecified, recurrent
C0156116|T020|AB|551.01|ICD9CM|Rec unil fem hern w gang|Rec unil fem hern w gang
C0156117|T020|AB|551.02|ICD9CM|Bilat fem hern w gang|Bilat fem hern w gang
C0156117|T020|PT|551.02|ICD9CM|Femoral hernia with gangrene, bilateral (not specified as recurrent)|Femoral hernia with gangrene, bilateral (not specified as recurrent)
C0156118|T047|PT|551.03|ICD9CM|Femoral hernia with gangrene, bilateral, recurrent|Femoral hernia with gangrene, bilateral, recurrent
C0156118|T047|AB|551.03|ICD9CM|Recur bil fem hern-gang|Recur bil fem hern-gang
C0156119|T047|AB|551.1|ICD9CM|Umbilical hernia w gangr|Umbilical hernia w gangr
C0156119|T047|PT|551.1|ICD9CM|Umbilical hernia with gangrene|Umbilical hernia with gangrene
C0156120|T047|HT|551.2|ICD9CM|Ventral hernia with gangrene|Ventral hernia with gangrene
C0156120|T047|AB|551.20|ICD9CM|Gangr ventral hernia NOS|Gangr ventral hernia NOS
C0156120|T047|PT|551.20|ICD9CM|Ventral hernia, unspecified, with gangrene|Ventral hernia, unspecified, with gangrene
C0156122|T047|AB|551.21|ICD9CM|Gangr incisional hernia|Gangr incisional hernia
C0156122|T047|PT|551.21|ICD9CM|Incisional ventral hernia, with gangrene|Incisional ventral hernia, with gangrene
C0156123|T020|AB|551.29|ICD9CM|Gang ventral hernia NEC|Gang ventral hernia NEC
C0156123|T020|PT|551.29|ICD9CM|Other ventral hernia with gangrene|Other ventral hernia with gangrene
C0156124|T047|AB|551.3|ICD9CM|Diaphragm hernia w gangr|Diaphragm hernia w gangr
C0156124|T047|PT|551.3|ICD9CM|Diaphragmatic hernia with gangrene|Diaphragmatic hernia with gangrene
C0156125|T020|PT|551.8|ICD9CM|Hernia of other specified sites, with gangrene|Hernia of other specified sites, with gangrene
C0156125|T020|AB|551.8|ICD9CM|Hernia, site NEC w gangr|Hernia, site NEC w gangr
C0267667|T047|PT|551.9|ICD9CM|Hernia of unspecified site, with gangrene|Hernia of unspecified site, with gangrene
C0267667|T047|AB|551.9|ICD9CM|Hernia, site NOS w gangr|Hernia, site NOS w gangr
C0156127|T020|HT|552|ICD9CM|Other hernia of abdominal cavity, with obstruction, but without mention of gangrene|Other hernia of abdominal cavity, with obstruction, but without mention of gangrene
C0156128|T020|HT|552.0|ICD9CM|Femoral hernia with obstruction|Femoral hernia with obstruction
C0156129|T020|PT|552.00|ICD9CM|Femoral hernia with obstruction, unilateral or unspecified (not specified as recurrent)|Femoral hernia with obstruction, unilateral or unspecified (not specified as recurrent)
C0156129|T020|AB|552.00|ICD9CM|Unil femoral hern w obst|Unil femoral hern w obst
C0156130|T020|PT|552.01|ICD9CM|Femoral hernia with obstruction, unilateral or unspecified, recurrent|Femoral hernia with obstruction, unilateral or unspecified, recurrent
C0156130|T020|AB|552.01|ICD9CM|Rec unil fem hern w obst|Rec unil fem hern w obst
C0156131|T020|AB|552.02|ICD9CM|Bil femoral hern w obstr|Bil femoral hern w obstr
C0156131|T020|PT|552.02|ICD9CM|Femoral hernia with obstruction, bilateral (not specified as recurrent)|Femoral hernia with obstruction, bilateral (not specified as recurrent)
C3665334|T190|PT|552.03|ICD9CM|Femoral hernia with obstruction, bilateral, recurrent|Femoral hernia with obstruction, bilateral, recurrent
C3665334|T190|AB|552.03|ICD9CM|Rec bil fem hern w obstr|Rec bil fem hern w obstr
C0156133|T020|AB|552.1|ICD9CM|Umbilical hernia w obstr|Umbilical hernia w obstr
C0156133|T020|PT|552.1|ICD9CM|Umbilical hernia with obstruction|Umbilical hernia with obstruction
C1532669|T020|HT|552.2|ICD9CM|Ventral hernia with obstruction|Ventral hernia with obstruction
C1532669|T020|AB|552.20|ICD9CM|Obstr ventral hernia NOS|Obstr ventral hernia NOS
C1532669|T020|PT|552.20|ICD9CM|Ventral, unspecified, hernia with obstruction|Ventral, unspecified, hernia with obstruction
C1442980|T020|PT|552.21|ICD9CM|Incisional ventral hernia with obstruction|Incisional ventral hernia with obstruction
C1442980|T020|AB|552.21|ICD9CM|Obstr incisional hernia|Obstr incisional hernia
C0156137|T020|AB|552.29|ICD9CM|Obstr ventral hernia NEC|Obstr ventral hernia NEC
C0156137|T020|PT|552.29|ICD9CM|Other ventral hernia with obstruction|Other ventral hernia with obstruction
C0700510|T020|AB|552.3|ICD9CM|Diaphragm hernia w obstr|Diaphragm hernia w obstr
C0700510|T020|PT|552.3|ICD9CM|Diaphragmatic hernia with obstruction|Diaphragmatic hernia with obstruction
C0156139|T020|PT|552.8|ICD9CM|Hernia of other specified sites, with obstruction|Hernia of other specified sites, with obstruction
C0156139|T020|AB|552.8|ICD9CM|Hernia, site NEC w obstr|Hernia, site NEC w obstr
C0156140|T020|PT|552.9|ICD9CM|Hernia of unspecified site, with obstruction|Hernia of unspecified site, with obstruction
C0156140|T020|AB|552.9|ICD9CM|Hernia, site NOS w obstr|Hernia, site NOS w obstr
C0156141|T020|HT|553|ICD9CM|Other hernia of abdominal cavity without mention of obstruction or gangrene|Other hernia of abdominal cavity without mention of obstruction or gangrene
C0520569|T020|HT|553.0|ICD9CM|Femoral hernia without mention of obstruction or gangrene|Femoral hernia without mention of obstruction or gangrene
C0041688|T020|AB|553.00|ICD9CM|Unilat femoral hernia|Unilat femoral hernia
C0156142|T020|PT|553.01|ICD9CM|Femoral hernia without mention of obstruction or gangrene, unilateral or unspecified, recurrent|Femoral hernia without mention of obstruction or gangrene, unilateral or unspecified, recurrent
C0156142|T020|AB|553.01|ICD9CM|Recur unil femoral hern|Recur unil femoral hern
C0401094|T020|AB|553.02|ICD9CM|Bilateral femoral hernia|Bilateral femoral hernia
C0401094|T020|PT|553.02|ICD9CM|Femoral hernia without mention of obstruction or gangrene, bilateral (not specified as recurrent)|Femoral hernia without mention of obstruction or gangrene, bilateral (not specified as recurrent)
C0156144|T020|PT|553.03|ICD9CM|Femoral hernia without mention of obstruction or gangrene, bilateral,recurrent|Femoral hernia without mention of obstruction or gangrene, bilateral,recurrent
C0156144|T020|AB|553.03|ICD9CM|Recur bilat femoral hern|Recur bilat femoral hern
C0041636|T020|AB|553.1|ICD9CM|Umbilical hernia|Umbilical hernia
C0041636|T020|PT|553.1|ICD9CM|Umbilical hernia without mention of obstruction or gangrene|Umbilical hernia without mention of obstruction or gangrene
C0042505|T020|HT|553.2|ICD9CM|Ventral hernia without mention of obstruction or gangrene|Ventral hernia without mention of obstruction or gangrene
C0041893|T020|AB|553.20|ICD9CM|Ventral hernia NOS|Ventral hernia NOS
C0041893|T020|PT|553.20|ICD9CM|Ventral, unspecified, hernia without mention of obstruction or gangrene|Ventral, unspecified, hernia without mention of obstruction or gangrene
C0156145|T020|AB|553.21|ICD9CM|Incisional hernia|Incisional hernia
C0156145|T020|PT|553.21|ICD9CM|Incisional hernia without mention of obstruction or gangrene|Incisional hernia without mention of obstruction or gangrene
C0029870|T020|PT|553.29|ICD9CM|Other ventral hernia without mention of obstruction or gangrene|Other ventral hernia without mention of obstruction or gangrene
C0029870|T020|AB|553.29|ICD9CM|Ventral hernia NEC|Ventral hernia NEC
C0494752|T047|AB|553.3|ICD9CM|Diaphragmatic hernia|Diaphragmatic hernia
C0494752|T047|PT|553.3|ICD9CM|Diaphragmatic hernia without mention of obstruction or gangrene|Diaphragmatic hernia without mention of obstruction or gangrene
C0019275|T190|AB|553.8|ICD9CM|Hernia NEC|Hernia NEC
C0019275|T190|PT|553.8|ICD9CM|Hernia of other specified sites without mention of obstruction or gangrene|Hernia of other specified sites without mention of obstruction or gangrene
C0019275|T190|AB|553.9|ICD9CM|Hernia NOS|Hernia NOS
C0019275|T190|PT|553.9|ICD9CM|Hernia of unspecified site without mention of obstruction or gangrene|Hernia of unspecified site without mention of obstruction or gangrene
C0678202|T047|HT|555|ICD9CM|Regional enteritis|Regional enteritis
C0178283|T047|HT|555-558.99|ICD9CM|NONINFECTIOUS ENTERITIS AND COLITIS|NONINFECTIOUS ENTERITIS AND COLITIS
C0156146|T047|AB|555.0|ICD9CM|Reg enteritis, sm intest|Reg enteritis, sm intest
C0156146|T047|PT|555.0|ICD9CM|Regional enteritis of small intestine|Regional enteritis of small intestine
C0156147|T047|AB|555.1|ICD9CM|Reg enteritis, lg intest|Reg enteritis, lg intest
C0156147|T047|PT|555.1|ICD9CM|Regional enteritis of large intestine|Regional enteritis of large intestine
C0267383|T047|AB|555.2|ICD9CM|Reg enterit sm/lg intest|Reg enterit sm/lg intest
C0267383|T047|PT|555.2|ICD9CM|Regional enteritis of small intestine with large intestine|Regional enteritis of small intestine with large intestine
C0678202|T047|AB|555.9|ICD9CM|Regional enteritis NOS|Regional enteritis NOS
C0678202|T047|PT|555.9|ICD9CM|Regional enteritis of unspecified site|Regional enteritis of unspecified site
C0009324|T047|HT|556|ICD9CM|Ulcerative colitis|Ulcerative colitis
C0267388|T047|PT|556.0|ICD9CM|Ulcerative (chronic) enterocolitis|Ulcerative (chronic) enterocolitis
C0267388|T047|AB|556.0|ICD9CM|Ulcerative enterocolitis|Ulcerative enterocolitis
C0267389|T047|PT|556.1|ICD9CM|Ulcerative (chronic) ileocolitis|Ulcerative (chronic) ileocolitis
C0267389|T047|AB|556.1|ICD9CM|Ulcerative ileocolitis|Ulcerative ileocolitis
C2937222|T047|PT|556.2|ICD9CM|Ulcerative (chronic) proctitis|Ulcerative (chronic) proctitis
C2937222|T047|AB|556.2|ICD9CM|Ulcerative proctitis|Ulcerative proctitis
C0267390|T047|PT|556.3|ICD9CM|Ulcerative (chronic) proctosigmoiditis|Ulcerative (chronic) proctosigmoiditis
C0267390|T047|AB|556.3|ICD9CM|Ulcertve prctosigmoidtis|Ulcertve prctosigmoidtis
C0267392|T047|AB|556.4|ICD9CM|Pseudopolyposis colon|Pseudopolyposis colon
C0267392|T047|PT|556.4|ICD9CM|Pseudopolyposis of colon|Pseudopolyposis of colon
C0375359|T047|PT|556.5|ICD9CM|Left-sided ulcerative (chronic) colitis|Left-sided ulcerative (chronic) colitis
C0375359|T047|AB|556.5|ICD9CM|Lftsded ulcertve colitis|Lftsded ulcertve colitis
C0375360|T047|PT|556.6|ICD9CM|Universal ulcerative (chronic) colitis|Universal ulcerative (chronic) colitis
C0375360|T047|AB|556.6|ICD9CM|Univrsl ulcertve colitis|Univrsl ulcertve colitis
C0348737|T047|AB|556.8|ICD9CM|Other ulcerative colitis|Other ulcerative colitis
C0348737|T047|PT|556.8|ICD9CM|Other ulcerative colitis|Other ulcerative colitis
C0009324|T047|PT|556.9|ICD9CM|Ulcerative colitis, unspecified|Ulcerative colitis, unspecified
C0009324|T047|AB|556.9|ICD9CM|Ulceratve colitis unspcf|Ulceratve colitis unspcf
C2004435|T047|HT|557|ICD9CM|Vascular insufficiency of intestine|Vascular insufficiency of intestine
C0001363|T047|AB|557.0|ICD9CM|Ac vasc insuff intestine|Ac vasc insuff intestine
C0001363|T047|PT|557.0|ICD9CM|Acute vascular insufficiency of intestine|Acute vascular insufficiency of intestine
C0311262|T047|AB|557.1|ICD9CM|Chr vasc insuff intest|Chr vasc insuff intest
C0311262|T047|PT|557.1|ICD9CM|Chronic vascular insufficiency of intestine|Chronic vascular insufficiency of intestine
C2004435|T047|PT|557.9|ICD9CM|Unspecified vascular insufficiency of intestine|Unspecified vascular insufficiency of intestine
C2004435|T047|AB|557.9|ICD9CM|Vasc insuff intest NOS|Vasc insuff intest NOS
C0029512|T047|HT|558|ICD9CM|Other and unspecified noninfectious gastroenteritis and colitis|Other and unspecified noninfectious gastroenteritis and colitis
C0156153|T047|PT|558.1|ICD9CM|Gastroenteritis and colitis due to radiation|Gastroenteritis and colitis due to radiation
C0156153|T047|AB|558.1|ICD9CM|Radiation gastroenterit|Radiation gastroenterit
C0156154|T047|AB|558.2|ICD9CM|Toxic gastroenteritis|Toxic gastroenteritis
C0156154|T047|PT|558.2|ICD9CM|Toxic gastroenteritis and colitis|Toxic gastroenteritis and colitis
C0401143|T047|PT|558.3|ICD9CM|Allergic gastroenteritis and colitis|Allergic gastroenteritis and colitis
C0401143|T047|AB|558.3|ICD9CM|Allrgic gastro & colitis|Allrgic gastro & colitis
C2349567|T047|HT|558.4|ICD9CM|Eosinophilic gastroenteritis and colitis|Eosinophilic gastroenteritis and colitis
C1262481|T047|AB|558.41|ICD9CM|Eosinophilic gastroent|Eosinophilic gastroent
C1262481|T047|PT|558.41|ICD9CM|Eosinophilic gastroenteritis|Eosinophilic gastroenteritis
C0267448|T047|PT|558.42|ICD9CM|Eosinophilic colitis|Eosinophilic colitis
C0267448|T047|AB|558.42|ICD9CM|Eosinophilic colitis|Eosinophilic colitis
C0029512|T047|AB|558.9|ICD9CM|Noninf gastroenterit NEC|Noninf gastroenterit NEC
C0029512|T047|PT|558.9|ICD9CM|Other and unspecified noninfectious gastroenteritis and colitis|Other and unspecified noninfectious gastroenteritis and colitis
C0021844|T020|HT|560|ICD9CM|Intestinal obstruction without mention of hernia|Intestinal obstruction without mention of hernia
C0178284|T047|HT|560-569.99|ICD9CM|OTHER DISEASES OF INTESTINES AND PERITONEUM|OTHER DISEASES OF INTESTINES AND PERITONEUM
C0021933|T047|AB|560.0|ICD9CM|Intussusception|Intussusception
C0021933|T047|PT|560.0|ICD9CM|Intussusception|Intussusception
C0030446|T047|AB|560.1|ICD9CM|Paralytic ileus|Paralytic ileus
C0030446|T047|PT|560.1|ICD9CM|Paralytic ileus|Paralytic ileus
C0042961|T047|PT|560.2|ICD9CM|Volvulus|Volvulus
C0042961|T047|AB|560.2|ICD9CM|Volvulus of intestine|Volvulus of intestine
C0392503|T033|HT|560.3|ICD9CM|Impaction of intestine|Impaction of intestine
C0392503|T033|AB|560.30|ICD9CM|Impaction intestine NOS|Impaction intestine NOS
C0392503|T033|PT|560.30|ICD9CM|Impaction of intestine, unspecified|Impaction of intestine, unspecified
C0156156|T047|AB|560.31|ICD9CM|Gallstone ileus|Gallstone ileus
C0156156|T047|PT|560.31|ICD9CM|Gallstone ileus|Gallstone ileus
C0015734|T033|PT|560.32|ICD9CM|Fecal impaction|Fecal impaction
C0015734|T033|AB|560.32|ICD9CM|Fecal impaction|Fecal impaction
C0029640|T047|AB|560.39|ICD9CM|Impaction intestine NEC|Impaction intestine NEC
C0029640|T047|PT|560.39|ICD9CM|Other impaction of intestine|Other impaction of intestine
C0156157|T047|HT|560.8|ICD9CM|Other specified intestinal obstruction|Other specified intestinal obstruction
C0156158|T047|AB|560.81|ICD9CM|Intestinal adhes w obstr|Intestinal adhes w obstr
C0156158|T047|PT|560.81|ICD9CM|Intestinal or peritoneal adhesions with obstruction (postoperative) (postinfection)|Intestinal or peritoneal adhesions with obstruction (postoperative) (postinfection)
C0156157|T047|AB|560.89|ICD9CM|Intestinal obstruct NEC|Intestinal obstruct NEC
C0156157|T047|PT|560.89|ICD9CM|Other specified intestinal obstruction|Other specified intestinal obstruction
C0021843|T047|AB|560.9|ICD9CM|Intestinal obstruct NOS|Intestinal obstruct NOS
C0021843|T047|PT|560.9|ICD9CM|Unspecified intestinal obstruction|Unspecified intestinal obstruction
C1510475|T047|HT|562|ICD9CM|Diverticula of intestine|Diverticula of intestine
C0267498|T047|HT|562.0|ICD9CM|Diverticula of small intestine|Diverticula of small intestine
C0156162|T047|PT|562.00|ICD9CM|Diverticulosis of small intestine (without mention of hemorrhage)|Diverticulosis of small intestine (without mention of hemorrhage)
C0156162|T047|AB|562.00|ICD9CM|Dvrtclo sml int w/o hmrg|Dvrtclo sml int w/o hmrg
C0156163|T047|PT|562.01|ICD9CM|Diverticulitis of small intestine (without mention of hemorrhage)|Diverticulitis of small intestine (without mention of hemorrhage)
C0156163|T047|AB|562.01|ICD9CM|Dvrtcli sml int w/o hmrg|Dvrtcli sml int w/o hmrg
C4038618|T047|PT|562.02|ICD9CM|Diverticulosis of small intestine with hemorrhage|Diverticulosis of small intestine with hemorrhage
C4038618|T047|AB|562.02|ICD9CM|Dvrtclo sml int w hmrhg|Dvrtclo sml int w hmrhg
C0156165|T047|PT|562.03|ICD9CM|Diverticulitis of small intestine with hemorrhage|Diverticulitis of small intestine with hemorrhage
C0156165|T047|AB|562.03|ICD9CM|Dvrtcli sml int w hmrhg|Dvrtcli sml int w hmrhg
C0012811|T190|HT|562.1|ICD9CM|Diverticula of colon|Diverticula of colon
C0156166|T047|PT|562.10|ICD9CM|Diverticulosis of colon (without mention of hemorrhage)|Diverticulosis of colon (without mention of hemorrhage)
C0156166|T047|AB|562.10|ICD9CM|Dvrtclo colon w/o hmrhg|Dvrtclo colon w/o hmrhg
C0156167|T047|PT|562.11|ICD9CM|Diverticulitis of colon (without mention of hemorrhage)|Diverticulitis of colon (without mention of hemorrhage)
C0156167|T047|AB|562.11|ICD9CM|Dvrtcli colon w/o hmrhg|Dvrtcli colon w/o hmrhg
C0156168|T047|PT|562.12|ICD9CM|Diverticulosis of colon with hemorrhage|Diverticulosis of colon with hemorrhage
C0156168|T047|AB|562.12|ICD9CM|Dvrtclo colon w hmrhg|Dvrtclo colon w hmrhg
C0544793|T047|PT|562.13|ICD9CM|Diverticulitis of colon with hemorrhage|Diverticulitis of colon with hemorrhage
C0544793|T047|AB|562.13|ICD9CM|Dvrtcli colon w hmrhg|Dvrtcli colon w hmrhg
C0302382|T047|HT|564|ICD9CM|Functional digestive disorders, not elsewhere classified|Functional digestive disorders, not elsewhere classified
C0009806|T184|HT|564.0|ICD9CM|Constipation|Constipation
C0009806|T184|AB|564.00|ICD9CM|Constipation NOS|Constipation NOS
C0009806|T184|PT|564.00|ICD9CM|Constipation, unspecified|Constipation, unspecified
C0729262|T033|PT|564.01|ICD9CM|Slow transit constipation|Slow transit constipation
C0729262|T033|AB|564.01|ICD9CM|Slow transt constipation|Slow transt constipation
C0949134|T047|AB|564.02|ICD9CM|Outlet dysfnc constption|Outlet dysfnc constption
C0949134|T047|PT|564.02|ICD9CM|Outlet dysfunction constipation|Outlet dysfunction constipation
C0949135|T047|AB|564.09|ICD9CM|Constipation NEC|Constipation NEC
C0949135|T047|PT|564.09|ICD9CM|Other constipation|Other constipation
C0022104|T047|AB|564.1|ICD9CM|Irritable bowel syndrome|Irritable bowel syndrome
C0022104|T047|PT|564.1|ICD9CM|Irritable bowel syndrome|Irritable bowel syndrome
C0032763|T047|AB|564.2|ICD9CM|Postgastric surgery synd|Postgastric surgery synd
C0032763|T047|PT|564.2|ICD9CM|Postgastric surgery syndromes|Postgastric surgery syndromes
C0156171|T184|PT|564.3|ICD9CM|Vomiting following gastrointestinal surgery|Vomiting following gastrointestinal surgery
C0156171|T184|AB|564.3|ICD9CM|Vomiting post-gi surgery|Vomiting post-gi surgery
C0156172|T047|PT|564.4|ICD9CM|Other postoperative functional disorders|Other postoperative functional disorders
C0156172|T047|AB|564.4|ICD9CM|Postop GI funct dis NEC|Postop GI funct dis NEC
C0156173|T047|AB|564.5|ICD9CM|Functional diarrhea|Functional diarrhea
C0156173|T047|PT|564.5|ICD9CM|Functional diarrhea|Functional diarrhea
C0152167|T047|AB|564.6|ICD9CM|Anal spasm|Anal spasm
C0152167|T047|PT|564.6|ICD9CM|Anal spasm|Anal spasm
C0235904|T047|AB|564.7|ICD9CM|Megacolon NEC|Megacolon NEC
C0235904|T047|PT|564.7|ICD9CM|Megacolon, other than Hirschsprung's|Megacolon, other than Hirschsprung's
C0494776|T047|HT|564.8|ICD9CM|Other specified functional disorders of intestine|Other specified functional disorders of intestine
C0695242|T047|AB|564.81|ICD9CM|Neurogenic bowel|Neurogenic bowel
C0695242|T047|PT|564.81|ICD9CM|Neurogenic bowel|Neurogenic bowel
C0341089|T047|AB|564.89|ICD9CM|Funct dis intestine NEC|Funct dis intestine NEC
C0341089|T047|PT|564.89|ICD9CM|Other functional disorders of intestine|Other functional disorders of intestine
C0016807|T047|AB|564.9|ICD9CM|Funct dis intestine NOS|Funct dis intestine NOS
C0016807|T047|PT|564.9|ICD9CM|Unspecified functional disorder of intestine|Unspecified functional disorder of intestine
C0156175|T190|HT|565|ICD9CM|Anal fissure and fistula|Anal fissure and fistula
C0016167|T047|AB|565.0|ICD9CM|Anal fissure|Anal fissure
C0016167|T047|PT|565.0|ICD9CM|Anal fissure|Anal fissure
C0205929|T020|AB|565.1|ICD9CM|Anal fistula|Anal fistula
C0205929|T020|PT|565.1|ICD9CM|Anal fistula|Anal fistula
C0267567|T047|PT|566|ICD9CM|Abscess of anal and rectal regions|Abscess of anal and rectal regions
C0267567|T047|AB|566|ICD9CM|Anal & rectal abscess|Anal & rectal abscess
C1561637|T047|HT|567|ICD9CM|Peritonitis and retroperitoneal infections|Peritonitis and retroperitoneal infections
C0156177|T047|AB|567.0|ICD9CM|Peritonitis in infec dis|Peritonitis in infec dis
C0156177|T047|PT|567.0|ICD9CM|Peritonitis in infectious diseases classified elsewhere|Peritonitis in infectious diseases classified elsewhere
C0156178|T047|AB|567.1|ICD9CM|Pneumococcal peritonitis|Pneumococcal peritonitis
C0156178|T047|PT|567.1|ICD9CM|Pneumococcal peritonitis|Pneumococcal peritonitis
C0156179|T047|HT|567.2|ICD9CM|Other suppurative peritonitis|Other suppurative peritonitis
C0267751|T047|AB|567.21|ICD9CM|Peritonitis (acute) gen|Peritonitis (acute) gen
C0267751|T047|PT|567.21|ICD9CM|Peritonitis (acute) generalized|Peritonitis (acute) generalized
C0267756|T047|AB|567.22|ICD9CM|Peritoneal abscess|Peritoneal abscess
C0267756|T047|PT|567.22|ICD9CM|Peritoneal abscess|Peritoneal abscess
C0275551|T047|AB|567.23|ICD9CM|Spontan bact peritonitis|Spontan bact peritonitis
C0275551|T047|PT|567.23|ICD9CM|Spontaneous bacterial peritonitis|Spontaneous bacterial peritonitis
C0156179|T047|PT|567.29|ICD9CM|Other suppurative peritonitis|Other suppurative peritonitis
C0156179|T047|AB|567.29|ICD9CM|Suppurat peritonitis NEC|Suppurat peritonitis NEC
C0920049|T047|HT|567.3|ICD9CM|Retroperitoneal infections|Retroperitoneal infections
C0085222|T047|AB|567.31|ICD9CM|Psoas muscle abscess|Psoas muscle abscess
C0085222|T047|PT|567.31|ICD9CM|Psoas muscle abscess|Psoas muscle abscess
C1561633|T046|PT|567.38|ICD9CM|Other retroperitoneal abscess|Other retroperitoneal abscess
C1561633|T046|AB|567.38|ICD9CM|Retroperiton abscess NEC|Retroperiton abscess NEC
C1561634|T047|PT|567.39|ICD9CM|Other retroperitoneal infections|Other retroperitoneal infections
C1561634|T047|AB|567.39|ICD9CM|Retroperiton infect NEC|Retroperiton infect NEC
C0029823|T047|HT|567.8|ICD9CM|Other specified peritonitis|Other specified peritonitis
C0267768|T047|AB|567.81|ICD9CM|Choleperitonitis|Choleperitonitis
C0267768|T047|PT|567.81|ICD9CM|Choleperitonitis|Choleperitonitis
C0267770|T047|AB|567.82|ICD9CM|Sclerosing mesenteritis|Sclerosing mesenteritis
C0267770|T047|PT|567.82|ICD9CM|Sclerosing mesenteritis|Sclerosing mesenteritis
C0029823|T047|PT|567.89|ICD9CM|Other specified peritonitis|Other specified peritonitis
C0029823|T047|AB|567.89|ICD9CM|Peritonitis NEC|Peritonitis NEC
C0031154|T046|AB|567.9|ICD9CM|Peritonitis NOS|Peritonitis NOS
C0031154|T046|PT|567.9|ICD9CM|Unspecified peritonitis|Unspecified peritonitis
C0156180|T047|HT|568|ICD9CM|Other disorders of peritoneum|Other disorders of peritoneum
C0375362|T047|AB|568.0|ICD9CM|Peritoneal adhesions|Peritoneal adhesions
C0375362|T047|PT|568.0|ICD9CM|Peritoneal adhesions (postoperative) (postinfection)|Peritoneal adhesions (postoperative) (postinfection)
C0029786|T047|HT|568.8|ICD9CM|Other specified disorders of peritoneum|Other specified disorders of peritoneum
C0019066|T046|AB|568.81|ICD9CM|Hemoperitoneum|Hemoperitoneum
C0019066|T046|PT|568.81|ICD9CM|Hemoperitoneum (nontraumatic)|Hemoperitoneum (nontraumatic)
C0031144|T047|AB|568.82|ICD9CM|Peritoneal effusion|Peritoneal effusion
C0031144|T047|PT|568.82|ICD9CM|Peritoneal effusion (chronic)|Peritoneal effusion (chronic)
C0029786|T047|PT|568.89|ICD9CM|Other specified disorders of peritoneum|Other specified disorders of peritoneum
C0029786|T047|AB|568.89|ICD9CM|Peritoneal disorder NEC|Peritoneal disorder NEC
C0031142|T047|AB|568.9|ICD9CM|Peritoneal disorder NOS|Peritoneal disorder NOS
C0031142|T047|PT|568.9|ICD9CM|Unspecified disorder of peritoneum|Unspecified disorder of peritoneum
C0156182|T047|HT|569|ICD9CM|Other disorders of intestine|Other disorders of intestine
C0002753|T020|AB|569.0|ICD9CM|Anal & rectal polyp|Anal & rectal polyp
C0002753|T020|PT|569.0|ICD9CM|Anal and rectal polyp|Anal and rectal polyp
C0034888|T047|AB|569.1|ICD9CM|Rectal prolapse|Rectal prolapse
C0034888|T047|PT|569.1|ICD9CM|Rectal prolapse|Rectal prolapse
C0156183|T190|AB|569.2|ICD9CM|Rectal & anal stenosis|Rectal & anal stenosis
C0156183|T190|PT|569.2|ICD9CM|Stenosis of rectum and anus|Stenosis of rectum and anus
C0019081|T046|PT|569.3|ICD9CM|Hemorrhage of rectum and anus|Hemorrhage of rectum and anus
C0019081|T046|AB|569.3|ICD9CM|Rectal & anal hemorrhage|Rectal & anal hemorrhage
C0348742|T047|HT|569.4|ICD9CM|Other specified disorders of rectum and anus|Other specified disorders of rectum and anus
C0400832|T047|AB|569.41|ICD9CM|Rectal & anal ulcer|Rectal & anal ulcer
C0400832|T047|PT|569.41|ICD9CM|Ulcer of anus and rectum|Ulcer of anus and rectum
C0002758|T184|AB|569.42|ICD9CM|Anal or rectal pain|Anal or rectal pain
C0002758|T184|PT|569.42|ICD9CM|Anal or rectal pain|Anal or rectal pain
C1955814|T047|PT|569.43|ICD9CM|Anal sphincter tear (healed) (old)|Anal sphincter tear (healed) (old)
C1955814|T047|AB|569.43|ICD9CM|Anal sphincter tear-old|Anal sphincter tear-old
C0347129|T191|PT|569.44|ICD9CM|Dysplasia of anus|Dysplasia of anus
C0347129|T191|AB|569.44|ICD9CM|Dysplasia of anus|Dysplasia of anus
C0348742|T047|PT|569.49|ICD9CM|Other specified disorders of rectum and anus|Other specified disorders of rectum and anus
C0348742|T047|AB|569.49|ICD9CM|Rectal & anal dis NEC|Rectal & anal dis NEC
C0156185|T047|PT|569.5|ICD9CM|Abscess of intestine|Abscess of intestine
C0156185|T047|AB|569.5|ICD9CM|Intestinal abscess|Intestinal abscess
C0156186|T046|HT|569.6|ICD9CM|Colostomy and enterostomy complications|Colostomy and enterostomy complications
C0156186|T046|PT|569.60|ICD9CM|Colostomy and enterostomy complication, unspecified|Colostomy and enterostomy complication, unspecified
C0156186|T046|AB|569.60|ICD9CM|Colstomy/enter comp NOS|Colstomy/enter comp NOS
C0375363|T047|AB|569.61|ICD9CM|Colosty/enterost infectn|Colosty/enterost infectn
C0375363|T047|PT|569.61|ICD9CM|Infection of colostomy or enterostomy|Infection of colostomy or enterostomy
C0695243|T046|AB|569.62|ICD9CM|Colosty/enter comp-mech|Colosty/enter comp-mech
C0695243|T046|PT|569.62|ICD9CM|Mechanical complication of colostomy and enterostomy|Mechanical complication of colostomy and enterostomy
C0375364|T047|AB|569.69|ICD9CM|Colstmy/enteros comp NEC|Colstmy/enteros comp NEC
C0375364|T047|PT|569.69|ICD9CM|Other colostomy and enterostomy complication|Other colostomy and enterostomy complication
C2712967|T046|HT|569.7|ICD9CM|Complications of intestinal pouch|Complications of intestinal pouch
C0376620|T047|AB|569.71|ICD9CM|Pouchitis|Pouchitis
C0376620|T047|PT|569.71|ICD9CM|Pouchitis|Pouchitis
C2712860|T046|AB|569.79|ICD9CM|Comp intest pouch NEC|Comp intest pouch NEC
C2712860|T046|PT|569.79|ICD9CM|Other complications of intestinal pouch|Other complications of intestinal pouch
C0348743|T047|HT|569.8|ICD9CM|Other specified disorders of intestine|Other specified disorders of intestine
C0016171|T190|PT|569.81|ICD9CM|Fistula of intestine, excluding rectum and anus|Fistula of intestine, excluding rectum and anus
C0016171|T190|AB|569.81|ICD9CM|Intestinal fistula|Intestinal fistula
C0151971|T047|AB|569.82|ICD9CM|Ulceration of intestine|Ulceration of intestine
C0151971|T047|PT|569.82|ICD9CM|Ulceration of intestine|Ulceration of intestine
C0021845|T047|AB|569.83|ICD9CM|Perforation of intestine|Perforation of intestine
C0021845|T047|PT|569.83|ICD9CM|Perforation of intestine|Perforation of intestine
C0267367|T047|AB|569.84|ICD9CM|Angio intes w/o hmrhg|Angio intes w/o hmrhg
C0267367|T047|PT|569.84|ICD9CM|Angiodysplasia of intestine (without mention of hemorrhage)|Angiodysplasia of intestine (without mention of hemorrhage)
C0156188|T047|AB|569.85|ICD9CM|Angio intes w hmrhg|Angio intes w hmrhg
C0156188|T047|PT|569.85|ICD9CM|Angiodysplasia of intestine with hemorrhage|Angiodysplasia of intestine with hemorrhage
C2183395|T047|AB|569.86|ICD9CM|Dieulafoy les, intestine|Dieulafoy les, intestine
C2183395|T047|PT|569.86|ICD9CM|Dieulafoy lesion (hemorrhagic) of intestine|Dieulafoy lesion (hemorrhagic) of intestine
C3874311|T047|PT|569.87|ICD9CM|Vomiting of fecal matter|Vomiting of fecal matter
C3874311|T047|AB|569.87|ICD9CM|Vomiting of fecal matter|Vomiting of fecal matter
C0348743|T047|AB|569.89|ICD9CM|Intestinal disorders NEC|Intestinal disorders NEC
C0348743|T047|PT|569.89|ICD9CM|Other specified disorders of intestine|Other specified disorders of intestine
C0021831|T047|AB|569.9|ICD9CM|Intestinal disorder NOS|Intestinal disorder NOS
C0021831|T047|PT|569.9|ICD9CM|Unspecified disorder of intestine|Unspecified disorder of intestine
C0001308|T047|PT|570|ICD9CM|Acute and subacute necrosis of liver|Acute and subacute necrosis of liver
C0001308|T047|AB|570|ICD9CM|Acute necrosis of liver|Acute necrosis of liver
C0178285|T047|HT|570-579.99|ICD9CM|OTHER DISEASES OF DIGESTIVE SYSTEM|OTHER DISEASES OF DIGESTIVE SYSTEM
C0156189|T047|HT|571|ICD9CM|Chronic liver disease and cirrhosis|Chronic liver disease and cirrhosis
C0015696|T047|AB|571.0|ICD9CM|Alcoholic fatty liver|Alcoholic fatty liver
C0015696|T047|PT|571.0|ICD9CM|Alcoholic fatty liver|Alcoholic fatty liver
C0001306|T047|AB|571.1|ICD9CM|Ac alcoholic hepatitis|Ac alcoholic hepatitis
C0001306|T047|PT|571.1|ICD9CM|Acute alcoholic hepatitis|Acute alcoholic hepatitis
C0023891|T047|AB|571.2|ICD9CM|Alcohol cirrhosis liver|Alcohol cirrhosis liver
C0023891|T047|PT|571.2|ICD9CM|Alcoholic cirrhosis of liver|Alcoholic cirrhosis of liver
C1442981|T047|AB|571.3|ICD9CM|Alcohol liver damage NOS|Alcohol liver damage NOS
C1442981|T047|PT|571.3|ICD9CM|Alcoholic liver damage, unspecified|Alcoholic liver damage, unspecified
C0019189|T047|HT|571.4|ICD9CM|Chronic hepatitis|Chronic hepatitis
C0019189|T047|AB|571.40|ICD9CM|Chronic hepatitis NOS|Chronic hepatitis NOS
C0019189|T047|PT|571.40|ICD9CM|Chronic hepatitis, unspecified|Chronic hepatitis, unspecified
C0149519|T047|AB|571.41|ICD9CM|Chr persistent hepatitis|Chr persistent hepatitis
C0149519|T047|PT|571.41|ICD9CM|Chronic persistent hepatitis|Chronic persistent hepatitis
C0241910|T047|AB|571.42|ICD9CM|Autoimmune hepatitis|Autoimmune hepatitis
C0241910|T047|PT|571.42|ICD9CM|Autoimmune hepatitis|Autoimmune hepatitis
C0029545|T047|AB|571.49|ICD9CM|Chronic hepatitis NEC|Chronic hepatitis NEC
C0029545|T047|PT|571.49|ICD9CM|Other chronic hepatitis|Other chronic hepatitis
C0008827|T047|AB|571.5|ICD9CM|Cirrhosis of liver NOS|Cirrhosis of liver NOS
C0008827|T047|PT|571.5|ICD9CM|Cirrhosis of liver without mention of alcohol|Cirrhosis of liver without mention of alcohol
C0023892|T047|AB|571.6|ICD9CM|Biliary cirrhosis|Biliary cirrhosis
C0023892|T047|PT|571.6|ICD9CM|Biliary cirrhosis|Biliary cirrhosis
C0029546|T047|AB|571.8|ICD9CM|Chronic liver dis NEC|Chronic liver dis NEC
C0029546|T047|PT|571.8|ICD9CM|Other chronic nonalcoholic liver disease|Other chronic nonalcoholic liver disease
C0687718|T047|AB|571.9|ICD9CM|Chronic liver dis NOS|Chronic liver dis NOS
C0687718|T047|PT|571.9|ICD9CM|Unspecified chronic liver disease without mention of alcohol|Unspecified chronic liver disease without mention of alcohol
C0156191|T047|HT|572|ICD9CM|Liver abscess and sequelae of chronic liver disease|Liver abscess and sequelae of chronic liver disease
C0023885|T047|AB|572.0|ICD9CM|Abscess of liver|Abscess of liver
C0023885|T047|PT|572.0|ICD9CM|Abscess of liver|Abscess of liver
C0156192|T047|AB|572.1|ICD9CM|Portal pyemia|Portal pyemia
C0156192|T047|PT|572.1|ICD9CM|Portal pyemia|Portal pyemia
C0019151|T047|PT|572.2|ICD9CM|Hepatic encephalopathy|Hepatic encephalopathy
C0019151|T047|AB|572.2|ICD9CM|Hepatic encephalopathy|Hepatic encephalopathy
C0020541|T047|AB|572.3|ICD9CM|Portal hypertension|Portal hypertension
C0020541|T047|PT|572.3|ICD9CM|Portal hypertension|Portal hypertension
C0019212|T047|AB|572.4|ICD9CM|Hepatorenal syndrome|Hepatorenal syndrome
C0019212|T047|PT|572.4|ICD9CM|Hepatorenal syndrome|Hepatorenal syndrome
C0156193|T047|AB|572.8|ICD9CM|Oth sequela, chr liv dis|Oth sequela, chr liv dis
C0156193|T047|PT|572.8|ICD9CM|Other sequelae of chronic liver disease|Other sequelae of chronic liver disease
C0156194|T047|HT|573|ICD9CM|Other disorders of liver|Other disorders of liver
C0156195|T047|AB|573.0|ICD9CM|Chr passiv congest liver|Chr passiv congest liver
C0156195|T047|PT|573.0|ICD9CM|Chronic passive congestion of liver|Chronic passive congestion of liver
C0156196|T047|AB|573.1|ICD9CM|Hepatitis in viral dis|Hepatitis in viral dis
C0156196|T047|PT|573.1|ICD9CM|Hepatitis in viral diseases classified elsewhere|Hepatitis in viral diseases classified elsewhere
C0156197|T047|AB|573.2|ICD9CM|Hepatitis in oth inf dis|Hepatitis in oth inf dis
C0156197|T047|PT|573.2|ICD9CM|Hepatitis in other infectious diseases classified elsewhere|Hepatitis in other infectious diseases classified elsewhere
C0019158|T047|AB|573.3|ICD9CM|Hepatitis NOS|Hepatitis NOS
C0019158|T047|PT|573.3|ICD9CM|Hepatitis, unspecified|Hepatitis, unspecified
C0151731|T047|AB|573.4|ICD9CM|Hepatic infarction|Hepatic infarction
C0151731|T047|PT|573.4|ICD9CM|Hepatic infarction|Hepatic infarction
C0600452|T047|PT|573.5|ICD9CM|Hepatopulmonary syndrome|Hepatopulmonary syndrome
C0600452|T047|AB|573.5|ICD9CM|Hepatopulmonary syndrome|Hepatopulmonary syndrome
C0348751|T047|AB|573.8|ICD9CM|Liver disorders NEC|Liver disorders NEC
C0348751|T047|PT|573.8|ICD9CM|Other specified disorders of liver|Other specified disorders of liver
C0023895|T047|AB|573.9|ICD9CM|Liver disorder NOS|Liver disorder NOS
C0023895|T047|PT|573.9|ICD9CM|Unspecified disorder of liver|Unspecified disorder of liver
C0008350|T047|HT|574|ICD9CM|Cholelithiasis|Cholelithiasis
C0156199|T047|HT|574.0|ICD9CM|Calculus of gallbladder with acute cholecystitis|Calculus of gallbladder with acute cholecystitis
C0400985|T047|PT|574.00|ICD9CM|Calculus of gallbladder with acute cholecystitis, without mention of obstruction|Calculus of gallbladder with acute cholecystitis, without mention of obstruction
C0400985|T047|AB|574.00|ICD9CM|Cholelith w ac cholecyst|Cholelith w ac cholecyst
C0156201|T047|PT|574.01|ICD9CM|Calculus of gallbladder with acute cholecystitis, with obstruction|Calculus of gallbladder with acute cholecystitis, with obstruction
C0156201|T047|AB|574.01|ICD9CM|Cholelith/ac gb inf-obst|Cholelith/ac gb inf-obst
C0156202|T047|HT|574.1|ICD9CM|Calculus of gallbladder with other cholecystitis|Calculus of gallbladder with other cholecystitis
C0156203|T047|PT|574.10|ICD9CM|Calculus of gallbladder with other cholecystitis, without mention of obstruction|Calculus of gallbladder with other cholecystitis, without mention of obstruction
C0156203|T047|AB|574.10|ICD9CM|Cholelith w cholecys NEC|Cholelith w cholecys NEC
C0156204|T047|PT|574.11|ICD9CM|Calculus of gallbladder with other cholecystitis, with obstruction|Calculus of gallbladder with other cholecystitis, with obstruction
C0156204|T047|AB|574.11|ICD9CM|Cholelith/gb inf NEC-obs|Cholelith/gb inf NEC-obs
C0006741|T047|HT|574.2|ICD9CM|Calculus of gallbladder without mention of cholecystitis|Calculus of gallbladder without mention of cholecystitis
C0006742|T047|PT|574.20|ICD9CM|Calculus of gallbladder without mention of cholecystitis, without mention of obstruction|Calculus of gallbladder without mention of cholecystitis, without mention of obstruction
C0006742|T047|AB|574.20|ICD9CM|Cholelithiasis NOS|Cholelithiasis NOS
C0156205|T047|PT|574.21|ICD9CM|Calculus of gallbladder without mention of cholecystitis, with obstruction|Calculus of gallbladder without mention of cholecystitis, with obstruction
C0156205|T047|AB|574.21|ICD9CM|Cholelithias NOS w obstr|Cholelithias NOS w obstr
C0156206|T047|HT|574.3|ICD9CM|Calculus of bile duct with acute cholecystitis|Calculus of bile duct with acute cholecystitis
C0156207|T047|PT|574.30|ICD9CM|Calculus of bile duct with acute cholecystitis, without mention of obstruction|Calculus of bile duct with acute cholecystitis, without mention of obstruction
C0156207|T047|AB|574.30|ICD9CM|Choledocholith/ac gb inf|Choledocholith/ac gb inf
C0156208|T047|PT|574.31|ICD9CM|Calculus of bile duct with acute cholecystitis, with obstruction|Calculus of bile duct with acute cholecystitis, with obstruction
C0156208|T047|AB|574.31|ICD9CM|Choledochlith/ac gb-obst|Choledochlith/ac gb-obst
C0156209|T047|HT|574.4|ICD9CM|Calculus of bile duct with other cholecystitis|Calculus of bile duct with other cholecystitis
C0156210|T047|PT|574.40|ICD9CM|Calculus of bile duct with other cholecystitis, without mention of obstruction|Calculus of bile duct with other cholecystitis, without mention of obstruction
C0156210|T047|AB|574.40|ICD9CM|Choledochlith/gb inf NEC|Choledochlith/gb inf NEC
C0156211|T047|PT|574.41|ICD9CM|Calculus of bile duct with other cholecystitis, with obstruction|Calculus of bile duct with other cholecystitis, with obstruction
C0156211|T047|AB|574.41|ICD9CM|Choledochlith/gb NEC-obs|Choledochlith/gb NEC-obs
C0006739|T047|HT|574.5|ICD9CM|Calculus of bile duct without mention of cholecystitis|Calculus of bile duct without mention of cholecystitis
C0156212|T047|PT|574.50|ICD9CM|Calculus of bile duct without mention of cholecystitis, without mention of obstruction|Calculus of bile duct without mention of cholecystitis, without mention of obstruction
C0156212|T047|AB|574.50|ICD9CM|Choledocholithiasis NOS|Choledocholithiasis NOS
C0375365|T047|HT|574.6|ICD9CM|Calculus of gallbladder and bile duct with acute cholecystitis|Calculus of gallbladder and bile duct with acute cholecystitis
C0375366|T047|PT|574.60|ICD9CM|Calculus of gallbladder and bile duct with acute cholecystitis, without mention of obstruction|Calculus of gallbladder and bile duct with acute cholecystitis, without mention of obstruction
C0375366|T047|AB|574.60|ICD9CM|Gall&bil cal w/ac w/o ob|Gall&bil cal w/ac w/o ob
C0375367|T047|PT|574.61|ICD9CM|Calculus of gallbladder and bile duct with acute cholecystitis, with obstruction|Calculus of gallbladder and bile duct with acute cholecystitis, with obstruction
C0375367|T047|AB|574.61|ICD9CM|Gall&bil cal w/ac w obs|Gall&bil cal w/ac w obs
C0375368|T047|HT|574.7|ICD9CM|Calculus of gallbladder and bile duct with other cholecystitis|Calculus of gallbladder and bile duct with other cholecystitis
C0375369|T047|PT|574.70|ICD9CM|Calculus of gallbladder and bile duct with other cholecystitis, without mention of obstruction|Calculus of gallbladder and bile duct with other cholecystitis, without mention of obstruction
C0375369|T047|AB|574.70|ICD9CM|Gal&bil cal w/oth w/o ob|Gal&bil cal w/oth w/o ob
C0375370|T047|PT|574.71|ICD9CM|Calculus of gallbladder and bile duct with other cholecystitis, with obstruction|Calculus of gallbladder and bile duct with other cholecystitis, with obstruction
C0375370|T047|AB|574.71|ICD9CM|Gall&bil cal w/oth w obs|Gall&bil cal w/oth w obs
C0375371|T047|HT|574.8|ICD9CM|Calculus of gallbladder and bile duct with acute and chronic cholecystitis|Calculus of gallbladder and bile duct with acute and chronic cholecystitis
C0375372|T047|AB|574.80|ICD9CM|Gal&bil cal w/ac&chr w/o|Gal&bil cal w/ac&chr w/o
C0375373|T047|PT|574.81|ICD9CM|Calculus of gallbladder and bile duct with acute and chronic cholecystitis, with obstruction|Calculus of gallbladder and bile duct with acute and chronic cholecystitis, with obstruction
C0375373|T047|AB|574.81|ICD9CM|Gal&bil cal w/ac&ch w ob|Gal&bil cal w/ac&ch w ob
C0375374|T047|HT|574.9|ICD9CM|Calculus of gallbladder and bile duct without cholecystitis|Calculus of gallbladder and bile duct without cholecystitis
C0375375|T047|PT|574.90|ICD9CM|Calculus of gallbladder and bile duct without cholecystitis, without mention of obstruction|Calculus of gallbladder and bile duct without cholecystitis, without mention of obstruction
C0375375|T047|AB|574.90|ICD9CM|Gall&bil cal w/o cho w/o|Gall&bil cal w/o cho w/o
C0375376|T047|PT|574.91|ICD9CM|Calculus of gallbladder and bile duct without cholecystitis, with obstruction|Calculus of gallbladder and bile duct without cholecystitis, with obstruction
C0375376|T047|AB|574.91|ICD9CM|Gall&bil cal w/o ch w ob|Gall&bil cal w/o ch w ob
C0156213|T047|HT|575|ICD9CM|Other disorders of gallbladder|Other disorders of gallbladder
C0149520|T047|AB|575.0|ICD9CM|Acute cholecystitis|Acute cholecystitis
C0149520|T047|PT|575.0|ICD9CM|Acute cholecystitis|Acute cholecystitis
C0029539|T047|HT|575.1|ICD9CM|Other cholecystitis|Other cholecystitis
C0008325|T047|AB|575.10|ICD9CM|Cholecystitis NOS|Cholecystitis NOS
C0008325|T047|PT|575.10|ICD9CM|Cholecystitis, unspecified|Cholecystitis, unspecified
C0085694|T047|AB|575.11|ICD9CM|Chronic cholecystitis|Chronic cholecystitis
C0085694|T047|PT|575.11|ICD9CM|Chronic cholecystitis|Chronic cholecystitis
C0302472|T047|AB|575.12|ICD9CM|Acte & chr cholecystitis|Acte & chr cholecystitis
C0302472|T047|PT|575.12|ICD9CM|Acute and chronic cholecystitis|Acute and chronic cholecystitis
C0156214|T047|AB|575.2|ICD9CM|Obstruction gallbladder|Obstruction gallbladder
C0156214|T047|PT|575.2|ICD9CM|Obstruction of gallbladder|Obstruction of gallbladder
C0152445|T047|AB|575.3|ICD9CM|Hydrops of gallbladder|Hydrops of gallbladder
C0152445|T047|PT|575.3|ICD9CM|Hydrops of gallbladder|Hydrops of gallbladder
C0156215|T037|AB|575.4|ICD9CM|Perforation gallbladder|Perforation gallbladder
C0156215|T037|PT|575.4|ICD9CM|Perforation of gallbladder|Perforation of gallbladder
C0156216|T190|AB|575.5|ICD9CM|Fistula of gallbladder|Fistula of gallbladder
C0156216|T190|PT|575.5|ICD9CM|Fistula of gallbladder|Fistula of gallbladder
C0152456|T047|PT|575.6|ICD9CM|Cholesterolosis of gallbladder|Cholesterolosis of gallbladder
C0152456|T047|AB|575.6|ICD9CM|Gb cholesterolosis|Gb cholesterolosis
C0348758|T047|AB|575.8|ICD9CM|Dis of gallbladder NEC|Dis of gallbladder NEC
C0348758|T047|PT|575.8|ICD9CM|Other specified disorders of gallbladder|Other specified disorders of gallbladder
C0016977|T047|AB|575.9|ICD9CM|Dis of gallbladder NOS|Dis of gallbladder NOS
C0016977|T047|PT|575.9|ICD9CM|Unspecified disorder of gallbladder|Unspecified disorder of gallbladder
C0156217|T047|HT|576|ICD9CM|Other disorders of biliary tract|Other disorders of biliary tract
C0152099|T047|AB|576.0|ICD9CM|Postcholecystectomy synd|Postcholecystectomy synd
C0152099|T047|PT|576.0|ICD9CM|Postcholecystectomy syndrome|Postcholecystectomy syndrome
C0008311|T047|AB|576.1|ICD9CM|Cholangitis|Cholangitis
C0008311|T047|PT|576.1|ICD9CM|Cholangitis|Cholangitis
C0008370|T047|AB|576.2|ICD9CM|Obstruction of bile duct|Obstruction of bile duct
C0008370|T047|PT|576.2|ICD9CM|Obstruction of bile duct|Obstruction of bile duct
C0156218|T047|AB|576.3|ICD9CM|Perforation of bile duct|Perforation of bile duct
C0156218|T047|PT|576.3|ICD9CM|Perforation of bile duct|Perforation of bile duct
C0005417|T046|AB|576.4|ICD9CM|Fistula of bile duct|Fistula of bile duct
C0005417|T046|PT|576.4|ICD9CM|Fistula of bile duct|Fistula of bile duct
C0152168|T046|PT|576.5|ICD9CM|Spasm of sphincter of Oddi|Spasm of sphincter of Oddi
C0152168|T046|AB|576.5|ICD9CM|Spasm sphincter of oddi|Spasm sphincter of oddi
C0348759|T047|AB|576.8|ICD9CM|Dis of biliary tract NEC|Dis of biliary tract NEC
C0348759|T047|PT|576.8|ICD9CM|Other specified disorders of biliary tract|Other specified disorders of biliary tract
C0005424|T047|AB|576.9|ICD9CM|Dis of biliary tract NOS|Dis of biliary tract NOS
C0005424|T047|PT|576.9|ICD9CM|Unspecified disorder of biliary tract|Unspecified disorder of biliary tract
C0030286|T047|HT|577|ICD9CM|Diseases of pancreas|Diseases of pancreas
C0001339|T047|AB|577.0|ICD9CM|Acute pancreatitis|Acute pancreatitis
C0001339|T047|PT|577.0|ICD9CM|Acute pancreatitis|Acute pancreatitis
C0149521|T047|AB|577.1|ICD9CM|Chronic pancreatitis|Chronic pancreatitis
C0149521|T047|PT|577.1|ICD9CM|Chronic pancreatitis|Chronic pancreatitis
C0010623|T190|PT|577.2|ICD9CM|Cyst and pseudocyst of pancreas|Cyst and pseudocyst of pancreas
C0010623|T190|AB|577.2|ICD9CM|Pancreat cyst/pseudocyst|Pancreat cyst/pseudocyst
C0029771|T047|PT|577.8|ICD9CM|Other specified diseases of pancreas|Other specified diseases of pancreas
C0029771|T047|AB|577.8|ICD9CM|Pancreatic disease NEC|Pancreatic disease NEC
C0030286|T047|AB|577.9|ICD9CM|Pancreatic disease NOS|Pancreatic disease NOS
C0030286|T047|PT|577.9|ICD9CM|Unspecified disease of pancreas|Unspecified disease of pancreas
C0017181|T046|HT|578|ICD9CM|Gastrointestinal hemorrhage|Gastrointestinal hemorrhage
C0018926|T184|AB|578.0|ICD9CM|Hematemesis|Hematemesis
C0018926|T184|PT|578.0|ICD9CM|Hematemesis|Hematemesis
C1321898|T184|AB|578.1|ICD9CM|Blood in stool|Blood in stool
C1321898|T184|PT|578.1|ICD9CM|Blood in stool|Blood in stool
C0017181|T046|AB|578.9|ICD9CM|Gastrointest hemorr NOS|Gastrointest hemorr NOS
C0017181|T046|PT|578.9|ICD9CM|Hemorrhage of gastrointestinal tract, unspecified|Hemorrhage of gastrointestinal tract, unspecified
C0024523|T047|HT|579|ICD9CM|Intestinal malabsorption|Intestinal malabsorption
C0007570|T047|AB|579.0|ICD9CM|Celiac disease|Celiac disease
C0007570|T047|PT|579.0|ICD9CM|Celiac disease|Celiac disease
C0038054|T047|AB|579.1|ICD9CM|Tropical sprue|Tropical sprue
C0038054|T047|PT|579.1|ICD9CM|Tropical sprue|Tropical sprue
C0005750|T047|AB|579.2|ICD9CM|Blind loop syndrome|Blind loop syndrome
C0005750|T047|PT|579.2|ICD9CM|Blind loop syndrome|Blind loop syndrome
C0029515|T033|AB|579.3|ICD9CM|Intest postop nonabsorb|Intest postop nonabsorb
C0029515|T033|PT|579.3|ICD9CM|Other and unspecified postsurgical nonabsorption|Other and unspecified postsurgical nonabsorption
C0152166|T047|AB|579.4|ICD9CM|Pancreatic steatorrhea|Pancreatic steatorrhea
C0152166|T047|PT|579.4|ICD9CM|Pancreatic steatorrhea|Pancreatic steatorrhea
C0029809|T047|AB|579.8|ICD9CM|Intest malabsorption NEC|Intest malabsorption NEC
C0029809|T047|PT|579.8|ICD9CM|Other specified intestinal malabsorption|Other specified intestinal malabsorption
C0024523|T047|AB|579.9|ICD9CM|Intest malabsorption NOS|Intest malabsorption NOS
C0024523|T047|PT|579.9|ICD9CM|Unspecified intestinal malabsorption|Unspecified intestinal malabsorption
C0156221|T047|HT|580|ICD9CM|Acute glomerulonephritis|Acute glomerulonephritis
C0178287|T047|HT|580-589.99|ICD9CM|NEPHRITIS, NEPHROTIC SYNDROME, AND NEPHROSIS|NEPHRITIS, NEPHROTIC SYNDROME, AND NEPHROSIS
C0080276|T047|HT|580-629.99|ICD9CM|DISEASES OF THE GENITOURINARY SYSTEM|DISEASES OF THE GENITOURINARY SYSTEM
C0341692|T047|AB|580.0|ICD9CM|Ac proliferat nephritis|Ac proliferat nephritis
C0341692|T047|PT|580.0|ICD9CM|Acute glomerulonephritis with lesion of proliferative glomerulonephritis|Acute glomerulonephritis with lesion of proliferative glomerulonephritis
C0156223|T047|AB|580.4|ICD9CM|Ac rapidly progr nephrit|Ac rapidly progr nephrit
C0156223|T047|PT|580.4|ICD9CM|Acute glomerulonephritis with lesion of rapidly progressive glomerulonephritis|Acute glomerulonephritis with lesion of rapidly progressive glomerulonephritis
C0156224|T047|HT|580.8|ICD9CM|Acute glomerulonephritis with other specified pathological lesion in kidney|Acute glomerulonephritis with other specified pathological lesion in kidney
C0156225|T047|AB|580.81|ICD9CM|Ac nephritis in oth dis|Ac nephritis in oth dis
C0156225|T047|PT|580.81|ICD9CM|Acute glomerulonephritis in diseases classified elsewhere|Acute glomerulonephritis in diseases classified elsewhere
C0156224|T047|PT|580.89|ICD9CM|Acute glomerulonephritis with other specified pathological lesion in kidney|Acute glomerulonephritis with other specified pathological lesion in kidney
C0156224|T047|AB|580.89|ICD9CM|Acute nephritis NEC|Acute nephritis NEC
C0156226|T047|PT|580.9|ICD9CM|Acute glomerulonephritis with unspecified pathological lesion in kidney|Acute glomerulonephritis with unspecified pathological lesion in kidney
C0156226|T047|AB|580.9|ICD9CM|Acute nephritis NOS|Acute nephritis NOS
C0027726|T047|HT|581|ICD9CM|Nephrotic syndrome|Nephrotic syndrome
C0156227|T047|AB|581.0|ICD9CM|Nephrotic syn, prolifer|Nephrotic syn, prolifer
C0156227|T047|PT|581.0|ICD9CM|Nephrotic syndrome with lesion of proliferative glomerulonephritis|Nephrotic syndrome with lesion of proliferative glomerulonephritis
C0156228|T047|AB|581.1|ICD9CM|Epimembranous nephritis|Epimembranous nephritis
C0156228|T047|PT|581.1|ICD9CM|Nephrotic syndrome with lesion of membranous glomerulonephritis|Nephrotic syndrome with lesion of membranous glomerulonephritis
C0156229|T047|AB|581.2|ICD9CM|Membranoprolif nephrosis|Membranoprolif nephrosis
C0156229|T047|PT|581.2|ICD9CM|Nephrotic syndrome with lesion of membranoproliferative glomerulonephritis|Nephrotic syndrome with lesion of membranoproliferative glomerulonephritis
C1704321|T047|AB|581.3|ICD9CM|Minimal change nephrosis|Minimal change nephrosis
C1704321|T047|PT|581.3|ICD9CM|Nephrotic syndrome with lesion of minimal change glomerulonephritis|Nephrotic syndrome with lesion of minimal change glomerulonephritis
C0027729|T047|HT|581.8|ICD9CM|Nephrotic syndrome with other specified pathological lesion in kidney|Nephrotic syndrome with other specified pathological lesion in kidney
C0156230|T047|AB|581.81|ICD9CM|Nephrotic syn in oth dis|Nephrotic syn in oth dis
C0156230|T047|PT|581.81|ICD9CM|Nephrotic syndrome in diseases classified elsewhere|Nephrotic syndrome in diseases classified elsewhere
C0027729|T047|AB|581.89|ICD9CM|Nephrotic syndrome NEC|Nephrotic syndrome NEC
C0027729|T047|PT|581.89|ICD9CM|Nephrotic syndrome with other specified pathological lesion in kidney|Nephrotic syndrome with other specified pathological lesion in kidney
C0027730|T047|AB|581.9|ICD9CM|Nephrotic syndrome NOS|Nephrotic syndrome NOS
C0027730|T047|PT|581.9|ICD9CM|Nephrotic syndrome with unspecified pathological lesion in kidney|Nephrotic syndrome with unspecified pathological lesion in kidney
C0152451|T047|HT|582|ICD9CM|Chronic glomerulonephritis|Chronic glomerulonephritis
C0156231|T047|AB|582.0|ICD9CM|Chr proliferat nephritis|Chr proliferat nephritis
C0156231|T047|PT|582.0|ICD9CM|Chronic glomerulonephritis with lesion of proliferative glomerulonephritis|Chronic glomerulonephritis with lesion of proliferative glomerulonephritis
C0008686|T047|AB|582.1|ICD9CM|Chr membranous nephritis|Chr membranous nephritis
C0008686|T047|PT|582.1|ICD9CM|Chronic glomerulonephritis with lesion of membranous glomerulonephritis|Chronic glomerulonephritis with lesion of membranous glomerulonephritis
C0008685|T047|AB|582.2|ICD9CM|Chr membranoprolif nephr|Chr membranoprolif nephr
C0008685|T047|PT|582.2|ICD9CM|Chronic glomerulonephritis with lesion of membranoproliferative glomerulonephritis|Chronic glomerulonephritis with lesion of membranoproliferative glomerulonephritis
C0341694|T047|AB|582.4|ICD9CM|Chr rapid progr nephrit|Chr rapid progr nephrit
C0341694|T047|PT|582.4|ICD9CM|Chronic glomerulonephritis with lesion of rapidly progressive glomerulonephritis|Chronic glomerulonephritis with lesion of rapidly progressive glomerulonephritis
C0156233|T047|HT|582.8|ICD9CM|Chronic glomerulonephritis with other specified pathological lesion in kidney|Chronic glomerulonephritis with other specified pathological lesion in kidney
C0156234|T047|AB|582.81|ICD9CM|Chr nephritis in oth dis|Chr nephritis in oth dis
C0156234|T047|PT|582.81|ICD9CM|Chronic glomerulonephritis in diseases classified elsewhere|Chronic glomerulonephritis in diseases classified elsewhere
C0156233|T047|PT|582.89|ICD9CM|Chronic glomerulonephritis with other specified pathological lesion in kidney|Chronic glomerulonephritis with other specified pathological lesion in kidney
C0156233|T047|AB|582.89|ICD9CM|Chronic nephritis NEC|Chronic nephritis NEC
C0156235|T047|PT|582.9|ICD9CM|Chronic glomerulonephritis with unspecified pathological lesion in kidney|Chronic glomerulonephritis with unspecified pathological lesion in kidney
C0156235|T047|AB|582.9|ICD9CM|Chronic nephritis NOS|Chronic nephritis NOS
C0027698|T047|HT|583|ICD9CM|Nephritis and nephropathy, not specified as acute or chronic|Nephritis and nephropathy, not specified as acute or chronic
C0156236|T047|AB|583.0|ICD9CM|Proliferat nephritis NOS|Proliferat nephritis NOS
C0027701|T047|AB|583.1|ICD9CM|Membranous nephritis NOS|Membranous nephritis NOS
C0027700|T047|AB|583.2|ICD9CM|Membranoprolif nephr NOS|Membranoprolif nephr NOS
C0156237|T047|AB|583.4|ICD9CM|Rapidly prog nephrit NOS|Rapidly prog nephrit NOS
C0156238|T047|PT|583.6|ICD9CM|Nephritis and nephropathy, not specified as acute or chronic, with lesion of renal cortical necrosis|Nephritis and nephropathy, not specified as acute or chronic, with lesion of renal cortical necrosis
C0156238|T047|AB|583.6|ICD9CM|Renal cort necrosis NOS|Renal cort necrosis NOS
C0156239|T047|AB|583.7|ICD9CM|Nephr NOS/medull necros|Nephr NOS/medull necros
C0027699|T047|PT|583.81|ICD9CM|Nephritis and nephropathy, not specified as acute or chronic, in diseases classified elsewhere|Nephritis and nephropathy, not specified as acute or chronic, in diseases classified elsewhere
C0027699|T047|AB|583.81|ICD9CM|Nephritis NOS in oth dis|Nephritis NOS in oth dis
C0027702|T047|AB|583.89|ICD9CM|Nephritis NEC|Nephritis NEC
C0027703|T047|AB|583.9|ICD9CM|Nephritis NOS|Nephritis NOS
C0022660|T047|HT|584|ICD9CM|Acute kidney failure|Acute kidney failure
C2712977|T047|AB|584.5|ICD9CM|Ac kidny fail, tubr necr|Ac kidny fail, tubr necr
C2712977|T047|PT|584.5|ICD9CM|Acute kidney failure with lesion of tubular necrosis|Acute kidney failure with lesion of tubular necrosis
C2712983|T047|AB|584.6|ICD9CM|Ac kidny fail, cort necr|Ac kidny fail, cort necr
C2712983|T047|PT|584.6|ICD9CM|Acute kidney failure with lesion of renal cortical necrosis|Acute kidney failure with lesion of renal cortical necrosis
C2712745|T047|AB|584.7|ICD9CM|Ac kidny fail, medu necr|Ac kidny fail, medu necr
C2712745|T047|PT|584.7|ICD9CM|Acute kidney failure with lesion of renal medullary [papillary] necrosis|Acute kidney failure with lesion of renal medullary [papillary] necrosis
C2712988|T047|AB|584.8|ICD9CM|Acute kidney failure NEC|Acute kidney failure NEC
C2712988|T047|PT|584.8|ICD9CM|Acute kidney failure with other specified pathological lesion in kidney|Acute kidney failure with other specified pathological lesion in kidney
C0022660|T047|AB|584.9|ICD9CM|Acute kidney failure NOS|Acute kidney failure NOS
C0022660|T047|PT|584.9|ICD9CM|Acute kidney failure, unspecified|Acute kidney failure, unspecified
C1561643|T047|HT|585|ICD9CM|Chronic kidney disease (CKD)|Chronic kidney disease (CKD)
C1561638|T047|AB|585.1|ICD9CM|Chro kidney dis stage I|Chro kidney dis stage I
C1561638|T047|PT|585.1|ICD9CM|Chronic kidney disease, Stage I|Chronic kidney disease, Stage I
C1561639|T047|AB|585.2|ICD9CM|Chro kidney dis stage II|Chro kidney dis stage II
C1561639|T047|PT|585.2|ICD9CM|Chronic kidney disease, Stage II (mild)|Chronic kidney disease, Stage II (mild)
C1561640|T047|AB|585.3|ICD9CM|Chr kidney dis stage III|Chr kidney dis stage III
C1561640|T047|PT|585.3|ICD9CM|Chronic kidney disease, Stage III (moderate)|Chronic kidney disease, Stage III (moderate)
C1561641|T047|AB|585.4|ICD9CM|Chr kidney dis stage IV|Chr kidney dis stage IV
C1561641|T047|PT|585.4|ICD9CM|Chronic kidney disease, Stage IV (severe)|Chronic kidney disease, Stage IV (severe)
C1561642|T047|AB|585.5|ICD9CM|Chron kidney dis stage V|Chron kidney dis stage V
C1561642|T047|PT|585.5|ICD9CM|Chronic kidney disease, Stage V|Chronic kidney disease, Stage V
C0022661|T047|AB|585.6|ICD9CM|End stage renal disease|End stage renal disease
C0022661|T047|PT|585.6|ICD9CM|End stage renal disease|End stage renal disease
C1561643|T047|AB|585.9|ICD9CM|Chronic kidney dis NOS|Chronic kidney dis NOS
C1561643|T047|PT|585.9|ICD9CM|Chronic kidney disease, unspecified|Chronic kidney disease, unspecified
C0035078|T047|AB|586|ICD9CM|Renal failure NOS|Renal failure NOS
C0035078|T047|PT|586|ICD9CM|Renal failure, unspecified|Renal failure, unspecified
C0027719|T047|AB|587|ICD9CM|Renal sclerosis NOS|Renal sclerosis NOS
C0027719|T047|PT|587|ICD9CM|Renal sclerosis, unspecified|Renal sclerosis, unspecified
C0341677|T047|HT|588|ICD9CM|Disorders resulting from impaired renal function|Disorders resulting from impaired renal function
C0035086|T047|AB|588.0|ICD9CM|Renal osteodystrophy|Renal osteodystrophy
C0035086|T047|PT|588.0|ICD9CM|Renal osteodystrophy|Renal osteodystrophy
C0162283|T047|AB|588.1|ICD9CM|Nephrogen diabetes insip|Nephrogen diabetes insip
C0162283|T047|PT|588.1|ICD9CM|Nephrogenic diabetes insipidus|Nephrogenic diabetes insipidus
C0029791|T047|HT|588.8|ICD9CM|Other specified disorders resulting from impaired renal function|Other specified disorders resulting from impaired renal function
C0271847|T047|AB|588.81|ICD9CM|Sec hyperparathyrd-renal|Sec hyperparathyrd-renal
C0271847|T047|PT|588.81|ICD9CM|Secondary hyperparathyroidism (of renal origin)|Secondary hyperparathyroidism (of renal origin)
C0029791|T047|AB|588.89|ICD9CM|Impair ren funct dis NEC|Impair ren funct dis NEC
C0029791|T047|PT|588.89|ICD9CM|Other specified disorders resulting from impaired renal function|Other specified disorders resulting from impaired renal function
C0341677|T047|AB|588.9|ICD9CM|Impaired renal funct NOS|Impaired renal funct NOS
C0341677|T047|PT|588.9|ICD9CM|Unspecified disorder resulting from impaired renal function|Unspecified disorder resulting from impaired renal function
C0156247|T033|HT|589|ICD9CM|Small kidney of unknown cause|Small kidney of unknown cause
C0156245|T019|AB|589.0|ICD9CM|Unilateral small kidney|Unilateral small kidney
C0156245|T019|PT|589.0|ICD9CM|Unilateral small kidney|Unilateral small kidney
C0156246|T190|AB|589.1|ICD9CM|Bilateral small kidneys|Bilateral small kidneys
C0156246|T190|PT|589.1|ICD9CM|Bilateral small kidneys|Bilateral small kidneys
C0156247|T033|AB|589.9|ICD9CM|Small kidney NOS|Small kidney NOS
C0156247|T033|PT|589.9|ICD9CM|Small kidney, unspecified|Small kidney, unspecified
C0021313|T047|HT|590|ICD9CM|Infections of kidney|Infections of kidney
C0178288|T047|HT|590-599.99|ICD9CM|OTHER DISEASES OF URINARY SYSTEM|OTHER DISEASES OF URINARY SYSTEM
C0085697|T047|HT|590.0|ICD9CM|Chronic pyelonephritis|Chronic pyelonephritis
C0156249|T047|AB|590.00|ICD9CM|Chr pyelonephritis NOS|Chr pyelonephritis NOS
C0156249|T047|PT|590.00|ICD9CM|Chronic pyelonephritis without lesion of renal medullary necrosis|Chronic pyelonephritis without lesion of renal medullary necrosis
C0156250|T047|AB|590.01|ICD9CM|Chr pyeloneph w med necr|Chr pyeloneph w med necr
C0156250|T047|PT|590.01|ICD9CM|Chronic pyelonephritis with lesion of renal medullary necrosis|Chronic pyelonephritis with lesion of renal medullary necrosis
C0520575|T047|HT|590.1|ICD9CM|Acute pyelonephritis|Acute pyelonephritis
C0156251|T047|AB|590.10|ICD9CM|Ac pyelonephritis NOS|Ac pyelonephritis NOS
C0156251|T047|PT|590.10|ICD9CM|Acute pyelonephritis without lesion of renal medullary necrosis|Acute pyelonephritis without lesion of renal medullary necrosis
C0156252|T047|AB|590.11|ICD9CM|Ac pyelonephr w med necr|Ac pyelonephr w med necr
C0156252|T047|PT|590.11|ICD9CM|Acute pyelonephritis with lesion of renal medullary necrosis|Acute pyelonephritis with lesion of renal medullary necrosis
C0156253|T047|PT|590.2|ICD9CM|Renal and perinephric abscess|Renal and perinephric abscess
C0156253|T047|AB|590.2|ICD9CM|Renal/perirenal abscess|Renal/perirenal abscess
C0156254|T047|AB|590.3|ICD9CM|Pyeloureteritis cystica|Pyeloureteritis cystica
C0156254|T047|PT|590.3|ICD9CM|Pyeloureteritis cystica|Pyeloureteritis cystica
C0156255|T047|HT|590.8|ICD9CM|Other pyelonephritis or pyonephrosis, not specified as acute or chronic|Other pyelonephritis or pyonephrosis, not specified as acute or chronic
C0034186|T047|AB|590.80|ICD9CM|Pyelonephritis NOS|Pyelonephritis NOS
C0034186|T047|PT|590.80|ICD9CM|Pyelonephritis, unspecified|Pyelonephritis, unspecified
C0156256|T047|PT|590.81|ICD9CM|Pyelitis or pyelonephritis in diseases classified elsewhere|Pyelitis or pyelonephritis in diseases classified elsewhere
C0156256|T047|AB|590.81|ICD9CM|Pyelonephrit in oth dis|Pyelonephrit in oth dis
C0021313|T047|AB|590.9|ICD9CM|Infection of kidney NOS|Infection of kidney NOS
C0021313|T047|PT|590.9|ICD9CM|Infection of kidney, unspecified|Infection of kidney, unspecified
C0020295|T047|AB|591|ICD9CM|Hydronephrosis|Hydronephrosis
C0020295|T047|PT|591|ICD9CM|Hydronephrosis|Hydronephrosis
C0156257|T047|HT|592|ICD9CM|Calculus of kidney and ureter|Calculus of kidney and ureter
C0022650|T047|AB|592.0|ICD9CM|Calculus of kidney|Calculus of kidney
C0022650|T047|PT|592.0|ICD9CM|Calculus of kidney|Calculus of kidney
C0041952|T047|AB|592.1|ICD9CM|Calculus of ureter|Calculus of ureter
C0041952|T047|PT|592.1|ICD9CM|Calculus of ureter|Calculus of ureter
C4759702|T047|AB|592.9|ICD9CM|Urinary calculus NOS|Urinary calculus NOS
C4759702|T047|PT|592.9|ICD9CM|Urinary calculus, unspecified|Urinary calculus, unspecified
C0156258|T047|HT|593|ICD9CM|Other disorders of kidney and ureter|Other disorders of kidney and ureter
C1384594|T047|AB|593.0|ICD9CM|Nephroptosis|Nephroptosis
C1384594|T047|PT|593.0|ICD9CM|Nephroptosis|Nephroptosis
C0156259|T047|AB|593.1|ICD9CM|Hypertrophy of kidney|Hypertrophy of kidney
C0156259|T047|PT|593.1|ICD9CM|Hypertrophy of kidney|Hypertrophy of kidney
C0268799|T047|AB|593.2|ICD9CM|Cyst of kidney, acquired|Cyst of kidney, acquired
C0268799|T047|PT|593.2|ICD9CM|Cyst of kidney, acquired|Cyst of kidney, acquired
C0156261|T020|AB|593.3|ICD9CM|Stricture of ureter|Stricture of ureter
C0156261|T020|PT|593.3|ICD9CM|Stricture or kinking of ureter|Stricture or kinking of ureter
C0029866|T190|PT|593.4|ICD9CM|Other ureteric obstruction|Other ureteric obstruction
C0029866|T190|AB|593.4|ICD9CM|Ureteric obstruction NEC|Ureteric obstruction NEC
C0521620|T190|AB|593.5|ICD9CM|Hydroureter|Hydroureter
C0521620|T190|PT|593.5|ICD9CM|Hydroureter|Hydroureter
C0232867|T047|AB|593.6|ICD9CM|Postural proteinuria|Postural proteinuria
C0232867|T047|PT|593.6|ICD9CM|Postural proteinuria|Postural proteinuria
C0042580|T047|HT|593.7|ICD9CM|Vesicoureteral reflux|Vesicoureteral reflux
C0490048|T047|AB|593.70|ICD9CM|Vescouretrl rflux unspcf|Vescouretrl rflux unspcf
C0490048|T047|PT|593.70|ICD9CM|Vesicoureteral reflux unspecified or without reflux nephropathy|Vesicoureteral reflux unspecified or without reflux nephropathy
C0375377|T047|PT|593.71|ICD9CM|Vesicoureteral reflux with reflux nephropathy, unilateral|Vesicoureteral reflux with reflux nephropathy, unilateral
C0375377|T047|AB|593.71|ICD9CM|Vscurt rflx npht uniltrl|Vscurt rflx npht uniltrl
C0375378|T047|PT|593.72|ICD9CM|Vesicoureteral reflux with reflux nephropathy, bilateral|Vesicoureteral reflux with reflux nephropathy, bilateral
C0375378|T047|AB|593.72|ICD9CM|Vscourtl rflx npht bltrl|Vscourtl rflx npht bltrl
C0375379|T047|PT|593.73|ICD9CM|Other vesicoureteral reflux with reflux nephropathy NOS|Other vesicoureteral reflux with reflux nephropathy NOS
C0375379|T047|AB|593.73|ICD9CM|Vscourtl rflx w npht NOS|Vscourtl rflx w npht NOS
C0029781|T047|HT|593.8|ICD9CM|Other specified disorders of kidney and ureter|Other specified disorders of kidney and ureter
C0268790|T047|AB|593.81|ICD9CM|Renal vascular disorder|Renal vascular disorder
C0268790|T047|PT|593.81|ICD9CM|Vascular disorders of kidney|Vascular disorders of kidney
C0156263|T020|AB|593.82|ICD9CM|Ureteral fistula|Ureteral fistula
C0156263|T020|PT|593.82|ICD9CM|Ureteral fistula|Ureteral fistula
C0029781|T047|PT|593.89|ICD9CM|Other specified disorders of kidney and ureter|Other specified disorders of kidney and ureter
C0029781|T047|AB|593.89|ICD9CM|Renal & ureteral dis NEC|Renal & ureteral dis NEC
C0268701|T047|AB|593.9|ICD9CM|Renal & ureteral dis NOS|Renal & ureteral dis NOS
C0268701|T047|PT|593.9|ICD9CM|Unspecified disorder of kidney and ureter|Unspecified disorder of kidney and ureter
C0156264|T047|HT|594|ICD9CM|Calculus of lower urinary tract|Calculus of lower urinary tract
C0156265|T047|AB|594.0|ICD9CM|Blad diverticulum calcul|Blad diverticulum calcul
C0156265|T047|PT|594.0|ICD9CM|Calculus in diverticulum of bladder|Calculus in diverticulum of bladder
C1961101|T047|AB|594.1|ICD9CM|Bladder calculus NEC|Bladder calculus NEC
C1961101|T047|PT|594.1|ICD9CM|Other calculus in bladder|Other calculus in bladder
C0162301|T047|PT|594.2|ICD9CM|Calculus in urethra|Calculus in urethra
C0162301|T047|AB|594.2|ICD9CM|Urethral calculus|Urethral calculus
C0156266|T047|AB|594.8|ICD9CM|Lower urin calcul NEC|Lower urin calcul NEC
C0156266|T047|PT|594.8|ICD9CM|Other lower urinary tract calculus|Other lower urinary tract calculus
C0156264|T047|PT|594.9|ICD9CM|Calculus of lower urinary tract, unspecified|Calculus of lower urinary tract, unspecified
C0156264|T047|AB|594.9|ICD9CM|Lower urin calcul NOS|Lower urin calcul NOS
C0010692|T047|HT|595|ICD9CM|Cystitis|Cystitis
C0149523|T047|AB|595.0|ICD9CM|Acute cystitis|Acute cystitis
C0149523|T047|PT|595.0|ICD9CM|Acute cystitis|Acute cystitis
C0600040|T047|AB|595.1|ICD9CM|Chr interstit cystitis|Chr interstit cystitis
C0600040|T047|PT|595.1|ICD9CM|Chronic interstitial cystitis|Chronic interstitial cystitis
C0156268|T047|AB|595.2|ICD9CM|Chronic cystitis NEC|Chronic cystitis NEC
C0156268|T047|PT|595.2|ICD9CM|Other chronic cystitis|Other chronic cystitis
C1261278|T047|AB|595.3|ICD9CM|Trigonitis|Trigonitis
C1261278|T047|PT|595.3|ICD9CM|Trigonitis|Trigonitis
C0156269|T047|PT|595.4|ICD9CM|Cystitis in diseases classified elsewhere|Cystitis in diseases classified elsewhere
C0156269|T047|AB|595.4|ICD9CM|Cystitis in oth dis|Cystitis in oth dis
C0029836|T047|HT|595.8|ICD9CM|Other specified types of cystitis|Other specified types of cystitis
C0152262|T047|AB|595.81|ICD9CM|Cystitis cystica|Cystitis cystica
C0152262|T047|PT|595.81|ICD9CM|Cystitis cystica|Cystitis cystica
C0156270|T047|AB|595.82|ICD9CM|Irradiation cystitis|Irradiation cystitis
C0156270|T047|PT|595.82|ICD9CM|Irradiation cystitis|Irradiation cystitis
C0029836|T047|AB|595.89|ICD9CM|Cystitis NEC|Cystitis NEC
C0029836|T047|PT|595.89|ICD9CM|Other specified types of cystitis|Other specified types of cystitis
C0010692|T047|AB|595.9|ICD9CM|Cystitis NOS|Cystitis NOS
C0010692|T047|PT|595.9|ICD9CM|Cystitis, unspecified|Cystitis, unspecified
C0156271|T047|HT|596|ICD9CM|Other disorders of bladder|Other disorders of bladder
C0005694|T047|AB|596.0|ICD9CM|Bladder neck obstruction|Bladder neck obstruction
C0005694|T047|PT|596.0|ICD9CM|Bladder neck obstruction|Bladder neck obstruction
C0156272|T047|AB|596.1|ICD9CM|Intestinovesical fistula|Intestinovesical fistula
C0156272|T047|PT|596.1|ICD9CM|Intestinovesical fistula|Intestinovesical fistula
C0868850|T190|AB|596.2|ICD9CM|Vesical fistula NEC|Vesical fistula NEC
C0868850|T190|PT|596.2|ICD9CM|Vesical fistula, not elsewhere classified|Vesical fistula, not elsewhere classified
C0156273|T020|AB|596.3|ICD9CM|Diverticulum of bladder|Diverticulum of bladder
C0156273|T020|PT|596.3|ICD9CM|Diverticulum of bladder|Diverticulum of bladder
C0403645|T033|AB|596.4|ICD9CM|Atony of bladder|Atony of bladder
C0403645|T033|PT|596.4|ICD9CM|Atony of bladder|Atony of bladder
C0156274|T046|HT|596.5|ICD9CM|Other functional disorders of bladder|Other functional disorders of bladder
C0878773|T047|AB|596.51|ICD9CM|Hypertonicity of bladder|Hypertonicity of bladder
C0878773|T047|PT|596.51|ICD9CM|Hypertonicity of bladder|Hypertonicity of bladder
C0489967|T047|AB|596.52|ICD9CM|Low bladder compliance|Low bladder compliance
C0489967|T047|PT|596.52|ICD9CM|Low bladder compliance|Low bladder compliance
C0235093|T033|AB|596.53|ICD9CM|Paralysis of bladder|Paralysis of bladder
C0235093|T033|PT|596.53|ICD9CM|Paralysis of bladder|Paralysis of bladder
C0005697|T047|AB|596.54|ICD9CM|Neurogenic bladder NOS|Neurogenic bladder NOS
C0005697|T047|PT|596.54|ICD9CM|Neurogenic bladder NOS|Neurogenic bladder NOS
C0341747|T047|PT|596.55|ICD9CM|Detrusor sphincter dyssynergia|Detrusor sphincter dyssynergia
C0341747|T047|AB|596.55|ICD9CM|Detrusr sphinc dyssnrgia|Detrusr sphinc dyssnrgia
C0156274|T046|AB|596.59|ICD9CM|Oth func dsdr bladder|Oth func dsdr bladder
C0156274|T046|PT|596.59|ICD9CM|Other functional disorder of bladder|Other functional disorder of bladder
C0156275|T047|AB|596.6|ICD9CM|Bladder rupt, nontraum|Bladder rupt, nontraum
C0156275|T047|PT|596.6|ICD9CM|Rupture of bladder, nontraumatic|Rupture of bladder, nontraumatic
C0156276|T046|AB|596.7|ICD9CM|Bladder wall hemorrhage|Bladder wall hemorrhage
C0156276|T046|PT|596.7|ICD9CM|Hemorrhage into bladder wall|Hemorrhage into bladder wall
C0029776|T047|HT|596.8|ICD9CM|Other specified disorders of bladder|Other specified disorders of bladder
C2903163|T046|AB|596.81|ICD9CM|Infection of cystostomy|Infection of cystostomy
C2903163|T046|PT|596.81|ICD9CM|Infection of cystostomy|Infection of cystostomy
C3161117|T046|AB|596.82|ICD9CM|Mech comp of cystostomy|Mech comp of cystostomy
C3161117|T046|PT|596.82|ICD9CM|Mechanical complication of cystostomy|Mechanical complication of cystostomy
C2903164|T046|AB|596.83|ICD9CM|Other comp of cystostomy|Other comp of cystostomy
C2903164|T046|PT|596.83|ICD9CM|Other complication of cystostomy|Other complication of cystostomy
C0029776|T047|AB|596.89|ICD9CM|Disorders of bladder NEC|Disorders of bladder NEC
C0029776|T047|PT|596.89|ICD9CM|Other specified disorders of bladder|Other specified disorders of bladder
C0005686|T047|AB|596.9|ICD9CM|Bladder disorder NOS|Bladder disorder NOS
C0005686|T047|PT|596.9|ICD9CM|Unspecified disorder of bladder|Unspecified disorder of bladder
C0156277|T047|HT|597|ICD9CM|Urethritis, not sexually transmitted, and urethral syndrome|Urethritis, not sexually transmitted, and urethral syndrome
C0156278|T047|AB|597.0|ICD9CM|Urethral abscess|Urethral abscess
C0156278|T047|PT|597.0|ICD9CM|Urethral abscess|Urethral abscess
C0029867|T047|HT|597.8|ICD9CM|Other urethritis|Other urethritis
C0311389|T047|AB|597.80|ICD9CM|Urethritis NOS|Urethritis NOS
C0311389|T047|PT|597.80|ICD9CM|Urethritis, unspecified|Urethritis, unspecified
C0156279|T047|AB|597.81|ICD9CM|Urethral syndrome NOS|Urethral syndrome NOS
C0156279|T047|PT|597.81|ICD9CM|Urethral syndrome NOS|Urethral syndrome NOS
C0029867|T047|PT|597.89|ICD9CM|Other urethritis|Other urethritis
C0029867|T047|AB|597.89|ICD9CM|Urethritis NEC|Urethritis NEC
C4551691|T047|HT|598|ICD9CM|Urethral stricture|Urethral stricture
C0403696|T020|HT|598.0|ICD9CM|Urethral stricture due to infection|Urethral stricture due to infection
C0403696|T020|AB|598.00|ICD9CM|Urethr strict:infect NOS|Urethr strict:infect NOS
C0403696|T020|PT|598.00|ICD9CM|Urethral stricture due to unspecified infection|Urethral stricture due to unspecified infection
C0156282|T020|AB|598.01|ICD9CM|Ureth strict:oth infect|Ureth strict:oth infect
C0156282|T020|PT|598.01|ICD9CM|Urethral stricture due to infective diseases classified elsewhere|Urethral stricture due to infective diseases classified elsewhere
C0403698|T037|AB|598.1|ICD9CM|Traum urethral stricture|Traum urethral stricture
C0403698|T037|PT|598.1|ICD9CM|Traumatic urethral stricture|Traumatic urethral stricture
C0156284|T020|AB|598.2|ICD9CM|Postop urethral strictur|Postop urethral strictur
C0156284|T020|PT|598.2|ICD9CM|Postoperative urethral stricture|Postoperative urethral stricture
C0029752|T047|PT|598.8|ICD9CM|Other specified causes of urethral stricture|Other specified causes of urethral stricture
C0029752|T047|AB|598.8|ICD9CM|Urethral stricture NEC|Urethral stricture NEC
C4551691|T047|AB|598.9|ICD9CM|Urethral stricture NOS|Urethral stricture NOS
C4551691|T047|PT|598.9|ICD9CM|Urethral stricture, unspecified|Urethral stricture, unspecified
C0546812|T047|HT|599|ICD9CM|Other disorders of urethra and urinary tract|Other disorders of urethra and urinary tract
C0042029|T047|AB|599.0|ICD9CM|Urin tract infection NOS|Urin tract infection NOS
C0042029|T047|PT|599.0|ICD9CM|Urinary tract infection, site not specified|Urinary tract infection, site not specified
C0041970|T190|AB|599.1|ICD9CM|Urethral fistula|Urethral fistula
C0041970|T190|PT|599.1|ICD9CM|Urethral fistula|Urethral fistula
C0152443|T047|AB|599.2|ICD9CM|Urethral diverticulum|Urethral diverticulum
C0152443|T047|PT|599.2|ICD9CM|Urethral diverticulum|Urethral diverticulum
C0152247|T020|AB|599.3|ICD9CM|Urethral caruncle|Urethral caruncle
C0152247|T020|PT|599.3|ICD9CM|Urethral caruncle|Urethral caruncle
C0156286|T020|AB|599.4|ICD9CM|Urethral false passage|Urethral false passage
C0156286|T020|PT|599.4|ICD9CM|Urethral false passage|Urethral false passage
C0156287|T047|AB|599.5|ICD9CM|Prolapse urethral mucosa|Prolapse urethral mucosa
C0156287|T047|PT|599.5|ICD9CM|Prolapsed urethral mucosa|Prolapsed urethral mucosa
C0178879|T047|HT|599.6|ICD9CM|Urinary obstruction|Urinary obstruction
C0178879|T047|AB|599.60|ICD9CM|Urinary obstruction NOS|Urinary obstruction NOS
C0178879|T047|PT|599.60|ICD9CM|Urinary obstruction, unspecified|Urinary obstruction, unspecified
C1561646|T047|AB|599.69|ICD9CM|Urinary obstruction NEC|Urinary obstruction NEC
C1561646|T047|PT|599.69|ICD9CM|Urinary obstruction, not elsewhere classified|Urinary obstruction, not elsewhere classified
C0018965|T047|HT|599.7|ICD9CM|Hematuria|Hematuria
C0018965|T047|AB|599.70|ICD9CM|Hematuria NOS|Hematuria NOS
C0018965|T047|PT|599.70|ICD9CM|Hematuria, unspecified|Hematuria, unspecified
C0473237|T033|PT|599.71|ICD9CM|Gross hematuria|Gross hematuria
C0473237|T033|AB|599.71|ICD9CM|Gross hematuria|Gross hematuria
C0239937|T033|PT|599.72|ICD9CM|Microscopic hematuria|Microscopic hematuria
C0239937|T033|AB|599.72|ICD9CM|Microscopic hematuria|Microscopic hematuria
C0156288|T047|HT|599.8|ICD9CM|Other specified disorders of urethra and urinary tract|Other specified disorders of urethra and urinary tract
C0375380|T046|AB|599.81|ICD9CM|Urethral hypermobility|Urethral hypermobility
C0375380|T046|PT|599.81|ICD9CM|Urethral hypermobility|Urethral hypermobility
C0375381|T047|AB|599.82|ICD9CM|Intrinsc sphnctr dficncy|Intrinsc sphnctr dficncy
C0375381|T047|PT|599.82|ICD9CM|Intrinsic (urethral) sphincter deficiency [ISD]|Intrinsic (urethral) sphincter deficiency [ISD]
C0344436|T046|AB|599.83|ICD9CM|Urethral instability|Urethral instability
C0344436|T046|PT|599.83|ICD9CM|Urethral instability|Urethral instability
C0348769|T047|AB|599.84|ICD9CM|Oth spcf dsdr urethra|Oth spcf dsdr urethra
C0348769|T047|PT|599.84|ICD9CM|Other specified disorders of urethra|Other specified disorders of urethra
C0477758|T047|AB|599.89|ICD9CM|Oth spcf dsdr urnry trct|Oth spcf dsdr urnry trct
C0477758|T047|PT|599.89|ICD9CM|Other specified disorders of urinary tract|Other specified disorders of urinary tract
C0042075|T047|PT|599.9|ICD9CM|Unspecified disorder of urethra and urinary tract|Unspecified disorder of urethra and urinary tract
C0042075|T047|AB|599.9|ICD9CM|Urinary tract dis NOS|Urinary tract dis NOS
C2937421|T047|HT|600|ICD9CM|Hyperplasia of prostate|Hyperplasia of prostate
C0017412|T047|HT|600-608.99|ICD9CM|DISEASES OF MALE GENITAL ORGANS|DISEASES OF MALE GENITAL ORGANS
C0005001|T046|HT|600.0|ICD9CM|Hypertrophy (benign) of prostate|Hypertrophy (benign) of prostate
C1719538|T047|AB|600.00|ICD9CM|BPH w/o urinary obs/LUTS|BPH w/o urinary obs/LUTS
C1260419|T047|AB|600.01|ICD9CM|BPH w urinary obs/LUTS|BPH w urinary obs/LUTS
C0748012|T047|HT|600.1|ICD9CM|Nodular prostate|Nodular prostate
C1260421|T047|AB|600.10|ICD9CM|Nod prostate w/o ur obst|Nod prostate w/o ur obst
C1260421|T047|PT|600.10|ICD9CM|Nodular prostate without urinary obstruction|Nodular prostate without urinary obstruction
C1260422|T047|AB|600.11|ICD9CM|Nod prostate w ur obst|Nod prostate w ur obst
C1260422|T047|PT|600.11|ICD9CM|Nodular prostate with urinary obstruction|Nodular prostate with urinary obstruction
C0878697|T047|HT|600.2|ICD9CM|Benign localized hyperplasia of prostate|Benign localized hyperplasia of prostate
C1719539|T047|AB|600.20|ICD9CM|BPH loc w/o ur obs/LUTS|BPH loc w/o ur obs/LUTS
C1260424|T047|AB|600.21|ICD9CM|BPH loc w urin obs/LUTS|BPH loc w urin obs/LUTS
C1443972|T047|AB|600.3|ICD9CM|Cyst of prostate|Cyst of prostate
C1443972|T047|PT|600.3|ICD9CM|Cyst of prostate|Cyst of prostate
C2937421|T047|HT|600.9|ICD9CM|Hyperplasia of prostate, unspecified|Hyperplasia of prostate, unspecified
C1719540|T047|AB|600.90|ICD9CM|BPH NOS w/o ur obs/LUTS|BPH NOS w/o ur obs/LUTS
C1260426|T047|AB|600.91|ICD9CM|BPH NOS w ur obs/LUTS|BPH NOS w ur obs/LUTS
C0033581|T047|HT|601|ICD9CM|Inflammatory diseases of prostate|Inflammatory diseases of prostate
C0149524|T047|AB|601.0|ICD9CM|Acute prostatitis|Acute prostatitis
C0149524|T047|PT|601.0|ICD9CM|Acute prostatitis|Acute prostatitis
C0085696|T047|AB|601.1|ICD9CM|Chronic prostatitis|Chronic prostatitis
C0085696|T047|PT|601.1|ICD9CM|Chronic prostatitis|Chronic prostatitis
C0156290|T047|AB|601.2|ICD9CM|Abscess of prostate|Abscess of prostate
C0156290|T047|PT|601.2|ICD9CM|Abscess of prostate|Abscess of prostate
C0156291|T047|AB|601.3|ICD9CM|Prostatocystitis|Prostatocystitis
C0156291|T047|PT|601.3|ICD9CM|Prostatocystitis|Prostatocystitis
C1621349|T047|PT|601.4|ICD9CM|Prostatitis in diseases classified elsewhere|Prostatitis in diseases classified elsewhere
C1621349|T047|AB|601.4|ICD9CM|Prostatitis in oth dis|Prostatitis in oth dis
C0268882|T047|PT|601.8|ICD9CM|Other specified inflammatory diseases of prostate|Other specified inflammatory diseases of prostate
C0268882|T047|AB|601.8|ICD9CM|Prostatic inflam dis NEC|Prostatic inflam dis NEC
C0033581|T047|AB|601.9|ICD9CM|Prostatitis NOS|Prostatitis NOS
C0033581|T047|PT|601.9|ICD9CM|Prostatitis, unspecified|Prostatitis, unspecified
C0156294|T047|HT|602|ICD9CM|Other disorders of prostate|Other disorders of prostate
C0149525|T047|AB|602.0|ICD9CM|Calculus of prostate|Calculus of prostate
C0149525|T047|PT|602.0|ICD9CM|Calculus of prostate|Calculus of prostate
C0156295|T046|PT|602.1|ICD9CM|Congestion or hemorrhage of prostate|Congestion or hemorrhage of prostate
C0156295|T046|AB|602.1|ICD9CM|Prostatic congest/hemorr|Prostatic congest/hemorr
C0156296|T047|AB|602.2|ICD9CM|Atrophy of prostate|Atrophy of prostate
C0156296|T047|PT|602.2|ICD9CM|Atrophy of prostate|Atrophy of prostate
C0949136|T047|AB|602.3|ICD9CM|Dysplasia of prostate|Dysplasia of prostate
C0949136|T047|PT|602.3|ICD9CM|Dysplasia of prostate|Dysplasia of prostate
C0156297|T047|PT|602.8|ICD9CM|Other specified disorders of prostate|Other specified disorders of prostate
C0156297|T047|AB|602.8|ICD9CM|Prostatic disorders NEC|Prostatic disorders NEC
C0033575|T047|AB|602.9|ICD9CM|Prostatic disorder NOS|Prostatic disorder NOS
C0033575|T047|PT|602.9|ICD9CM|Unspecified disorder of prostate|Unspecified disorder of prostate
C1720771|T019|HT|603|ICD9CM|Hydrocele|Hydrocele
C0156299|T046|AB|603.0|ICD9CM|Encysted hydrocele|Encysted hydrocele
C0156299|T046|PT|603.0|ICD9CM|Encysted hydrocele|Encysted hydrocele
C0156300|T047|AB|603.1|ICD9CM|Infected hydrocele|Infected hydrocele
C0156300|T047|PT|603.1|ICD9CM|Infected hydrocele|Infected hydrocele
C0029837|T047|AB|603.8|ICD9CM|Hydrocele NEC|Hydrocele NEC
C0029837|T047|PT|603.8|ICD9CM|Other specified types of hydrocele|Other specified types of hydrocele
C1720771|T019|AB|603.9|ICD9CM|Hydrocele NOS|Hydrocele NOS
C1720771|T019|PT|603.9|ICD9CM|Hydrocele, unspecified|Hydrocele, unspecified
C0149881|T047|HT|604|ICD9CM|Orchitis and epididymitis|Orchitis and epididymitis
C0156301|T047|AB|604.0|ICD9CM|Orchitis with abscess|Orchitis with abscess
C0156301|T047|PT|604.0|ICD9CM|Orchitis, epididymitis, and epididymo-orchitis, with abscess|Orchitis, epididymitis, and epididymo-orchitis, with abscess
C0156302|T047|HT|604.9|ICD9CM|Other orchitis, epididymitis, and epididymo-orchitis, without mention of abscess|Other orchitis, epididymitis, and epididymo-orchitis, without mention of abscess
C0149881|T047|PT|604.90|ICD9CM|Orchitis and epididymitis, unspecified|Orchitis and epididymitis, unspecified
C0149881|T047|AB|604.90|ICD9CM|Orchitis/epididymit NOS|Orchitis/epididymit NOS
C0156303|T047|PT|604.91|ICD9CM|Orchitis and epididymitis in diseases classified elsewhere|Orchitis and epididymitis in diseases classified elsewhere
C0156303|T047|AB|604.91|ICD9CM|Orchitis in oth disease|Orchitis in oth disease
C0156302|T047|AB|604.99|ICD9CM|Orchitis/epididymit NEC|Orchitis/epididymit NEC
C0156302|T047|PT|604.99|ICD9CM|Other orchitis, epididymitis, and epididymo-orchitis, without mention of abscess|Other orchitis, epididymitis, and epididymo-orchitis, without mention of abscess
C0034919|T047|AB|605|ICD9CM|Redun prepuce & phimosis|Redun prepuce & phimosis
C0034919|T047|PT|605|ICD9CM|Redundant prepuce and phimosis|Redundant prepuce and phimosis
C0021364|T047|HT|606|ICD9CM|Infertility, male|Infertility, male
C0004509|T047|AB|606.0|ICD9CM|Azoospermia|Azoospermia
C0004509|T047|PT|606.0|ICD9CM|Azoospermia|Azoospermia
C0028960|T047|AB|606.1|ICD9CM|Oligospermia|Oligospermia
C0028960|T047|PT|606.1|ICD9CM|Oligospermia|Oligospermia
C0021360|T047|PT|606.8|ICD9CM|Infertility due to extratesticular causes|Infertility due to extratesticular causes
C0021360|T047|AB|606.8|ICD9CM|Male infertility NEC|Male infertility NEC
C0021364|T047|AB|606.9|ICD9CM|Male infertility NOS|Male infertility NOS
C0021364|T047|PT|606.9|ICD9CM|Male infertility, unspecified|Male infertility, unspecified
C0030846|T047|HT|607|ICD9CM|Disorders of penis|Disorders of penis
C0022782|T047|AB|607.0|ICD9CM|Leukoplakia of penis|Leukoplakia of penis
C0022782|T047|PT|607.0|ICD9CM|Leukoplakia of penis|Leukoplakia of penis
C0004691|T047|AB|607.1|ICD9CM|Balanoposthitis|Balanoposthitis
C0004691|T047|PT|607.1|ICD9CM|Balanoposthitis|Balanoposthitis
C0156306|T047|AB|607.2|ICD9CM|Inflam dis, penis NEC|Inflam dis, penis NEC
C0156306|T047|PT|607.2|ICD9CM|Other inflammatory disorders of penis|Other inflammatory disorders of penis
C0033117|T047|AB|607.3|ICD9CM|Priapism|Priapism
C0033117|T047|PT|607.3|ICD9CM|Priapism|Priapism
C0029785|T047|HT|607.8|ICD9CM|Other specified disorders of penis|Other specified disorders of penis
C0152460|T047|AB|607.81|ICD9CM|Balanitis xerotica oblit|Balanitis xerotica oblit
C0152460|T047|PT|607.81|ICD9CM|Balanitis xerotica obliterans|Balanitis xerotica obliterans
C0156307|T047|AB|607.82|ICD9CM|Vascular disorder, penis|Vascular disorder, penis
C0156307|T047|PT|607.82|ICD9CM|Vascular disorders of penis|Vascular disorders of penis
C0156308|T046|AB|607.83|ICD9CM|Edema of penis|Edema of penis
C0156308|T046|PT|607.83|ICD9CM|Edema of penis|Edema of penis
C0156309|T046|PT|607.84|ICD9CM|Impotence of organic origin|Impotence of organic origin
C0156309|T046|AB|607.84|ICD9CM|Impotence, organic orign|Impotence, organic orign
C0030848|T047|AB|607.85|ICD9CM|Peyronie's disease|Peyronie's disease
C0030848|T047|PT|607.85|ICD9CM|Peyronie's disease|Peyronie's disease
C0029785|T047|AB|607.89|ICD9CM|Disorder of penis NEC|Disorder of penis NEC
C0029785|T047|PT|607.89|ICD9CM|Other specified disorders of penis|Other specified disorders of penis
C0030846|T047|AB|607.9|ICD9CM|Disorder of penis NOS|Disorder of penis NOS
C0030846|T047|PT|607.9|ICD9CM|Unspecified disorder of penis|Unspecified disorder of penis
C0156311|T047|HT|608|ICD9CM|Other disorders of male genital organs|Other disorders of male genital organs
C0042588|T047|AB|608.0|ICD9CM|Seminal vesiculitis|Seminal vesiculitis
C0042588|T047|PT|608.0|ICD9CM|Seminal vesiculitis|Seminal vesiculitis
C0037859|T047|AB|608.1|ICD9CM|Spermatocele|Spermatocele
C0037859|T047|PT|608.1|ICD9CM|Spermatocele|Spermatocele
C0037856|T047|HT|608.2|ICD9CM|Torsion of testis|Torsion of testis
C0037856|T047|AB|608.20|ICD9CM|Torsion of testis NOS|Torsion of testis NOS
C0037856|T047|PT|608.20|ICD9CM|Torsion of testis, unspecified|Torsion of testis, unspecified
C1719541|T046|AB|608.21|ICD9CM|Extravag tors sperm cord|Extravag tors sperm cord
C1719541|T046|PT|608.21|ICD9CM|Extravaginal torsion of spermatic cord|Extravaginal torsion of spermatic cord
C1719542|T047|AB|608.22|ICD9CM|Intravag tors sperm cord|Intravag tors sperm cord
C1719542|T047|PT|608.22|ICD9CM|Intravaginal torsion of spermatic cord|Intravaginal torsion of spermatic cord
C0392531|T190|AB|608.23|ICD9CM|Torsion appendix testis|Torsion appendix testis
C0392531|T190|PT|608.23|ICD9CM|Torsion of appendix testis|Torsion of appendix testis
C1997777|T047|AB|608.24|ICD9CM|Torsion appy epididymis|Torsion appy epididymis
C1997777|T047|PT|608.24|ICD9CM|Torsion of appendix epididymis|Torsion of appendix epididymis
C0156312|T047|AB|608.3|ICD9CM|Atrophy of testis|Atrophy of testis
C0156312|T047|PT|608.3|ICD9CM|Atrophy of testis|Atrophy of testis
C0156313|T047|AB|608.4|ICD9CM|Male gen inflam dis NEC|Male gen inflam dis NEC
C0156313|T047|PT|608.4|ICD9CM|Other inflammatory disorders of male genital organs|Other inflammatory disorders of male genital organs
C0029782|T047|HT|608.8|ICD9CM|Other specified disorders of male genital organs|Other specified disorders of male genital organs
C0156314|T047|PT|608.81|ICD9CM|Disorders of male genital organs in diseases classified elsewhere|Disorders of male genital organs in diseases classified elsewhere
C0156314|T047|AB|608.81|ICD9CM|Male gen dis in oth dis|Male gen dis in oth dis
C0149707|T033|AB|608.82|ICD9CM|Hematospermia|Hematospermia
C0149707|T033|PT|608.82|ICD9CM|Hematospermia|Hematospermia
C0042374|T047|AB|608.83|ICD9CM|Male gen vascul dis NEC|Male gen vascul dis NEC
C0042374|T047|PT|608.83|ICD9CM|Vascular disorders of male genital organs|Vascular disorders of male genital organs
C0156315|T047|PT|608.84|ICD9CM|Chylocele of tunica vaginalis|Chylocele of tunica vaginalis
C0156315|T047|AB|608.84|ICD9CM|Chylocele, tunic vaginal|Chylocele, tunic vaginal
C0156316|T190|PT|608.85|ICD9CM|Stricture of male genital organs|Stricture of male genital organs
C0156316|T190|AB|608.85|ICD9CM|Stricture, male gen orgn|Stricture, male gen orgn
C0156317|T184|PT|608.86|ICD9CM|Edema of male genital organs|Edema of male genital organs
C0156317|T184|AB|608.86|ICD9CM|Edema, male genital orgn|Edema, male genital orgn
C0403673|T046|AB|608.87|ICD9CM|Retrograde ejaculation|Retrograde ejaculation
C0403673|T046|PT|608.87|ICD9CM|Retrograde ejaculation|Retrograde ejaculation
C0029782|T047|AB|608.89|ICD9CM|Male genital dis NEC|Male genital dis NEC
C0029782|T047|PT|608.89|ICD9CM|Other specified disorders of male genital organs|Other specified disorders of male genital organs
C0017412|T047|AB|608.9|ICD9CM|Male genital dis NOS|Male genital dis NOS
C0017412|T047|PT|608.9|ICD9CM|Unspecified disorder of male genital organs|Unspecified disorder of male genital organs
C1305934|T046|HT|610|ICD9CM|Benign mammary dysplasias|Benign mammary dysplasias
C0006145|T047|HT|610-612.99|ICD9CM|DISORDERS OF BREAST|DISORDERS OF BREAST
C0037619|T190|AB|610.0|ICD9CM|Solitary cyst of breast|Solitary cyst of breast
C0037619|T190|PT|610.0|ICD9CM|Solitary cyst of breast|Solitary cyst of breast
C0016034|T047|AB|610.1|ICD9CM|Diffus cystic mastopathy|Diffus cystic mastopathy
C0016034|T047|PT|610.1|ICD9CM|Diffuse cystic mastopathy|Diffuse cystic mastopathy
C1305875|T047|AB|610.2|ICD9CM|Fibroadenosis of breast|Fibroadenosis of breast
C1305875|T047|PT|610.2|ICD9CM|Fibroadenosis of breast|Fibroadenosis of breast
C0156318|T047|AB|610.3|ICD9CM|Fibrosclerosis of breast|Fibrosclerosis of breast
C0156318|T047|PT|610.3|ICD9CM|Fibrosclerosis of breast|Fibrosclerosis of breast
C0152442|T047|AB|610.4|ICD9CM|Mammary duct ectasia|Mammary duct ectasia
C0152442|T047|PT|610.4|ICD9CM|Mammary duct ectasia|Mammary duct ectasia
C0156319|T047|AB|610.8|ICD9CM|Benign mamm dysplas NEC|Benign mamm dysplas NEC
C0156319|T047|PT|610.8|ICD9CM|Other specified benign mammary dysplasias|Other specified benign mammary dysplasias
C1305934|T046|AB|610.9|ICD9CM|Benign mamm dysplas NOS|Benign mamm dysplas NOS
C1305934|T046|PT|610.9|ICD9CM|Benign mammary dysplasia, unspecified|Benign mammary dysplasia, unspecified
C0156320|T047|HT|611|ICD9CM|Other disorders of breast|Other disorders of breast
C3495439|T047|AB|611.0|ICD9CM|Inflam disease of breast|Inflam disease of breast
C3495439|T047|PT|611.0|ICD9CM|Inflammatory disease of breast|Inflammatory disease of breast
C0020565|T046|AB|611.1|ICD9CM|Hypertrophy of breast|Hypertrophy of breast
C0020565|T046|PT|611.1|ICD9CM|Hypertrophy of breast|Hypertrophy of breast
C0152453|T033|AB|611.2|ICD9CM|Fissure of nipple|Fissure of nipple
C0152453|T033|PT|611.2|ICD9CM|Fissure of nipple|Fissure of nipple
C0156321|T047|AB|611.3|ICD9CM|Fat necrosis of breast|Fat necrosis of breast
C0156321|T047|PT|611.3|ICD9CM|Fat necrosis of breast|Fat necrosis of breast
C0151511|T020|AB|611.4|ICD9CM|Atrophy of breast|Atrophy of breast
C0151511|T020|PT|611.4|ICD9CM|Atrophy of breast|Atrophy of breast
C0152243|T020|AB|611.5|ICD9CM|Galactocele|Galactocele
C0152243|T020|PT|611.5|ICD9CM|Galactocele|Galactocele
C0235660|T047|PT|611.6|ICD9CM|Galactorrhea not associated with childbirth|Galactorrhea not associated with childbirth
C0235660|T047|AB|611.6|ICD9CM|Galactorrhea-nonobstet|Galactorrhea-nonobstet
C0156323|T184|HT|611.7|ICD9CM|Signs and symptoms in breast|Signs and symptoms in breast
C0024902|T184|AB|611.71|ICD9CM|Mastodynia|Mastodynia
C0024902|T184|PT|611.71|ICD9CM|Mastodynia|Mastodynia
C0024103|T033|AB|611.72|ICD9CM|Lump or mass in breast|Lump or mass in breast
C0024103|T033|PT|611.72|ICD9CM|Lump or mass in breast|Lump or mass in breast
C0156324|T184|PT|611.79|ICD9CM|Other signs and symptoms in breast|Other signs and symptoms in breast
C0156324|T184|AB|611.79|ICD9CM|Symptoms in breast NEC|Symptoms in breast NEC
C0156325|T047|HT|611.8|ICD9CM|Other specified disorders of breast|Other specified disorders of breast
C2233848|T033|PT|611.81|ICD9CM|Ptosis of breast|Ptosis of breast
C2233848|T033|AB|611.81|ICD9CM|Ptosis of breast|Ptosis of breast
C0266013|T019|PT|611.82|ICD9CM|Hypoplasia of breast|Hypoplasia of breast
C0266013|T019|AB|611.82|ICD9CM|Hypoplasia of breast|Hypoplasia of breast
C2349571|T047|AB|611.83|ICD9CM|Capslr contrctr brst imp|Capslr contrctr brst imp
C2349571|T047|PT|611.83|ICD9CM|Capsular contracture of breast implant|Capsular contracture of breast implant
C0156325|T047|AB|611.89|ICD9CM|Disorders breast NEC|Disorders breast NEC
C0156325|T047|PT|611.89|ICD9CM|Other specified disorders of breast|Other specified disorders of breast
C0006145|T047|AB|611.9|ICD9CM|Breast disorder NOS|Breast disorder NOS
C0006145|T047|PT|611.9|ICD9CM|Unspecified breast disorder|Unspecified breast disorder
C2349581|T047|HT|612|ICD9CM|Deformity and disproportion of reconstructed breast|Deformity and disproportion of reconstructed breast
C2349574|T047|PT|612.0|ICD9CM|Deformity of reconstructed breast|Deformity of reconstructed breast
C2349574|T047|AB|612.0|ICD9CM|Deformity reconst breast|Deformity reconst breast
C2349578|T047|PT|612.1|ICD9CM|Disproportion of reconstructed breast|Disproportion of reconstructed breast
C2349578|T047|AB|612.1|ICD9CM|Disproportn reconst brst|Disproportn reconst brst
C0156326|T047|HT|614|ICD9CM|Inflammatory disease of ovary, fallopian tube, pelvic cellular tissue, and peritoneum|Inflammatory disease of ovary, fallopian tube, pelvic cellular tissue, and peritoneum
C0242172|T047|HT|614-616.99|ICD9CM|INFLAMMATORY DISEASE OF FEMALE PELVIC ORGANS|INFLAMMATORY DISEASE OF FEMALE PELVIC ORGANS
C0156327|T047|AB|614.0|ICD9CM|Ac salpingo-oophoritis|Ac salpingo-oophoritis
C0156327|T047|PT|614.0|ICD9CM|Acute salpingitis and oophoritis|Acute salpingitis and oophoritis
C0156328|T047|AB|614.1|ICD9CM|Chr salpingo-oophoritis|Chr salpingo-oophoritis
C0156328|T047|PT|614.1|ICD9CM|Chronic salpingitis and oophoritis|Chronic salpingitis and oophoritis
C0036133|T047|PT|614.2|ICD9CM|Salpingitis and oophoritis not specified as acute, subacute, or chronic|Salpingitis and oophoritis not specified as acute, subacute, or chronic
C0036133|T047|AB|614.2|ICD9CM|Salpingo-oophoritis NOS|Salpingo-oophoritis NOS
C0156329|T047|AB|614.3|ICD9CM|Acute parametritis|Acute parametritis
C0156329|T047|PT|614.3|ICD9CM|Acute parametritis and pelvic cellulitis|Acute parametritis and pelvic cellulitis
C0404458|T047|PT|614.4|ICD9CM|Chronic or unspecified parametritis and pelvic cellulitis|Chronic or unspecified parametritis and pelvic cellulitis
C0404458|T047|AB|614.4|ICD9CM|Chronic parametritis|Chronic parametritis
C0269032|T047|AB|614.5|ICD9CM|Ac pelv peritonitis-fem|Ac pelv peritonitis-fem
C0269032|T047|PT|614.5|ICD9CM|Acute or unspecified pelvic peritonitis, female|Acute or unspecified pelvic peritonitis, female
C0375384|T020|AB|614.6|ICD9CM|Fem pelvic periton adhes|Fem pelvic periton adhes
C0375384|T020|PT|614.6|ICD9CM|Pelvic peritoneal adhesions, female (postoperative) (postinfection)|Pelvic peritoneal adhesions, female (postoperative) (postinfection)
C0156332|T047|AB|614.7|ICD9CM|Chr pelv periton NEC-fem|Chr pelv periton NEC-fem
C0156332|T047|PT|614.7|ICD9CM|Other chronic pelvic peritonitis, female|Other chronic pelvic peritonitis, female
C0029807|T047|AB|614.8|ICD9CM|Fem pelv inflam dis NEC|Fem pelv inflam dis NEC
C0029807|T047|PT|614.8|ICD9CM|Other specified inflammatory disease of female pelvic organs and tissues|Other specified inflammatory disease of female pelvic organs and tissues
C0242172|T047|AB|614.9|ICD9CM|Fem pelv inflam dis NOS|Fem pelv inflam dis NOS
C0242172|T047|PT|614.9|ICD9CM|Unspecified inflammatory disease of female pelvic organs and tissues|Unspecified inflammatory disease of female pelvic organs and tissues
C0156333|T047|HT|615|ICD9CM|Inflammatory diseases of uterus, except cervix|Inflammatory diseases of uterus, except cervix
C0156334|T047|AB|615.0|ICD9CM|Ac uterine inflammation|Ac uterine inflammation
C0156334|T047|PT|615.0|ICD9CM|Acute inflammatory diseases of uterus, except cervix|Acute inflammatory diseases of uterus, except cervix
C0156335|T047|AB|615.1|ICD9CM|Chr uterine inflammation|Chr uterine inflammation
C0156335|T047|PT|615.1|ICD9CM|Chronic inflammatory diseases of uterus, except cervix|Chronic inflammatory diseases of uterus, except cervix
C0269047|T047|PT|615.9|ICD9CM|Unspecified inflammatory disease of uterus|Unspecified inflammatory disease of uterus
C0269047|T047|AB|615.9|ICD9CM|Uterine inflam dis NOS|Uterine inflam dis NOS
C0156342|T047|HT|616|ICD9CM|Inflammatory disease of cervix, vagina, and vulva|Inflammatory disease of cervix, vagina, and vulva
C0007861|T047|AB|616.0|ICD9CM|Cervicitis|Cervicitis
C0007861|T047|PT|616.0|ICD9CM|Cervicitis and endocervicitis|Cervicitis and endocervicitis
C0042268|T047|HT|616.1|ICD9CM|Vaginitis and vulvovaginitis|Vaginitis and vulvovaginitis
C0042268|T047|PT|616.10|ICD9CM|Vaginitis and vulvovaginitis, unspecified|Vaginitis and vulvovaginitis, unspecified
C0042268|T047|AB|616.10|ICD9CM|Vaginitis NOS|Vaginitis NOS
C0156337|T047|PT|616.11|ICD9CM|Vaginitis and vulvovaginitis in diseases classified elsewhere|Vaginitis and vulvovaginitis in diseases classified elsewhere
C0156337|T047|AB|616.11|ICD9CM|Vaginitis in oth disease|Vaginitis in oth disease
C0004767|T047|AB|616.2|ICD9CM|Bartholin's gland cyst|Bartholin's gland cyst
C0004767|T047|PT|616.2|ICD9CM|Cyst of Bartholin's gland|Cyst of Bartholin's gland
C0004766|T046|PT|616.3|ICD9CM|Abscess of Bartholin's gland|Abscess of Bartholin's gland
C0004766|T046|AB|616.3|ICD9CM|Bartholin's glnd abscess|Bartholin's glnd abscess
C0156338|T047|AB|616.4|ICD9CM|Abscess of vulva NEC|Abscess of vulva NEC
C0156338|T047|PT|616.4|ICD9CM|Other abscess of vulva|Other abscess of vulva
C0156339|T047|HT|616.5|ICD9CM|Ulceration of vulva|Ulceration of vulva
C0156339|T047|AB|616.50|ICD9CM|Ulceration of vulva NOS|Ulceration of vulva NOS
C0156339|T047|PT|616.50|ICD9CM|Ulceration of vulva, unspecified|Ulceration of vulva, unspecified
C0156340|T047|PT|616.51|ICD9CM|Ulceration of vulva in diseases classified elsewhere|Ulceration of vulva in diseases classified elsewhere
C0156340|T047|AB|616.51|ICD9CM|Vulvar ulcer in oth dis|Vulvar ulcer in oth dis
C0156341|T047|HT|616.8|ICD9CM|Other specified inflammatory diseases of cervix, vagina, and vulva|Other specified inflammatory diseases of cervix, vagina, and vulva
C1719543|T047|PT|616.81|ICD9CM|Mucositis (ulcerative) of cervix, vagina, and vulva|Mucositis (ulcerative) of cervix, vagina, and vulva
C1719543|T047|AB|616.81|ICD9CM|Mucositis cerv,vag,vulva|Mucositis cerv,vag,vulva
C1719544|T047|AB|616.89|ICD9CM|Inflm cerv,vag,vulva NEC|Inflm cerv,vag,vulva NEC
C1719544|T047|PT|616.89|ICD9CM|Other inflammatory disease of cervix, vagina and vulva|Other inflammatory disease of cervix, vagina and vulva
C0156342|T047|AB|616.9|ICD9CM|Female gen inflam NOS|Female gen inflam NOS
C0156342|T047|PT|616.9|ICD9CM|Unspecified inflammatory disease of cervix, vagina, and vulva|Unspecified inflammatory disease of cervix, vagina, and vulva
C0014175|T047|HT|617|ICD9CM|Endometriosis|Endometriosis
C0178291|T047|HT|617-629.99|ICD9CM|OTHER DISORDERS OF FEMALE GENITAL TRACT|OTHER DISORDERS OF FEMALE GENITAL TRACT
C0341858|T047|PT|617.0|ICD9CM|Endometriosis of uterus|Endometriosis of uterus
C0341858|T047|AB|617.0|ICD9CM|Uterine endometriosis|Uterine endometriosis
C0156344|T047|PT|617.1|ICD9CM|Endometriosis of ovary|Endometriosis of ovary
C0156344|T047|AB|617.1|ICD9CM|Ovarian endometriosis|Ovarian endometriosis
C0014177|T047|PT|617.2|ICD9CM|Endometriosis of fallopian tube|Endometriosis of fallopian tube
C0014177|T047|AB|617.2|ICD9CM|Tubal endometriosis|Tubal endometriosis
C0156345|T047|PT|617.3|ICD9CM|Endometriosis of pelvic peritoneum|Endometriosis of pelvic peritoneum
C0156345|T047|AB|617.3|ICD9CM|Pelv perit endometriosis|Pelv perit endometriosis
C0156346|T047|PT|617.4|ICD9CM|Endometriosis of rectovaginal septum and vagina|Endometriosis of rectovaginal septum and vagina
C0156346|T047|AB|617.4|ICD9CM|Vaginal endometriosis|Vaginal endometriosis
C0156347|T047|PT|617.5|ICD9CM|Endometriosis of intestine|Endometriosis of intestine
C0156347|T047|AB|617.5|ICD9CM|Intestinal endometriosis|Intestinal endometriosis
C0156348|T047|AB|617.6|ICD9CM|Endometriosis in scar|Endometriosis in scar
C0156348|T047|PT|617.6|ICD9CM|Endometriosis in scar of skin|Endometriosis in scar of skin
C0014178|T047|AB|617.8|ICD9CM|Endometriosis NEC|Endometriosis NEC
C0014178|T047|PT|617.8|ICD9CM|Endometriosis of other specified sites|Endometriosis of other specified sites
C0014175|T047|AB|617.9|ICD9CM|Endometriosis NOS|Endometriosis NOS
C0014175|T047|PT|617.9|ICD9CM|Endometriosis, site unspecified|Endometriosis, site unspecified
C0156349|T047|HT|618|ICD9CM|Genital prolapse|Genital prolapse
C0156350|T020|HT|618.0|ICD9CM|Prolapse of vaginal walls without mention of uterine prolapse|Prolapse of vaginal walls without mention of uterine prolapse
C1456247|T047|PT|618.00|ICD9CM|Unspecified prolapse of vaginal walls|Unspecified prolapse of vaginal walls
C1456247|T047|AB|618.00|ICD9CM|Vaginal wall prolpse NOS|Vaginal wall prolpse NOS
C1456248|T047|AB|618.01|ICD9CM|Cystocele, midline|Cystocele, midline
C1456248|T047|PT|618.01|ICD9CM|Cystocele, midline|Cystocele, midline
C2711750|T047|AB|618.02|ICD9CM|Cystocele, lateral|Cystocele, lateral
C2711750|T047|PT|618.02|ICD9CM|Cystocele, lateral|Cystocele, lateral
C0238502|T047|AB|618.03|ICD9CM|Urethrocele|Urethrocele
C0238502|T047|PT|618.03|ICD9CM|Urethrocele|Urethrocele
C0149771|T020|AB|618.04|ICD9CM|Rectocele|Rectocele
C0149771|T020|PT|618.04|ICD9CM|Rectocele|Rectocele
C1456251|T047|AB|618.05|ICD9CM|Perineocele|Perineocele
C1456251|T047|PT|618.05|ICD9CM|Perineocele|Perineocele
C1456252|T047|AB|618.09|ICD9CM|Cystourethrocele|Cystourethrocele
C1456252|T047|PT|618.09|ICD9CM|Other prolapse of vaginal walls without mention of uterine prolapse|Other prolapse of vaginal walls without mention of uterine prolapse
C0553716|T020|AB|618.1|ICD9CM|Uterine prolapse|Uterine prolapse
C0553716|T020|PT|618.1|ICD9CM|Uterine prolapse without mention of vaginal wall prolapse|Uterine prolapse without mention of vaginal wall prolapse
C0156351|T020|AB|618.2|ICD9CM|Uterovag prolaps-incompl|Uterovag prolaps-incompl
C0156351|T020|PT|618.2|ICD9CM|Uterovaginal prolapse, incomplete|Uterovaginal prolapse, incomplete
C0392530|T020|AB|618.3|ICD9CM|Uterovag prolaps-complet|Uterovag prolaps-complet
C0392530|T020|PT|618.3|ICD9CM|Uterovaginal prolapse, complete|Uterovaginal prolapse, complete
C0156353|T020|PT|618.4|ICD9CM|Uterovaginal prolapse, unspecified|Uterovaginal prolapse, unspecified
C0156353|T020|AB|618.4|ICD9CM|Utervaginal prolapse NOS|Utervaginal prolapse NOS
C0156354|T020|AB|618.5|ICD9CM|Postop vaginal prolapse|Postop vaginal prolapse
C0156354|T020|PT|618.5|ICD9CM|Prolapse of vaginal vault after hysterectomy|Prolapse of vaginal vault after hysterectomy
C0205792|T190|AB|618.6|ICD9CM|Vaginal enterocele|Vaginal enterocele
C0205792|T190|PT|618.6|ICD9CM|Vaginal enterocele, congenital or acquired|Vaginal enterocele, congenital or acquired
C0156355|T037|AB|618.7|ICD9CM|Old lacer pelvic muscle|Old lacer pelvic muscle
C0156355|T037|PT|618.7|ICD9CM|Old laceration of muscles of pelvic floor|Old laceration of muscles of pelvic floor
C0029801|T047|HT|618.8|ICD9CM|Other specified genital prolapse|Other specified genital prolapse
C1456253|T047|PT|618.81|ICD9CM|Incompetence or weakening of pubocervical tissue|Incompetence or weakening of pubocervical tissue
C1456253|T047|AB|618.81|ICD9CM|Incomptnce pubocerv tiss|Incomptnce pubocerv tiss
C1456254|T047|PT|618.82|ICD9CM|Incompetence or weakening of rectovaginal tissue|Incompetence or weakening of rectovaginal tissue
C1456254|T047|AB|618.82|ICD9CM|Incomptnce rectovag tiss|Incomptnce rectovag tiss
C1456255|T047|AB|618.83|ICD9CM|Pelvic muscle wasting|Pelvic muscle wasting
C1456255|T047|PT|618.83|ICD9CM|Pelvic muscle wasting|Pelvic muscle wasting
C1719546|T020|PT|618.84|ICD9CM|Cervical stump prolapse|Cervical stump prolapse
C1719546|T020|AB|618.84|ICD9CM|Cervical stump prolapse|Cervical stump prolapse
C0029801|T047|AB|618.89|ICD9CM|Genital prolapse NEC|Genital prolapse NEC
C0029801|T047|PT|618.89|ICD9CM|Other specified genital prolapse|Other specified genital prolapse
C0156356|T020|AB|618.9|ICD9CM|Genital prolapse NOS|Genital prolapse NOS
C0156356|T020|PT|618.9|ICD9CM|Unspecified genital prolapse|Unspecified genital prolapse
C0156357|T190|HT|619|ICD9CM|Fistula involving female genital tract|Fistula involving female genital tract
C0042033|T047|AB|619.0|ICD9CM|Urin-genital fistul, fem|Urin-genital fistul, fem
C0042033|T047|PT|619.0|ICD9CM|Urinary-genital tract fistula, female|Urinary-genital tract fistula, female
C0012246|T190|AB|619.1|ICD9CM|Digest-genit fistul, fem|Digest-genit fistul, fem
C0012246|T190|PT|619.1|ICD9CM|Digestive-genital tract fistula, female|Digestive-genital tract fistula, female
C0156358|T020|PT|619.2|ICD9CM|Genital tract-skin fistula, female|Genital tract-skin fistula, female
C0156358|T020|AB|619.2|ICD9CM|Genital-skin fistul, fem|Genital-skin fistul, fem
C0029797|T190|AB|619.8|ICD9CM|Fem genital fistula NEC|Fem genital fistula NEC
C0029797|T190|PT|619.8|ICD9CM|Other specified fistulas involving female genital tract|Other specified fistulas involving female genital tract
C0269131|T190|AB|619.9|ICD9CM|Fem genital fistula NOS|Fem genital fistula NOS
C0269131|T190|PT|619.9|ICD9CM|Unspecified fistula involving female genital tract|Unspecified fistula involving female genital tract
C0156367|T047|HT|620|ICD9CM|Noninflammatory disorders of ovary, fallopian tube, and broad ligament|Noninflammatory disorders of ovary, fallopian tube, and broad ligament
C0016429|T047|AB|620.0|ICD9CM|Follicular cyst of ovary|Follicular cyst of ovary
C0016429|T047|PT|620.0|ICD9CM|Follicular cyst of ovary|Follicular cyst of ovary
C0156361|T047|AB|620.1|ICD9CM|Corpus luteum cyst|Corpus luteum cyst
C0156361|T047|PT|620.1|ICD9CM|Corpus luteum cyst or hematoma|Corpus luteum cyst or hematoma
C0029513|T020|PT|620.2|ICD9CM|Other and unspecified ovarian cyst|Other and unspecified ovarian cyst
C0029513|T020|AB|620.2|ICD9CM|Ovarian cyst NEC/NOS|Ovarian cyst NEC/NOS
C0156362|T020|AB|620.3|ICD9CM|Acq atrophy ovary & tube|Acq atrophy ovary & tube
C0156362|T020|PT|620.3|ICD9CM|Acquired atrophy of ovary and fallopian tube|Acquired atrophy of ovary and fallopian tube
C0495094|T020|AB|620.4|ICD9CM|Prolapse of ovary & tube|Prolapse of ovary & tube
C0495094|T020|PT|620.4|ICD9CM|Prolapse or hernia of ovary and fallopian tube|Prolapse or hernia of ovary and fallopian tube
C0156364|T190|AB|620.5|ICD9CM|Torsion of ovary or tube|Torsion of ovary or tube
C0156364|T190|PT|620.5|ICD9CM|Torsion of ovary, ovarian pedicle, or fallopian tube|Torsion of ovary, ovarian pedicle, or fallopian tube
C0152079|T047|AB|620.6|ICD9CM|Broad ligament lacer syn|Broad ligament lacer syn
C0152079|T047|PT|620.6|ICD9CM|Broad ligament laceration syndrome|Broad ligament laceration syndrome
C0156365|T046|AB|620.7|ICD9CM|Broad ligament hematoma|Broad ligament hematoma
C0156365|T046|PT|620.7|ICD9CM|Hematoma of broad ligament|Hematoma of broad ligament
C0156366|T047|AB|620.8|ICD9CM|Noninfl dis ova/adnx NEC|Noninfl dis ova/adnx NEC
C0156366|T047|PT|620.8|ICD9CM|Other noninflammatory disorders of ovary, fallopian tube, and broad ligament|Other noninflammatory disorders of ovary, fallopian tube, and broad ligament
C0156367|T047|AB|620.9|ICD9CM|Noninfl dis ova/adnx NOS|Noninfl dis ova/adnx NOS
C0156367|T047|PT|620.9|ICD9CM|Unspecified noninflammatory disorder of ovary, fallopian tube, and broad ligament|Unspecified noninflammatory disorder of ovary, fallopian tube, and broad ligament
C0868853|T047|HT|621|ICD9CM|Disorders of uterus, not elsewhere classified|Disorders of uterus, not elsewhere classified
C0156369|T191|AB|621.0|ICD9CM|Polyp of corpus uteri|Polyp of corpus uteri
C0156369|T191|PT|621.0|ICD9CM|Polyp of corpus uteri|Polyp of corpus uteri
C0156370|T047|AB|621.1|ICD9CM|Chr uterine subinvolutn|Chr uterine subinvolutn
C0156370|T047|PT|621.1|ICD9CM|Chronic subinvolution of uterus|Chronic subinvolution of uterus
C0156371|T033|AB|621.2|ICD9CM|Hypertrophy of uterus|Hypertrophy of uterus
C0156371|T033|PT|621.2|ICD9CM|Hypertrophy of uterus|Hypertrophy of uterus
C0014173|T047|HT|621.3|ICD9CM|Endometrial hyperplasia|Endometrial hyperplasia
C0014173|T047|AB|621.30|ICD9CM|Endometrial hyperpla NOS|Endometrial hyperpla NOS
C0014173|T047|PT|621.30|ICD9CM|Endometrial hyperplasia, unspecified|Endometrial hyperplasia, unspecified
C1335967|T046|AB|621.31|ICD9CM|Simp endo hyper w/o atyp|Simp endo hyper w/o atyp
C1335967|T046|PT|621.31|ICD9CM|Simple endometrial hyperplasia without atypia|Simple endometrial hyperplasia without atypia
C1333139|T046|AB|621.32|ICD9CM|Comp endo hyper w/o atyp|Comp endo hyper w/o atyp
C1333139|T046|PT|621.32|ICD9CM|Complex endometrial hyperplasia without atypia|Complex endometrial hyperplasia without atypia
C0349579|T047|AB|621.33|ICD9CM|Endomet hyperpla w atyp|Endomet hyperpla w atyp
C0349579|T047|PT|621.33|ICD9CM|Endometrial hyperplasia with atypia|Endometrial hyperplasia with atypia
C2712711|T047|AB|621.34|ICD9CM|Ben endomet hyperplasia|Ben endomet hyperplasia
C2712711|T047|PT|621.34|ICD9CM|Benign endometrial hyperplasia|Benign endometrial hyperplasia
C1333394|T191|AB|621.35|ICD9CM|Endomet intraepithl neop|Endomet intraepithl neop
C1333394|T191|PT|621.35|ICD9CM|Endometrial intraepithelial neoplasia [EIN]|Endometrial intraepithelial neoplasia [EIN]
C0018948|T046|AB|621.4|ICD9CM|Hematometra|Hematometra
C0018948|T046|PT|621.4|ICD9CM|Hematometra|Hematometra
C1704274|T047|AB|621.5|ICD9CM|Intrauterine synechiae|Intrauterine synechiae
C1704274|T047|PT|621.5|ICD9CM|Intrauterine synechiae|Intrauterine synechiae
C0156373|T033|AB|621.6|ICD9CM|Malposition of uterus|Malposition of uterus
C0156373|T033|PT|621.6|ICD9CM|Malposition of uterus|Malposition of uterus
C0156374|T047|AB|621.7|ICD9CM|Chr inversion of uterus|Chr inversion of uterus
C0156374|T047|PT|621.7|ICD9CM|Chronic inversion of uterus|Chronic inversion of uterus
C0302384|T047|AB|621.8|ICD9CM|Disorders of uterus NEC|Disorders of uterus NEC
C0302384|T047|PT|621.8|ICD9CM|Other specified disorders of uterus, not elsewhere classified|Other specified disorders of uterus, not elsewhere classified
C0042131|T047|AB|621.9|ICD9CM|Disorder of uterus NOS|Disorder of uterus NOS
C0042131|T047|PT|621.9|ICD9CM|Unspecified disorder of uterus|Unspecified disorder of uterus
C0156377|T047|HT|622|ICD9CM|Noninflammatory disorders of cervix|Noninflammatory disorders of cervix
C0014719|T020|PT|622.0|ICD9CM|Erosion and ectropion of cervix|Erosion and ectropion of cervix
C0014719|T020|AB|622.0|ICD9CM|Erosion/ectropion cervix|Erosion/ectropion cervix
C0007868|T047|HT|622.1|ICD9CM|Dysplasia of cervix (uteri)|Dysplasia of cervix (uteri)
C0007868|T047|AB|622.10|ICD9CM|Dysplasia of cervix NOS|Dysplasia of cervix NOS
C0007868|T047|PT|622.10|ICD9CM|Dysplasia of cervix, unspecified|Dysplasia of cervix, unspecified
C0349458|T191|AB|622.11|ICD9CM|Mild dysplasia of cervix|Mild dysplasia of cervix
C0349458|T191|PT|622.11|ICD9CM|Mild dysplasia of cervix|Mild dysplasia of cervix
C0349459|T191|AB|622.12|ICD9CM|Mod dysplasia of cervix|Mod dysplasia of cervix
C0349459|T191|PT|622.12|ICD9CM|Moderate dysplasia of cervix|Moderate dysplasia of cervix
C0269194|T191|AB|622.2|ICD9CM|Leukoplakia of cervix|Leukoplakia of cervix
C0269194|T191|PT|622.2|ICD9CM|Leukoplakia of cervix (uteri)|Leukoplakia of cervix (uteri)
C0156379|T037|AB|622.3|ICD9CM|Old laceration of cervix|Old laceration of cervix
C0156379|T037|PT|622.3|ICD9CM|Old laceration of cervix|Old laceration of cervix
C0156380|T190|PT|622.4|ICD9CM|Stricture and stenosis of cervix|Stricture and stenosis of cervix
C0156380|T190|AB|622.4|ICD9CM|Stricture of cervix|Stricture of cervix
C0007871|T046|AB|622.5|ICD9CM|Incompetence of cervix|Incompetence of cervix
C0007871|T046|PT|622.5|ICD9CM|Incompetence of cervix|Incompetence of cervix
C0020561|T047|AB|622.6|ICD9CM|Hypertrophic elong cervx|Hypertrophic elong cervx
C0020561|T047|PT|622.6|ICD9CM|Hypertrophic elongation of cervix|Hypertrophic elongation of cervix
C0026725|T191|AB|622.7|ICD9CM|Mucous polyp of cervix|Mucous polyp of cervix
C0026725|T191|PT|622.7|ICD9CM|Mucous polyp of cervix|Mucous polyp of cervix
C0477784|T047|AB|622.8|ICD9CM|Noninflam dis cervix NEC|Noninflam dis cervix NEC
C0477784|T047|PT|622.8|ICD9CM|Other specified noninflammatory disorders of cervix|Other specified noninflammatory disorders of cervix
C0156377|T047|AB|622.9|ICD9CM|Noninflam dis cervix NOS|Noninflam dis cervix NOS
C0156377|T047|PT|622.9|ICD9CM|Unspecified noninflammatory disorder of cervix|Unspecified noninflammatory disorder of cervix
C0156383|T047|HT|623|ICD9CM|Noninflammatory disorders of vagina|Noninflammatory disorders of vagina
C0156384|T046|AB|623.0|ICD9CM|Dysplasia of vagina|Dysplasia of vagina
C0156384|T046|PT|623.0|ICD9CM|Dysplasia of vagina|Dysplasia of vagina
C0156385|T191|AB|623.1|ICD9CM|Leukoplakia of vagina|Leukoplakia of vagina
C0156385|T191|PT|623.1|ICD9CM|Leukoplakia of vagina|Leukoplakia of vagina
C0156386|T190|AB|623.2|ICD9CM|Stricture of vagina|Stricture of vagina
C0156386|T190|PT|623.2|ICD9CM|Stricture or atresia of vagina|Stricture or atresia of vagina
C0156387|T190|AB|623.3|ICD9CM|Tight hymenal ring|Tight hymenal ring
C0156387|T190|PT|623.3|ICD9CM|Tight hymenal ring|Tight hymenal ring
C0156388|T033|AB|623.4|ICD9CM|Old vaginal laceration|Old vaginal laceration
C0156388|T033|PT|623.4|ICD9CM|Old vaginal laceration|Old vaginal laceration
C0023534|T047|PT|623.5|ICD9CM|Leukorrhea, not specified as infective|Leukorrhea, not specified as infective
C0023534|T047|AB|623.5|ICD9CM|Noninfect vag leukorrhea|Noninfect vag leukorrhea
C0156389|T046|AB|623.6|ICD9CM|Vaginal hematoma|Vaginal hematoma
C0156389|T046|PT|623.6|ICD9CM|Vaginal hematoma|Vaginal hematoma
C0156390|T191|AB|623.7|ICD9CM|Polyp of vagina|Polyp of vagina
C0156390|T191|PT|623.7|ICD9CM|Polyp of vagina|Polyp of vagina
C0029819|T047|AB|623.8|ICD9CM|Noninflam dis vagina NEC|Noninflam dis vagina NEC
C0029819|T047|PT|623.8|ICD9CM|Other specified noninflammatory disorders of vagina|Other specified noninflammatory disorders of vagina
C0156383|T047|AB|623.9|ICD9CM|Noninflam dis vagina NOS|Noninflam dis vagina NOS
C0156383|T047|PT|623.9|ICD9CM|Unspecified noninflammatory disorder of vagina|Unspecified noninflammatory disorder of vagina
C0156400|T047|HT|624|ICD9CM|Noninflammatory disorders of vulva and perineum|Noninflammatory disorders of vulva and perineum
C0013426|T047|HT|624.0|ICD9CM|Dystrophy of vulva|Dystrophy of vulva
C0495106|T191|AB|624.01|ICD9CM|Vulvar intraeph neopl I|Vulvar intraeph neopl I
C0495106|T191|PT|624.01|ICD9CM|Vulvar intraepithelial neoplasia I [VIN I]|Vulvar intraepithelial neoplasia I [VIN I]
C0495107|T191|PT|624.02|ICD9CM|Vulvar intraepithelial neoplasia II [VIN II]|Vulvar intraepithelial neoplasia II [VIN II]
C0495107|T191|AB|624.02|ICD9CM|Vulvr intraepth neopl II|Vulvr intraepth neopl II
C1955816|T047|AB|624.09|ICD9CM|Dystrophy of vulva NEC|Dystrophy of vulva NEC
C1955816|T047|PT|624.09|ICD9CM|Other dystrophy of vulva|Other dystrophy of vulva
C0156393|T047|AB|624.1|ICD9CM|Atrophy of vulva|Atrophy of vulva
C0156393|T047|PT|624.1|ICD9CM|Atrophy of vulva|Atrophy of vulva
C0156394|T047|AB|624.2|ICD9CM|Hypertrophy of clitoris|Hypertrophy of clitoris
C0156394|T047|PT|624.2|ICD9CM|Hypertrophy of clitoris|Hypertrophy of clitoris
C0404531|T046|AB|624.3|ICD9CM|Hypertrophy of labia|Hypertrophy of labia
C0404531|T046|PT|624.3|ICD9CM|Hypertrophy of labia|Hypertrophy of labia
C0269223|T037|AB|624.4|ICD9CM|Old laceration of vulva|Old laceration of vulva
C0269223|T037|PT|624.4|ICD9CM|Old laceration or scarring of vulva|Old laceration or scarring of vulva
C0156397|T046|AB|624.5|ICD9CM|Hematoma of vulva|Hematoma of vulva
C0156397|T046|PT|624.5|ICD9CM|Hematoma of vulva|Hematoma of vulva
C0156398|T047|AB|624.6|ICD9CM|Polyp of labia and vulva|Polyp of labia and vulva
C0156398|T047|PT|624.6|ICD9CM|Polyp of labia and vulva|Polyp of labia and vulva
C0156399|T047|AB|624.8|ICD9CM|Noninflam dis vulva NEC|Noninflam dis vulva NEC
C0156399|T047|PT|624.8|ICD9CM|Other specified noninflammatory disorders of vulva and perineum|Other specified noninflammatory disorders of vulva and perineum
C0156400|T047|AB|624.9|ICD9CM|Noninflam dis vulva NOS|Noninflam dis vulva NOS
C0156400|T047|PT|624.9|ICD9CM|Unspecified noninflammatory disorder of vulva and perineum|Unspecified noninflammatory disorder of vulva and perineum
C0156401|T184|HT|625|ICD9CM|Pain and other symptoms associated with female genital organs|Pain and other symptoms associated with female genital organs
C0013394|T047|AB|625.0|ICD9CM|Dyspareunia|Dyspareunia
C0013394|T047|PT|625.0|ICD9CM|Dyspareunia|Dyspareunia
C2004487|T047|AB|625.1|ICD9CM|Vaginismus|Vaginismus
C2004487|T047|PT|625.1|ICD9CM|Vaginismus|Vaginismus
C0152149|T184|AB|625.2|ICD9CM|Mittelschmerz|Mittelschmerz
C0152149|T184|PT|625.2|ICD9CM|Mittelschmerz|Mittelschmerz
C0013390|T047|AB|625.3|ICD9CM|Dysmenorrhea|Dysmenorrhea
C0013390|T047|PT|625.3|ICD9CM|Dysmenorrhea|Dysmenorrhea
C0376356|T047|AB|625.4|ICD9CM|Premenstrual tension|Premenstrual tension
C0376356|T047|PT|625.4|ICD9CM|Premenstrual tension syndromes|Premenstrual tension syndromes
C0152078|T047|AB|625.5|ICD9CM|Pelvic congestion synd|Pelvic congestion synd
C0152078|T047|PT|625.5|ICD9CM|Pelvic congestion syndrome|Pelvic congestion syndrome
C0038437|T047|AB|625.6|ICD9CM|Fem stress incontinence|Fem stress incontinence
C0038437|T047|PT|625.6|ICD9CM|Stress incontinence, female|Stress incontinence, female
C0406670|T047|HT|625.7|ICD9CM|Vulvodynia|Vulvodynia
C0406670|T047|AB|625.70|ICD9CM|Vulvodynia NOS|Vulvodynia NOS
C0406670|T047|PT|625.70|ICD9CM|Vulvodynia, unspecified|Vulvodynia, unspecified
C0269084|T047|PT|625.71|ICD9CM|Vulvar vestibulitis|Vulvar vestibulitis
C0269084|T047|AB|625.71|ICD9CM|Vulvar vestibulitis|Vulvar vestibulitis
C2349583|T047|PT|625.79|ICD9CM|Other vulvodynia|Other vulvodynia
C2349583|T047|AB|625.79|ICD9CM|Other vulvodynia|Other vulvodynia
C0156402|T184|AB|625.8|ICD9CM|Fem genital symptoms NEC|Fem genital symptoms NEC
C0156402|T184|PT|625.8|ICD9CM|Other specified symptoms associated with female genital organs|Other specified symptoms associated with female genital organs
C0041889|T184|AB|625.9|ICD9CM|Fem genital symptoms NOS|Fem genital symptoms NOS
C0041889|T184|PT|625.9|ICD9CM|Unspecified symptom associated with female genital organs|Unspecified symptom associated with female genital organs
C0041827|T047|HT|626|ICD9CM|Disorders of menstruation and other abnormal bleeding from female genital tract|Disorders of menstruation and other abnormal bleeding from female genital tract
C0002453|T033|AB|626.0|ICD9CM|Absence of menstruation|Absence of menstruation
C0002453|T033|PT|626.0|ICD9CM|Absence of menstruation|Absence of menstruation
C0404550|T033|AB|626.1|ICD9CM|Scanty menstruation|Scanty menstruation
C0404550|T033|PT|626.1|ICD9CM|Scanty or infrequent menstruation|Scanty or infrequent menstruation
C0341863|T046|AB|626.2|ICD9CM|Excessive menstruation|Excessive menstruation
C0341863|T046|PT|626.2|ICD9CM|Excessive or frequent menstruation|Excessive or frequent menstruation
C0156403|T046|AB|626.3|ICD9CM|Pubertal menorrhagia|Pubertal menorrhagia
C0156403|T046|PT|626.3|ICD9CM|Puberty bleeding|Puberty bleeding
C0156404|T033|PT|626.4|ICD9CM|Irregular menstrual cycle|Irregular menstrual cycle
C0156404|T033|AB|626.4|ICD9CM|Irregular menstruation|Irregular menstruation
C0156405|T184|AB|626.5|ICD9CM|Ovulation bleeding|Ovulation bleeding
C0156405|T184|PT|626.5|ICD9CM|Ovulation bleeding|Ovulation bleeding
C0025874|T046|AB|626.6|ICD9CM|Metrorrhagia|Metrorrhagia
C0025874|T046|PT|626.6|ICD9CM|Metrorrhagia|Metrorrhagia
C0156406|T046|AB|626.7|ICD9CM|Postcoital bleeding|Postcoital bleeding
C0156406|T046|PT|626.7|ICD9CM|Postcoital bleeding|Postcoital bleeding
C0029592|T033|AB|626.8|ICD9CM|Menstrual disorder NEC|Menstrual disorder NEC
C0029592|T033|PT|626.8|ICD9CM|Other disorders of menstruation and other abnormal bleeding from female genital tract|Other disorders of menstruation and other abnormal bleeding from female genital tract
C0041827|T047|AB|626.9|ICD9CM|Menstrual disorder NOS|Menstrual disorder NOS
C0041827|T047|PT|626.9|ICD9CM|Unspecified disorders of menstruation and other abnormal bleeding from female genital tract|Unspecified disorders of menstruation and other abnormal bleeding from female genital tract
C0156407|T047|HT|627|ICD9CM|Menopausal and postmenopausal disorders|Menopausal and postmenopausal disorders
C0156408|T046|PT|627.0|ICD9CM|Premenopausal menorrhagia|Premenopausal menorrhagia
C0156408|T046|AB|627.0|ICD9CM|Premenopause menorrhagia|Premenopause menorrhagia
C0032776|T046|AB|627.1|ICD9CM|Postmenopausal bleeding|Postmenopausal bleeding
C0032776|T046|PT|627.1|ICD9CM|Postmenopausal bleeding|Postmenopausal bleeding
C1135336|T047|AB|627.2|ICD9CM|Sympt fem climact state|Sympt fem climact state
C1135336|T047|PT|627.2|ICD9CM|Symptomatic menopausal or female climacteric states|Symptomatic menopausal or female climacteric states
C0156409|T047|AB|627.3|ICD9CM|Atrophic vaginitis|Atrophic vaginitis
C0156409|T047|PT|627.3|ICD9CM|Postmenopausal atrophic vaginitis|Postmenopausal atrophic vaginitis
C1135337|T047|AB|627.4|ICD9CM|Sympt state w artif meno|Sympt state w artif meno
C1135337|T047|PT|627.4|ICD9CM|Symptomatic states associated with artificial menopause|Symptomatic states associated with artificial menopause
C0156411|T047|AB|627.8|ICD9CM|Menopausal disorder NEC|Menopausal disorder NEC
C0156411|T047|PT|627.8|ICD9CM|Other specified menopausal and postmenopausal disorders|Other specified menopausal and postmenopausal disorders
C0156407|T047|AB|627.9|ICD9CM|Menopausal disorder NOS|Menopausal disorder NOS
C0156407|T047|PT|627.9|ICD9CM|Unspecified menopausal and postmenopausal disorder|Unspecified menopausal and postmenopausal disorder
C0021361|T046|HT|628|ICD9CM|Infertility, female|Infertility, female
C0404572|T047|AB|628.0|ICD9CM|Infertility-anovulation|Infertility-anovulation
C0404572|T047|PT|628.0|ICD9CM|Infertility, female, associated with anovulation|Infertility, female, associated with anovulation
C0156414|T047|AB|628.1|ICD9CM|Infertil-pituitary orig|Infertil-pituitary orig
C0156414|T047|PT|628.1|ICD9CM|Infertility, female, of pituitary-hypothalamic origin|Infertility, female, of pituitary-hypothalamic origin
C0156415|T047|AB|628.2|ICD9CM|Infertility-tubal origin|Infertility-tubal origin
C0156415|T047|PT|628.2|ICD9CM|Infertility, female, of tubal origin|Infertility, female, of tubal origin
C0156416|T046|AB|628.3|ICD9CM|Infertility-uterine orig|Infertility-uterine orig
C0156416|T046|PT|628.3|ICD9CM|Infertility, female, of uterine origin|Infertility, female, of uterine origin
C0156417|T047|AB|628.4|ICD9CM|Infertil-cervical orig|Infertil-cervical orig
C0156417|T047|PT|628.4|ICD9CM|Infertility, female, of cervical or vaginal origin|Infertility, female, of cervical or vaginal origin
C0021362|T033|AB|628.8|ICD9CM|Female infertility NEC|Female infertility NEC
C0021362|T033|PT|628.8|ICD9CM|Infertility, female, of other specified origin|Infertility, female, of other specified origin
C0021361|T046|AB|628.9|ICD9CM|Female infertility NOS|Female infertility NOS
C0021361|T046|PT|628.9|ICD9CM|Infertility, female, of unspecified origin|Infertility, female, of unspecified origin
C0156418|T047|HT|629|ICD9CM|Other disorders of female genital organs|Other disorders of female genital organs
C0869280|T047|AB|629.0|ICD9CM|Hematocele, female NEC|Hematocele, female NEC
C0869280|T047|PT|629.0|ICD9CM|Hematocele, female, not elsewhere classified|Hematocele, female, not elsewhere classified
C0156420|T190|AB|629.1|ICD9CM|Hydrocele canal nuck-fem|Hydrocele canal nuck-fem
C0156420|T190|PT|629.1|ICD9CM|Hydrocele, canal of nuck|Hydrocele, canal of nuck
C0744374|T033|HT|629.2|ICD9CM|Female genital mutilation status|Female genital mutilation status
C0744374|T033|PT|629.20|ICD9CM|Female genital mutilation status, unspecified|Female genital mutilation status, unspecified
C0744374|T033|AB|629.20|ICD9CM|Genital mutilation NOS|Genital mutilation NOS
C1456059|T047|PT|629.21|ICD9CM|Female genital mutilation Type I status|Female genital mutilation Type I status
C1456059|T047|AB|629.21|ICD9CM|Genital mutilatn type I|Genital mutilatn type I
C1456061|T047|PT|629.22|ICD9CM|Female genital mutilation Type II status|Female genital mutilation Type II status
C1456061|T047|AB|629.22|ICD9CM|Genital mutilatn type II|Genital mutilatn type II
C1456063|T047|PT|629.23|ICD9CM|Female genital mutilation Type III status|Female genital mutilation Type III status
C1456063|T047|AB|629.23|ICD9CM|Genital muilatn type III|Genital muilatn type III
C1719551|T033|AB|629.29|ICD9CM|Fem genital mutilate NEC|Fem genital mutilate NEC
C1719551|T033|PT|629.29|ICD9CM|Other female genital mutilation status|Other female genital mutilation status
C3161257|T046|HT|629.3|ICD9CM|Complication of implanted vaginal mesh and other prosthetic materials|Complication of implanted vaginal mesh and other prosthetic materials
C3161118|T046|AB|629.31|ICD9CM|Eros imp vag mesh in tis|Eros imp vag mesh in tis
C3161118|T046|PT|629.31|ICD9CM|Erosion of implanted vaginal mesh and other prosthetic materials to surrounding organ or tissue|Erosion of implanted vaginal mesh and other prosthetic materials to surrounding organ or tissue
C3161119|T046|AB|629.32|ICD9CM|Exp imp vag mesh-vagina|Exp imp vag mesh-vagina
C3161119|T046|PT|629.32|ICD9CM|Exposure of implanted vaginal mesh and other prosthetic materials into vagina|Exposure of implanted vaginal mesh and other prosthetic materials into vagina
C0156421|T047|HT|629.8|ICD9CM|Other specified disorders of female genital organs|Other specified disorders of female genital organs
C2921105|T046|AB|629.81|ICD9CM|Rec preg loss wo cur prg|Rec preg loss wo cur prg
C2921105|T046|PT|629.81|ICD9CM|Recurrent pregnancy loss without current pregnancy|Recurrent pregnancy loss without current pregnancy
C0156421|T047|AB|629.89|ICD9CM|Female genital disor NEC|Female genital disor NEC
C0156421|T047|PT|629.89|ICD9CM|Other specified disorders of female genital organs|Other specified disorders of female genital organs
C0017411|T047|AB|629.9|ICD9CM|Female genital dis NOS|Female genital dis NOS
C0017411|T047|PT|629.9|ICD9CM|Unspecified disorder of female genital organs|Unspecified disorder of female genital organs
C0020217|T191|AB|630|ICD9CM|Hydatidiform mole|Hydatidiform mole
C0020217|T191|PT|630|ICD9CM|Hydatidiform mole|Hydatidiform mole
C0178293|T047|HT|630-633.99|ICD9CM|ECTOPIC AND MOLAR PREGNANCY|ECTOPIC AND MOLAR PREGNANCY
C0178292|T046|HT|630-679.99|ICD9CM|COMPLICATIONS OF PREGNANCY, CHILDBIRTH, AND THE PUERPERIUM|COMPLICATIONS OF PREGNANCY, CHILDBIRTH, AND THE PUERPERIUM
C0156422|T047|HT|631|ICD9CM|Other abnormal product of conception|Other abnormal product of conception
C3161120|T033|AB|631.0|ICD9CM|Inapp chg hCG early preg|Inapp chg hCG early preg
C3161120|T033|PT|631.0|ICD9CM|Inappropriate change in quantitative human chorionic gonadotropin (hCG) in early pregnancy|Inappropriate change in quantitative human chorionic gonadotropin (hCG) in early pregnancy
C0156422|T047|AB|631.8|ICD9CM|Oth abn prod conception|Oth abn prod conception
C0156422|T047|PT|631.8|ICD9CM|Other abnormal products of conception|Other abnormal products of conception
C0000814|T047|AB|632|ICD9CM|Missed abortion|Missed abortion
C0000814|T047|PT|632|ICD9CM|Missed abortion|Missed abortion
C0032987|T046|HT|633|ICD9CM|Ectopic pregnancy|Ectopic pregnancy
C0032984|T046|HT|633.0|ICD9CM|Abdominal pregnancy|Abdominal pregnancy
C1135231|T046|AB|633.00|ICD9CM|Abd preg w/o intrau preg|Abd preg w/o intrau preg
C1135231|T046|PT|633.00|ICD9CM|Abdominal pregnancy without intrauterine pregnancy|Abdominal pregnancy without intrauterine pregnancy
C1135232|T046|AB|633.01|ICD9CM|Abd preg w intraut preg|Abd preg w intraut preg
C1135232|T046|PT|633.01|ICD9CM|Abdominal pregnancy with intrauterine pregnancy|Abdominal pregnancy with intrauterine pregnancy
C0032994|T046|HT|633.1|ICD9CM|Tubal pregnancy|Tubal pregnancy
C1135233|T046|AB|633.10|ICD9CM|Tubal preg w/o intra prg|Tubal preg w/o intra prg
C1135233|T046|PT|633.10|ICD9CM|Tubal pregnancy without intrauterine pregnancy|Tubal pregnancy without intrauterine pregnancy
C1135234|T046|AB|633.11|ICD9CM|Tubal preg w intra preg|Tubal preg w intra preg
C1135234|T046|PT|633.11|ICD9CM|Tubal pregnancy with intrauterine pregnancy|Tubal pregnancy with intrauterine pregnancy
C0032991|T046|HT|633.2|ICD9CM|Ovarian pregnancy|Ovarian pregnancy
C1135235|T046|PT|633.20|ICD9CM|Ovarian pregnancy without intrauterine pregnancy|Ovarian pregnancy without intrauterine pregnancy
C1135235|T046|AB|633.20|ICD9CM|Ovarn preg w/o intra prg|Ovarn preg w/o intra prg
C1135236|T046|AB|633.21|ICD9CM|Ovarian preg w intra prg|Ovarian preg w intra prg
C1135236|T046|PT|633.21|ICD9CM|Ovarian pregnancy with intrauterine pregnancy|Ovarian pregnancy with intrauterine pregnancy
C0029604|T046|HT|633.8|ICD9CM|Other ectopic pregnancy|Other ectopic pregnancy
C1135237|T047|AB|633.80|ICD9CM|Ect preg NEC w/o int prg|Ect preg NEC w/o int prg
C1135237|T047|PT|633.80|ICD9CM|Other ectopic pregnancy without intrauterine pregnancy|Other ectopic pregnancy without intrauterine pregnancy
C1135238|T047|AB|633.81|ICD9CM|Ectpc prg NEC w int preg|Ectpc prg NEC w int preg
C1135238|T047|PT|633.81|ICD9CM|Other ectopic pregnancy with intrauterine pregnancy|Other ectopic pregnancy with intrauterine pregnancy
C0032987|T046|HT|633.9|ICD9CM|Unspecified ectopic pregnancy|Unspecified ectopic pregnancy
C1135239|T046|AB|633.90|ICD9CM|Ect preg NOS w/o int prg|Ect preg NOS w/o int prg
C1135239|T046|PT|633.90|ICD9CM|Unspecified ectopic pregnancy without intrauterine pregnancy|Unspecified ectopic pregnancy without intrauterine pregnancy
C1135240|T046|AB|633.91|ICD9CM|Ectp preg NOS w int preg|Ectp preg NOS w int preg
C1135240|T046|PT|633.91|ICD9CM|Unspecified ectopic pregnancy with intrauterine pregnancy|Unspecified ectopic pregnancy with intrauterine pregnancy
C0000786|T046|HT|634|ICD9CM|Spontaneous abortion|Spontaneous abortion
C0178294|T047|HT|634-639.99|ICD9CM|OTHER PREGNANCY WITH ABORTIVE OUTCOME|OTHER PREGNANCY WITH ABORTIVE OUTCOME
C0156424|T047|HT|634.0|ICD9CM|Spontaneous abortion complicated by genital tract and pelvic infection|Spontaneous abortion complicated by genital tract and pelvic infection
C0156424|T047|AB|634.00|ICD9CM|Spon abor w pel inf-unsp|Spon abor w pel inf-unsp
C0156424|T047|PT|634.00|ICD9CM|Spontaneous abortion, complicated by genital tract and pelvic infection, unspecified|Spontaneous abortion, complicated by genital tract and pelvic infection, unspecified
C0156425|T047|AB|634.01|ICD9CM|Spon abor w pelv inf-inc|Spon abor w pelv inf-inc
C0156425|T047|PT|634.01|ICD9CM|Spontaneous abortion, complicated by genital tract and pelvic infection, incomplete|Spontaneous abortion, complicated by genital tract and pelvic infection, incomplete
C0156426|T047|AB|634.02|ICD9CM|Spon abor w pel inf-comp|Spon abor w pel inf-comp
C0156426|T047|PT|634.02|ICD9CM|Spontaneous abortion, complicated by genital tract and pelvic infection, complete|Spontaneous abortion, complicated by genital tract and pelvic infection, complete
C0156427|T046|HT|634.1|ICD9CM|Spontaneous abortion complicated by delayed or excessive hemorrhage|Spontaneous abortion complicated by delayed or excessive hemorrhage
C0156428|T047|AB|634.10|ICD9CM|Spon abort w hemorr-unsp|Spon abort w hemorr-unsp
C0156428|T047|PT|634.10|ICD9CM|Spontaneous abortion, complicated by delayed or excessive hemorrhage, unspecified|Spontaneous abortion, complicated by delayed or excessive hemorrhage, unspecified
C0156429|T046|AB|634.11|ICD9CM|Spon abort w hemorr-inc|Spon abort w hemorr-inc
C0156429|T046|PT|634.11|ICD9CM|Spontaneous abortion, complicated by delayed or excessive hemorrhage, incomplete|Spontaneous abortion, complicated by delayed or excessive hemorrhage, incomplete
C0156430|T047|AB|634.12|ICD9CM|Spon abort w hemorr-comp|Spon abort w hemorr-comp
C0156430|T047|PT|634.12|ICD9CM|Spontaneous abortion, complicated by delayed or excessive hemorrhage, complete|Spontaneous abortion, complicated by delayed or excessive hemorrhage, complete
C0269403|T047|HT|634.2|ICD9CM|Spontaneous abortion complicated by damage to pelvic organs or tissues|Spontaneous abortion complicated by damage to pelvic organs or tissues
C0269403|T047|AB|634.20|ICD9CM|Spon ab w pel damag-unsp|Spon ab w pel damag-unsp
C0269403|T047|PT|634.20|ICD9CM|Spontaneous abortion, complicated by damage to pelvic organs or tissues, unspecified|Spontaneous abortion, complicated by damage to pelvic organs or tissues, unspecified
C0156433|T037|AB|634.21|ICD9CM|Spon ab w pelv damag-inc|Spon ab w pelv damag-inc
C0156433|T037|PT|634.21|ICD9CM|Spontaneous abortion, complicated by damage to pelvic organs or tissues, incomplete|Spontaneous abortion, complicated by damage to pelvic organs or tissues, incomplete
C0156434|T037|AB|634.22|ICD9CM|Spon ab w pel damag-comp|Spon ab w pel damag-comp
C0156434|T037|PT|634.22|ICD9CM|Spontaneous abortion, complicated by damage to pelvic organs or tissues, complete|Spontaneous abortion, complicated by damage to pelvic organs or tissues, complete
C0156435|T047|HT|634.3|ICD9CM|Spontaneous abortion complicated by renal failure|Spontaneous abortion complicated by renal failure
C0156436|T047|AB|634.30|ICD9CM|Spon ab w ren fail-unsp|Spon ab w ren fail-unsp
C0156436|T047|PT|634.30|ICD9CM|Spontaneous abortion, complicated by renal failure, unspecified|Spontaneous abortion, complicated by renal failure, unspecified
C0404922|T047|AB|634.31|ICD9CM|Spon ab w ren fail-inc|Spon ab w ren fail-inc
C0404922|T047|PT|634.31|ICD9CM|Spontaneous abortion, complicated by renal failure, incomplete|Spontaneous abortion, complicated by renal failure, incomplete
C0404905|T046|AB|634.32|ICD9CM|Spon ab w ren fail-comp|Spon ab w ren fail-comp
C0404905|T046|PT|634.32|ICD9CM|Spontaneous abortion, complicated by renal failure, complete|Spontaneous abortion, complicated by renal failure, complete
C0156439|T047|HT|634.4|ICD9CM|Spontaneous abortion complicated by metabolic disorder|Spontaneous abortion complicated by metabolic disorder
C0156439|T047|AB|634.40|ICD9CM|Spon ab w metab dis-unsp|Spon ab w metab dis-unsp
C0156439|T047|PT|634.40|ICD9CM|Spontaneous abortion, complicated by metabolic disorder, unspecified|Spontaneous abortion, complicated by metabolic disorder, unspecified
C0404921|T046|AB|634.41|ICD9CM|Spon ab w metab dis-inc|Spon ab w metab dis-inc
C0404921|T046|PT|634.41|ICD9CM|Spontaneous abortion, complicated by metabolic disorder, incomplete|Spontaneous abortion, complicated by metabolic disorder, incomplete
C0156442|T047|AB|634.42|ICD9CM|Spon ab w metab dis-comp|Spon ab w metab dis-comp
C0156442|T047|PT|634.42|ICD9CM|Spontaneous abortion, complicated by metabolic disorder, complete|Spontaneous abortion, complicated by metabolic disorder, complete
C0156443|T047|HT|634.5|ICD9CM|Spontaneous abortion complicated by shock|Spontaneous abortion complicated by shock
C0156444|T047|AB|634.50|ICD9CM|Spon abort w shock-unsp|Spon abort w shock-unsp
C0156444|T047|PT|634.50|ICD9CM|Spontaneous abortion, complicated by shock, unspecified|Spontaneous abortion, complicated by shock, unspecified
C0156445|T047|AB|634.51|ICD9CM|Spon abort w shock-inc|Spon abort w shock-inc
C0156445|T047|PT|634.51|ICD9CM|Spontaneous abortion, complicated by shock, incomplete|Spontaneous abortion, complicated by shock, incomplete
C0404903|T046|AB|634.52|ICD9CM|Spon abort w shock-comp|Spon abort w shock-comp
C0404903|T046|PT|634.52|ICD9CM|Spontaneous abortion, complicated by shock, complete|Spontaneous abortion, complicated by shock, complete
C0156447|T047|HT|634.6|ICD9CM|Spontaneous abortion complicated by embolism|Spontaneous abortion complicated by embolism
C0156448|T047|AB|634.60|ICD9CM|Spon abort w embol-unsp|Spon abort w embol-unsp
C0156448|T047|PT|634.60|ICD9CM|Spontaneous abortion, complicated by embolism, unspecified|Spontaneous abortion, complicated by embolism, unspecified
C0404919|T046|AB|634.61|ICD9CM|Spon abort w embol-inc|Spon abort w embol-inc
C0404919|T046|PT|634.61|ICD9CM|Spontaneous abortion, complicated by embolism, incomplete|Spontaneous abortion, complicated by embolism, incomplete
C0404902|T046|AB|634.62|ICD9CM|Spon abort w embol-comp|Spon abort w embol-comp
C0404902|T046|PT|634.62|ICD9CM|Spontaneous abortion, complicated by embolism, complete|Spontaneous abortion, complicated by embolism, complete
C0156452|T047|HT|634.7|ICD9CM|Spontaneous abortion with other specified complications|Spontaneous abortion with other specified complications
C0156452|T047|AB|634.70|ICD9CM|Spon ab w compl NEC-unsp|Spon ab w compl NEC-unsp
C0156452|T047|PT|634.70|ICD9CM|Spontaneous abortion, with other specified complications, unspecified|Spontaneous abortion, with other specified complications, unspecified
C0156453|T047|AB|634.71|ICD9CM|Spon ab w compl NEC-inc|Spon ab w compl NEC-inc
C0156453|T047|PT|634.71|ICD9CM|Spontaneous abortion, with other specified complications, incomplete|Spontaneous abortion, with other specified complications, incomplete
C0156454|T047|AB|634.72|ICD9CM|Spon ab w compl NEC-comp|Spon ab w compl NEC-comp
C0156454|T047|PT|634.72|ICD9CM|Spontaneous abortion, with other specified complications, complete|Spontaneous abortion, with other specified complications, complete
C0156456|T046|HT|634.8|ICD9CM|Spontaneous abortion with unspecified complication|Spontaneous abortion with unspecified complication
C0156456|T046|AB|634.80|ICD9CM|Spon ab w compl NOS-unsp|Spon ab w compl NOS-unsp
C0156456|T046|PT|634.80|ICD9CM|Spontaneous abortion, with unspecified complication, unspecified|Spontaneous abortion, with unspecified complication, unspecified
C0156457|T046|AB|634.81|ICD9CM|Spon ab w compl NOS-inc|Spon ab w compl NOS-inc
C0156457|T046|PT|634.81|ICD9CM|Spontaneous abortion, with unspecified complication, incomplete|Spontaneous abortion, with unspecified complication, incomplete
C0156458|T047|AB|634.82|ICD9CM|Spon ab w compl NOS-comp|Spon ab w compl NOS-comp
C0156458|T047|PT|634.82|ICD9CM|Spontaneous abortion, with unspecified complication, complete|Spontaneous abortion, with unspecified complication, complete
C0156459|T046|HT|634.9|ICD9CM|Spontaneous abortion without mention of complication|Spontaneous abortion without mention of complication
C0156459|T046|AB|634.90|ICD9CM|Spon abort uncompl-unsp|Spon abort uncompl-unsp
C0156459|T046|PT|634.90|ICD9CM|Spontaneous abortion, without mention of complication, unspecified|Spontaneous abortion, without mention of complication, unspecified
C0729205|T046|AB|634.91|ICD9CM|Spon abort uncompl-inc|Spon abort uncompl-inc
C0729205|T046|PT|634.91|ICD9CM|Spontaneous abortion, without mention of complication, incomplete|Spontaneous abortion, without mention of complication, incomplete
C0156461|T047|AB|634.92|ICD9CM|Spon abort uncompl-comp|Spon abort uncompl-comp
C0156461|T047|PT|634.92|ICD9CM|Spontaneous abortion, without mention of complication, complete|Spontaneous abortion, without mention of complication, complete
C1456876|T033|HT|635|ICD9CM|Legally induced abortion|Legally induced abortion
C0156464|T047|HT|635.0|ICD9CM|Legally induced abortion complicated by genital tract and pelvic infection|Legally induced abortion complicated by genital tract and pelvic infection
C0156464|T047|AB|635.00|ICD9CM|Leg abor w pelv inf-unsp|Leg abor w pelv inf-unsp
C0156464|T047|PT|635.00|ICD9CM|Legally induced abortion, complicated by genital tract and pelvic infection, unspecified|Legally induced abortion, complicated by genital tract and pelvic infection, unspecified
C0156465|T046|AB|635.01|ICD9CM|Leg abor w pelv inf-inc|Leg abor w pelv inf-inc
C0156465|T046|PT|635.01|ICD9CM|Legally induced abortion, complicated by genital tract and pelvic infection, incomplete|Legally induced abortion, complicated by genital tract and pelvic infection, incomplete
C0156466|T046|AB|635.02|ICD9CM|Leg abor w pelv inf-comp|Leg abor w pelv inf-comp
C0156466|T046|PT|635.02|ICD9CM|Legally induced abortion, complicated by genital tract and pelvic infection, complete|Legally induced abortion, complicated by genital tract and pelvic infection, complete
C0269450|T046|HT|635.1|ICD9CM|Legally induced abortion complicated by delayed or excessive hemorrhage|Legally induced abortion complicated by delayed or excessive hemorrhage
C0269450|T046|AB|635.10|ICD9CM|Legal abor w hemorr-unsp|Legal abor w hemorr-unsp
C0269450|T046|PT|635.10|ICD9CM|Legally induced abortion, complicated by delayed or excessive hemorrhage, unspecified|Legally induced abortion, complicated by delayed or excessive hemorrhage, unspecified
C0156469|T046|AB|635.11|ICD9CM|Legal abort w hemorr-inc|Legal abort w hemorr-inc
C0156469|T046|PT|635.11|ICD9CM|Legally induced abortion, complicated by delayed or excessive hemorrhage, incomplete|Legally induced abortion, complicated by delayed or excessive hemorrhage, incomplete
C0156470|T046|AB|635.12|ICD9CM|Legal abor w hemorr-comp|Legal abor w hemorr-comp
C0156470|T046|PT|635.12|ICD9CM|Legally induced abortion, complicated by delayed or excessive hemorrhage, complete|Legally induced abortion, complicated by delayed or excessive hemorrhage, complete
C0156472|T046|HT|635.2|ICD9CM|Legally induced abortion complicated by damage to pelvic organs or tissues|Legally induced abortion complicated by damage to pelvic organs or tissues
C0156472|T046|AB|635.20|ICD9CM|Leg ab w pelv damag-unsp|Leg ab w pelv damag-unsp
C0156472|T046|PT|635.20|ICD9CM|Legally induced abortion, complicated by damage to pelvic organs or tissues, unspecified|Legally induced abortion, complicated by damage to pelvic organs or tissues, unspecified
C0156473|T046|AB|635.21|ICD9CM|Leg ab w pelv damag-inc|Leg ab w pelv damag-inc
C0156473|T046|PT|635.21|ICD9CM|Legally induced abortion, complicated by damage to pelvic organs or tissues, incomplete|Legally induced abortion, complicated by damage to pelvic organs or tissues, incomplete
C0156474|T037|AB|635.22|ICD9CM|Leg ab w pelv damag-comp|Leg ab w pelv damag-comp
C0156474|T037|PT|635.22|ICD9CM|Legally induced abortion, complicated by damage to pelvic organs or tissues, complete|Legally induced abortion, complicated by damage to pelvic organs or tissues, complete
C0269469|T046|HT|635.3|ICD9CM|Legally induced abortion complicated by renal failure|Legally induced abortion complicated by renal failure
C0269469|T046|AB|635.30|ICD9CM|Leg abor w ren fail-unsp|Leg abor w ren fail-unsp
C0269469|T046|PT|635.30|ICD9CM|Legally induced abortion, complicated by renal failure,unspecified|Legally induced abortion, complicated by renal failure,unspecified
C0156477|T046|AB|635.31|ICD9CM|Leg abor w ren fail-inc|Leg abor w ren fail-inc
C0156477|T046|PT|635.31|ICD9CM|Legally induced abortion, complicated by renal failure, incomplete|Legally induced abortion, complicated by renal failure, incomplete
C0156478|T046|AB|635.32|ICD9CM|Leg abor w ren fail-comp|Leg abor w ren fail-comp
C0156478|T046|PT|635.32|ICD9CM|Legally induced abortion, complicated by renal failure, complete|Legally induced abortion, complicated by renal failure, complete
C0269474|T046|HT|635.4|ICD9CM|Legally induced abortion complicated by metabolic disorder|Legally induced abortion complicated by metabolic disorder
C0269474|T046|AB|635.40|ICD9CM|Leg ab w metab dis-unsp|Leg ab w metab dis-unsp
C0269474|T046|PT|635.40|ICD9CM|Legally induced abortion, complicated by metabolic disorder, unspecified|Legally induced abortion, complicated by metabolic disorder, unspecified
C0156481|T046|AB|635.41|ICD9CM|Leg ab w metab dis-inc|Leg ab w metab dis-inc
C0156481|T046|PT|635.41|ICD9CM|Legally induced abortion, complicated by metabolic disorder, incomplete|Legally induced abortion, complicated by metabolic disorder, incomplete
C0156482|T046|AB|635.42|ICD9CM|Leg ab w metab dis-comp|Leg ab w metab dis-comp
C0156482|T046|PT|635.42|ICD9CM|Legally induced abortion, complicated by metabolic disorder, complete|Legally induced abortion, complicated by metabolic disorder, complete
C0269476|T046|HT|635.5|ICD9CM|Legally induced abortion complicated by shock|Legally induced abortion complicated by shock
C0269476|T046|AB|635.50|ICD9CM|Legal abort w shock-unsp|Legal abort w shock-unsp
C0269476|T046|PT|635.50|ICD9CM|Legally induced abortion, complicated by shock, unspecified|Legally induced abortion, complicated by shock, unspecified
C0156485|T046|AB|635.51|ICD9CM|Legal abort w shock-inc|Legal abort w shock-inc
C0156485|T046|PT|635.51|ICD9CM|Legally induced abortion, complicated by shock, incomplete|Legally induced abortion, complicated by shock, incomplete
C0156486|T046|AB|635.52|ICD9CM|Legal abort w shock-comp|Legal abort w shock-comp
C0156486|T046|PT|635.52|ICD9CM|Legally induced abortion, complicated by shock, complete|Legally induced abortion, complicated by shock, complete
C0269479|T046|HT|635.6|ICD9CM|Legally induced abortion complicated by embolism|Legally induced abortion complicated by embolism
C0269479|T046|AB|635.60|ICD9CM|Legal abort w embol-unsp|Legal abort w embol-unsp
C0269479|T046|PT|635.60|ICD9CM|Legally induced abortion, complicated by embolism, unspecified|Legally induced abortion, complicated by embolism, unspecified
C0156489|T046|AB|635.61|ICD9CM|Legal abort w embol-inc|Legal abort w embol-inc
C0156489|T046|PT|635.61|ICD9CM|Legally induced abortion, complicated by embolism, incomplete|Legally induced abortion, complicated by embolism, incomplete
C0156490|T046|AB|635.62|ICD9CM|Legal abort w embol-comp|Legal abort w embol-comp
C0156490|T046|PT|635.62|ICD9CM|Legally induced abortion, complicated by embolism, complete|Legally induced abortion, complicated by embolism, complete
C0156492|T046|HT|635.7|ICD9CM|Legally induced abortion with other specified complications|Legally induced abortion with other specified complications
C0156492|T046|AB|635.70|ICD9CM|Leg ab w compl NEC-unsp|Leg ab w compl NEC-unsp
C0156492|T046|PT|635.70|ICD9CM|Legally induced abortion, with other specified complications, unspecified|Legally induced abortion, with other specified complications, unspecified
C0156493|T046|AB|635.71|ICD9CM|Leg ab w compl NEC-inc|Leg ab w compl NEC-inc
C0156493|T046|PT|635.71|ICD9CM|Legally induced abortion, with other specified complications, incomplete|Legally induced abortion, with other specified complications, incomplete
C0156494|T046|AB|635.72|ICD9CM|Leg ab w compl NEC-comp|Leg ab w compl NEC-comp
C0156494|T046|PT|635.72|ICD9CM|Legally induced abortion, with other specified complications, complete|Legally induced abortion, with other specified complications, complete
C0269441|T046|HT|635.8|ICD9CM|Legally induced abortion with unspecified complication|Legally induced abortion with unspecified complication
C0269441|T046|AB|635.80|ICD9CM|Leg ab w compl NOS-unsp|Leg ab w compl NOS-unsp
C0269441|T046|PT|635.80|ICD9CM|Legally induced abortion, with unspecified complication, unspecified|Legally induced abortion, with unspecified complication, unspecified
C0600042|T046|AB|635.81|ICD9CM|Leg ab w compl NOS-inc|Leg ab w compl NOS-inc
C0600042|T046|PT|635.81|ICD9CM|Legally induced abortion, with unspecified complication, incomplete|Legally induced abortion, with unspecified complication, incomplete
C0156498|T046|AB|635.82|ICD9CM|Leg ab w compl NOS-comp|Leg ab w compl NOS-comp
C0156498|T046|PT|635.82|ICD9CM|Legally induced abortion, with unspecified complication, complete|Legally induced abortion, with unspecified complication, complete
C0156499|T033|HT|635.9|ICD9CM|Legally induced abortion without mention of complication|Legally induced abortion without mention of complication
C0156499|T033|AB|635.90|ICD9CM|Legal abort uncompl-unsp|Legal abort uncompl-unsp
C0156499|T033|PT|635.90|ICD9CM|Legally induced abortion, without mention of complication, unspecified|Legally induced abortion, without mention of complication, unspecified
C0600043|T046|AB|635.91|ICD9CM|Legal abort uncompl-inc|Legal abort uncompl-inc
C0600043|T046|PT|635.91|ICD9CM|Legally induced abortion, without mention of complication, incomplete|Legally induced abortion, without mention of complication, incomplete
C1261319|T047|AB|635.92|ICD9CM|Legal abort uncompl-comp|Legal abort uncompl-comp
C1261319|T047|PT|635.92|ICD9CM|Legally induced abortion, without mention of complication, complete|Legally induced abortion, without mention of complication, complete
C0000804|T033|HT|636|ICD9CM|Illegally induced abortion|Illegally induced abortion
C0156504|T046|HT|636.0|ICD9CM|Illegally induced abortion complicated by genital tract and pelvic infection|Illegally induced abortion complicated by genital tract and pelvic infection
C0156504|T046|AB|636.00|ICD9CM|Illeg ab w pelv inf-unsp|Illeg ab w pelv inf-unsp
C0156504|T046|PT|636.00|ICD9CM|Illegally induced abortion, complicated by genital tract and pelvic infection, unspecified|Illegally induced abortion, complicated by genital tract and pelvic infection, unspecified
C0156505|T046|AB|636.01|ICD9CM|Illeg ab w pelv inf-inc|Illeg ab w pelv inf-inc
C0156505|T046|PT|636.01|ICD9CM|Illegally induced abortion, complicated by genital tract and pelvic infection, incomplete|Illegally induced abortion, complicated by genital tract and pelvic infection, incomplete
C0156506|T037|AB|636.02|ICD9CM|Illeg ab w pelv inf-comp|Illeg ab w pelv inf-comp
C0156506|T037|PT|636.02|ICD9CM|Illegally induced abortion, complicated by genital tract and pelvic infection, complete|Illegally induced abortion, complicated by genital tract and pelvic infection, complete
C0269505|T033|HT|636.1|ICD9CM|Illegally induced abortion complicated by delayed or excessive hemorrhage|Illegally induced abortion complicated by delayed or excessive hemorrhage
C0269505|T033|AB|636.10|ICD9CM|Illeg ab w hemorr-unspec|Illeg ab w hemorr-unspec
C0269505|T033|PT|636.10|ICD9CM|Illegally induced abortion, complicated by delayed or excessive hemorrhage, unspecified|Illegally induced abortion, complicated by delayed or excessive hemorrhage, unspecified
C0156509|T047|AB|636.11|ICD9CM|Illeg ab w hemorr-inc|Illeg ab w hemorr-inc
C0156509|T047|PT|636.11|ICD9CM|Illegally induced abortion, complicated by delayed or excessive hemorrhage, incomplete|Illegally induced abortion, complicated by delayed or excessive hemorrhage, incomplete
C0156510|T047|AB|636.12|ICD9CM|Illeg ab w hemorr-comp|Illeg ab w hemorr-comp
C0156510|T047|PT|636.12|ICD9CM|Illegally induced abortion, complicated by delayed or excessive hemorrhage, complete|Illegally induced abortion, complicated by delayed or excessive hemorrhage, complete
C0269509|T046|HT|636.2|ICD9CM|Illegally induced abortion complicated by damage to pelvic organs or tissue|Illegally induced abortion complicated by damage to pelvic organs or tissue
C0269509|T046|AB|636.20|ICD9CM|Illeg ab w pel damg-unsp|Illeg ab w pel damg-unsp
C0269509|T046|PT|636.20|ICD9CM|Illegally induced abortion, complicated by damage to pelvic organs or tissues, unspecified|Illegally induced abortion, complicated by damage to pelvic organs or tissues, unspecified
C0156513|T037|AB|636.21|ICD9CM|Illeg ab w pel damag-inc|Illeg ab w pel damag-inc
C0156513|T037|PT|636.21|ICD9CM|Illegally induced abortion, complicated by damage to pelvic organs or tissues, incomplete|Illegally induced abortion, complicated by damage to pelvic organs or tissues, incomplete
C0156514|T037|AB|636.22|ICD9CM|Illeg ab w pel damg-comp|Illeg ab w pel damg-comp
C0156514|T037|PT|636.22|ICD9CM|Illegally induced abortion, complicated by damage to pelvic organs or tissues, complete|Illegally induced abortion, complicated by damage to pelvic organs or tissues, complete
C0269524|T046|HT|636.3|ICD9CM|Illegally induced abortion complicated by renal failure|Illegally induced abortion complicated by renal failure
C0269524|T046|AB|636.30|ICD9CM|Illeg ab w ren fail-unsp|Illeg ab w ren fail-unsp
C0269524|T046|PT|636.30|ICD9CM|Illegally induced abortion, complicated by renal failure, unspecified|Illegally induced abortion, complicated by renal failure, unspecified
C0156517|T047|AB|636.31|ICD9CM|Illeg ab w ren fail-inc|Illeg ab w ren fail-inc
C0156517|T047|PT|636.31|ICD9CM|Illegally induced abortion, complicated by renal failure, incomplete|Illegally induced abortion, complicated by renal failure, incomplete
C0156518|T047|AB|636.32|ICD9CM|Illeg ab w ren fail-comp|Illeg ab w ren fail-comp
C0156518|T047|PT|636.32|ICD9CM|Illegally induced abortion, complicated by renal failure, complete|Illegally induced abortion, complicated by renal failure, complete
C0269529|T046|HT|636.4|ICD9CM|Illegally induced abortion complicated by metabolic disorder|Illegally induced abortion complicated by metabolic disorder
C0269529|T046|AB|636.40|ICD9CM|Illeg ab w met dis-unsp|Illeg ab w met dis-unsp
C0269529|T046|PT|636.40|ICD9CM|Illegally induced abortion, complicated by metabolic disorder, unspecified|Illegally induced abortion, complicated by metabolic disorder, unspecified
C0156521|T047|AB|636.41|ICD9CM|Illeg ab w metab dis-inc|Illeg ab w metab dis-inc
C0156521|T047|PT|636.41|ICD9CM|Illegally induced abortion, complicated by metabolic disorder, incomplete|Illegally induced abortion, complicated by metabolic disorder, incomplete
C0156522|T047|AB|636.42|ICD9CM|Illeg ab w met dis-comp|Illeg ab w met dis-comp
C0156522|T047|PT|636.42|ICD9CM|Illegally induced abortion, complicated by metabolic disorder, complete|Illegally induced abortion, complicated by metabolic disorder, complete
C0269531|T046|HT|636.5|ICD9CM|Illegally induced abortion complicated by shock|Illegally induced abortion complicated by shock
C0269531|T046|AB|636.50|ICD9CM|Illeg abort w shock-unsp|Illeg abort w shock-unsp
C0269531|T046|PT|636.50|ICD9CM|Illegally induced abortion, complicated by shock, unspecified|Illegally induced abortion, complicated by shock, unspecified
C0156525|T037|AB|636.51|ICD9CM|Illeg abort w shock-inc|Illeg abort w shock-inc
C0156525|T037|PT|636.51|ICD9CM|Illegally induced abortion, complicated by shock, incomplete|Illegally induced abortion, complicated by shock, incomplete
C0156526|T037|AB|636.52|ICD9CM|Illeg abort w shock-comp|Illeg abort w shock-comp
C0156526|T037|PT|636.52|ICD9CM|Illegally induced abortion, complicated by shock, complete|Illegally induced abortion, complicated by shock, complete
C0269534|T046|HT|636.6|ICD9CM|Illegally induced abortion complicated by embolism|Illegally induced abortion complicated by embolism
C0269534|T046|AB|636.60|ICD9CM|Illeg ab w embolism-unsp|Illeg ab w embolism-unsp
C0269534|T046|PT|636.60|ICD9CM|Illegally induced abortion, complicated by embolism, unspecified|Illegally induced abortion, complicated by embolism, unspecified
C0156529|T037|AB|636.61|ICD9CM|Illeg ab w embolism-inc|Illeg ab w embolism-inc
C0156529|T037|PT|636.61|ICD9CM|Illegally induced abortion, complicated by embolism, incomplete|Illegally induced abortion, complicated by embolism, incomplete
C0156530|T037|AB|636.62|ICD9CM|Illeg ab w embolism-comp|Illeg ab w embolism-comp
C0156530|T037|PT|636.62|ICD9CM|Illegally induced abortion, complicated by embolism, complete|Illegally induced abortion, complicated by embolism, complete
C0156532|T046|HT|636.7|ICD9CM|Illegally induced abortion with other specified complications|Illegally induced abortion with other specified complications
C0156532|T046|PT|636.70|ICD9CM|Illegally induced abortion, with other specified complications, unspecified|Illegally induced abortion, with other specified complications, unspecified
C0156532|T046|AB|636.70|ICD9CM|Illg ab w compl NEC-unsp|Illg ab w compl NEC-unsp
C0156533|T046|AB|636.71|ICD9CM|Illeg ab w compl NEC-inc|Illeg ab w compl NEC-inc
C0156533|T046|PT|636.71|ICD9CM|Illegally induced abortion, with other specified complications, incomplete|Illegally induced abortion, with other specified complications, incomplete
C0156534|T046|PT|636.72|ICD9CM|Illegally induced abortion, with other specified complications, complete|Illegally induced abortion, with other specified complications, complete
C0156534|T046|AB|636.72|ICD9CM|Illg ab w compl NEC-comp|Illg ab w compl NEC-comp
C0269496|T046|HT|636.8|ICD9CM|Illegally induced abortion with unspecified complication|Illegally induced abortion with unspecified complication
C0269496|T046|PT|636.80|ICD9CM|Illegally induced abortion, with unspecified complication, unspecified|Illegally induced abortion, with unspecified complication, unspecified
C0269496|T046|AB|636.80|ICD9CM|Illg ab w compl NOS-unsp|Illg ab w compl NOS-unsp
C0156537|T037|AB|636.81|ICD9CM|Illeg ab w compl NOS-inc|Illeg ab w compl NOS-inc
C0156537|T037|PT|636.81|ICD9CM|Illegally induced abortion, with unspecified complication, incomplete|Illegally induced abortion, with unspecified complication, incomplete
C0156538|T037|PT|636.82|ICD9CM|Illegally induced abortion, with unspecified complication, complete|Illegally induced abortion, with unspecified complication, complete
C0156538|T037|AB|636.82|ICD9CM|Illg ab w compl NOS-comp|Illg ab w compl NOS-comp
C0260335|T046|HT|636.9|ICD9CM|Illegally induced abortion without mention of complication|Illegally induced abortion without mention of complication
C0260335|T046|AB|636.90|ICD9CM|Illeg abort uncompl-unsp|Illeg abort uncompl-unsp
C0260335|T046|PT|636.90|ICD9CM|Illegally induced abortion, without mention of complication, unspecified|Illegally induced abortion, without mention of complication, unspecified
C0156541|T037|AB|636.91|ICD9CM|Illeg abort uncompl-inc|Illeg abort uncompl-inc
C0156541|T037|PT|636.91|ICD9CM|Illegally induced abortion, without mention of complication, incomplete|Illegally induced abortion, without mention of complication, incomplete
C0156542|T046|AB|636.92|ICD9CM|Illeg abort uncompl-comp|Illeg abort uncompl-comp
C0156542|T046|PT|636.92|ICD9CM|Illegally induced abortion, without mention of complication, complete|Illegally induced abortion, without mention of complication, complete
C0156543|T033|HT|637|ICD9CM|Unspecified abortion|Unspecified abortion
C0156545|T046|HT|637.0|ICD9CM|Unspecified abortion complicated by genital tract and pelvic infection|Unspecified abortion complicated by genital tract and pelvic infection
C0156545|T046|AB|637.00|ICD9CM|Abort NOS w pel inf-unsp|Abort NOS w pel inf-unsp
C0156545|T046|PT|637.00|ICD9CM|Unspecified abortion, complicated by genital tract and pelvic infection, unspecified|Unspecified abortion, complicated by genital tract and pelvic infection, unspecified
C0156546|T047|AB|637.01|ICD9CM|Abort NOS w pel inf-inc|Abort NOS w pel inf-inc
C0156546|T047|PT|637.01|ICD9CM|Unspecified abortion, complicated by genital tract and pelvic infection, incomplete|Unspecified abortion, complicated by genital tract and pelvic infection, incomplete
C0156547|T037|AB|637.02|ICD9CM|Abort NOS w pel inf-comp|Abort NOS w pel inf-comp
C0156547|T037|PT|637.02|ICD9CM|Unspecified abortion, complicated by genital tract and pelvic infection, complete|Unspecified abortion, complicated by genital tract and pelvic infection, complete
C0156548|T033|HT|637.1|ICD9CM|Unspecified abortion complicated by delayed or excessive hemorrhage|Unspecified abortion complicated by delayed or excessive hemorrhage
C0156548|T033|AB|637.10|ICD9CM|Abort NOS w hemorr-unsp|Abort NOS w hemorr-unsp
C0156548|T033|PT|637.10|ICD9CM|Unspecified abortion, complicated by delayed or excessive hemorrhage, unspecified|Unspecified abortion, complicated by delayed or excessive hemorrhage, unspecified
C0156550|T046|AB|637.11|ICD9CM|Abort NOS w hemorr-inc|Abort NOS w hemorr-inc
C0156550|T046|PT|637.11|ICD9CM|Unspecified abortion, complicated by delayed or excessive hemorrhage, incomplete|Unspecified abortion, complicated by delayed or excessive hemorrhage, incomplete
C0156551|T037|AB|637.12|ICD9CM|Abort NOS w hemorr-comp|Abort NOS w hemorr-comp
C0156551|T037|PT|637.12|ICD9CM|Unspecified abortion, complicated by delayed or excessive hemorrhage, complete|Unspecified abortion, complicated by delayed or excessive hemorrhage, complete
C1263817|T037|HT|637.2|ICD9CM|Unspecified abortion complicated by damage to pelvic organs or tissues|Unspecified abortion complicated by damage to pelvic organs or tissues
C1263817|T037|AB|637.20|ICD9CM|Ab NOS w pelv damag-unsp|Ab NOS w pelv damag-unsp
C1263817|T037|PT|637.20|ICD9CM|Unspecified abortion, complicated by damage to pelvic organs or tissues, unspecified|Unspecified abortion, complicated by damage to pelvic organs or tissues, unspecified
C0156554|T037|AB|637.21|ICD9CM|Ab NOS w pelv damag-inc|Ab NOS w pelv damag-inc
C0156554|T037|PT|637.21|ICD9CM|Unspecified abortion, complicated by damage to pelvic organs or tissues, incomplete|Unspecified abortion, complicated by damage to pelvic organs or tissues, incomplete
C0156555|T037|AB|637.22|ICD9CM|Ab NOS w pelv damag-comp|Ab NOS w pelv damag-comp
C0156555|T037|PT|637.22|ICD9CM|Unspecified abortion, complicated by damage to pelvic organs or tissues, complete|Unspecified abortion, complicated by damage to pelvic organs or tissues, complete
C0156556|T046|HT|637.3|ICD9CM|Unspecified abortion complicated by renal failure|Unspecified abortion complicated by renal failure
C0156556|T046|AB|637.30|ICD9CM|Ab NOS w renal fail-unsp|Ab NOS w renal fail-unsp
C0156556|T046|PT|637.30|ICD9CM|Unspecified abortion, complicated by renal failure, unspecified|Unspecified abortion, complicated by renal failure, unspecified
C0156558|T037|AB|637.31|ICD9CM|Ab NOS w renal fail-inc|Ab NOS w renal fail-inc
C0156558|T037|PT|637.31|ICD9CM|Unspecified abortion, complicated by renal failure, incomplete|Unspecified abortion, complicated by renal failure, incomplete
C0156559|T037|AB|637.32|ICD9CM|Ab NOS w renal fail-comp|Ab NOS w renal fail-comp
C0156559|T037|PT|637.32|ICD9CM|Unspecified abortion, complicated by renal failure, complete|Unspecified abortion, complicated by renal failure, complete
C0156560|T047|HT|637.4|ICD9CM|Unspecified abortion complicated by metabolic disorder|Unspecified abortion complicated by metabolic disorder
C0156561|T037|AB|637.40|ICD9CM|Ab NOS w metab dis-unsp|Ab NOS w metab dis-unsp
C0156561|T037|PT|637.40|ICD9CM|Unspecified abortion, complicated by metabolic disorder, unspecified|Unspecified abortion, complicated by metabolic disorder, unspecified
C0156562|T037|AB|637.41|ICD9CM|Ab NOS w metab dis-inc|Ab NOS w metab dis-inc
C0156562|T037|PT|637.41|ICD9CM|Unspecified abortion, complicated by metabolic disorder, incomplete|Unspecified abortion, complicated by metabolic disorder, incomplete
C0156563|T037|AB|637.42|ICD9CM|Ab NOS w metab dis-comp|Ab NOS w metab dis-comp
C0156563|T037|PT|637.42|ICD9CM|Unspecified abortion, complicated by metabolic disorder, complete|Unspecified abortion, complicated by metabolic disorder, complete
C0156564|T046|HT|637.5|ICD9CM|Unspecified abortion complicated by shock|Unspecified abortion complicated by shock
C0156564|T046|AB|637.50|ICD9CM|Abort NOS w shock-unsp|Abort NOS w shock-unsp
C0156564|T046|PT|637.50|ICD9CM|Unspecified abortion, complicated by shock, unspecified|Unspecified abortion, complicated by shock, unspecified
C0156566|T037|AB|637.51|ICD9CM|Abort NOS w shock-inc|Abort NOS w shock-inc
C0156566|T037|PT|637.51|ICD9CM|Unspecified abortion, complicated by shock, incomplete|Unspecified abortion, complicated by shock, incomplete
C0156567|T037|AB|637.52|ICD9CM|Abort NOS w shock-comp|Abort NOS w shock-comp
C0156567|T037|PT|637.52|ICD9CM|Unspecified abortion, complicated by shock, complete|Unspecified abortion, complicated by shock, complete
C0156568|T047|HT|637.6|ICD9CM|Unspecified abortion complicated by embolism|Unspecified abortion complicated by embolism
C0156568|T047|AB|637.60|ICD9CM|Ab NOS w embolism-unsp|Ab NOS w embolism-unsp
C0156568|T047|PT|637.60|ICD9CM|Unspecified abortion, complicated by embolism, unspecified|Unspecified abortion, complicated by embolism, unspecified
C0156570|T047|AB|637.61|ICD9CM|Ab NOS w embolism-inc|Ab NOS w embolism-inc
C0156570|T047|PT|637.61|ICD9CM|Unspecified abortion, complicated by embolism, incomplete|Unspecified abortion, complicated by embolism, incomplete
C0156571|T037|AB|637.62|ICD9CM|Ab NOS w embolism-comp|Ab NOS w embolism-comp
C0156571|T037|PT|637.62|ICD9CM|Unspecified abortion, complicated by embolism, complete|Unspecified abortion, complicated by embolism, complete
C0156572|T046|HT|637.7|ICD9CM|Unspecified abortion with other specified complications|Unspecified abortion with other specified complications
C0156573|T037|AB|637.70|ICD9CM|Ab NOS w compl NEC-unsp|Ab NOS w compl NEC-unsp
C0156573|T037|PT|637.70|ICD9CM|Unspecified abortion, with other specified complications, unspecified|Unspecified abortion, with other specified complications, unspecified
C0156574|T046|AB|637.71|ICD9CM|Ab NOS w compl NEC-inc|Ab NOS w compl NEC-inc
C0156574|T046|PT|637.71|ICD9CM|Unspecified abortion, with other specified complications, incomplete|Unspecified abortion, with other specified complications, incomplete
C0156575|T046|AB|637.72|ICD9CM|Ab NOS w compl NEC-comp|Ab NOS w compl NEC-comp
C0156575|T046|PT|637.72|ICD9CM|Unspecified abortion, with other specified complications, complete|Unspecified abortion, with other specified complications, complete
C1299558|T046|HT|637.8|ICD9CM|Unspecified abortion with unspecified complication|Unspecified abortion with unspecified complication
C1299558|T046|AB|637.80|ICD9CM|Ab NOS w compl NOS-unsp|Ab NOS w compl NOS-unsp
C1299558|T046|PT|637.80|ICD9CM|Unspecified abortion, with unspecified complication, unspecified|Unspecified abortion, with unspecified complication, unspecified
C0156578|T046|AB|637.81|ICD9CM|Ab NOS w compl NOS-inc|Ab NOS w compl NOS-inc
C0156578|T046|PT|637.81|ICD9CM|Unspecified abortion, with unspecified complication, incomplete|Unspecified abortion, with unspecified complication, incomplete
C0156579|T046|AB|637.82|ICD9CM|Ab NOS w compl NOS-comp|Ab NOS w compl NOS-comp
C0156579|T046|PT|637.82|ICD9CM|Unspecified abortion, with unspecified complication, complete|Unspecified abortion, with unspecified complication, complete
C0156580|T046|HT|637.9|ICD9CM|Unspecified abortion without mention of complication|Unspecified abortion without mention of complication
C0156580|T046|AB|637.90|ICD9CM|Ab NOS uncomplicat-unsp|Ab NOS uncomplicat-unsp
C0156580|T046|PT|637.90|ICD9CM|Unspecified abortion, without mention of complication, unspecified|Unspecified abortion, without mention of complication, unspecified
C0156581|T037|AB|637.91|ICD9CM|Ab NOS uncomplicat-inc|Ab NOS uncomplicat-inc
C0156581|T037|PT|637.91|ICD9CM|Unspecified abortion, without mention of complication, incomplete|Unspecified abortion, without mention of complication, incomplete
C0156582|T037|AB|637.92|ICD9CM|Ab NOS uncomplicat-comp|Ab NOS uncomplicat-comp
C0156582|T037|PT|637.92|ICD9CM|Unspecified abortion, without mention of complication, complete|Unspecified abortion, without mention of complication, complete
C0392536|T046|HT|638|ICD9CM|Failed attempted abortion|Failed attempted abortion
C0156584|T037|AB|638.0|ICD9CM|Attem abort w pelvic inf|Attem abort w pelvic inf
C0156584|T037|PT|638.0|ICD9CM|Failed attempted abortion complicated by genital tract and pelvic infection|Failed attempted abortion complicated by genital tract and pelvic infection
C0156585|T046|AB|638.1|ICD9CM|Attem abort w hemorrhage|Attem abort w hemorrhage
C0156585|T046|PT|638.1|ICD9CM|Failed attempted abortion complicated by delayed or excessive hemorrhage|Failed attempted abortion complicated by delayed or excessive hemorrhage
C0269561|T037|AB|638.2|ICD9CM|Attem abort w pelv damag|Attem abort w pelv damag
C0269561|T037|PT|638.2|ICD9CM|Failed attempted abortion complicated by damage to pelvic organs or tissues|Failed attempted abortion complicated by damage to pelvic organs or tissues
C0156587|T046|AB|638.3|ICD9CM|Attem abort w renal fail|Attem abort w renal fail
C0156587|T046|PT|638.3|ICD9CM|Failed attempted abortion complicated by renal failure|Failed attempted abortion complicated by renal failure
C0156588|T047|AB|638.4|ICD9CM|Attem abor w metabol dis|Attem abor w metabol dis
C0156588|T047|PT|638.4|ICD9CM|Failed attempted abortion complicated by metabolic disorder|Failed attempted abortion complicated by metabolic disorder
C0156589|T046|AB|638.5|ICD9CM|Attem abortion w shock|Attem abortion w shock
C0156589|T046|PT|638.5|ICD9CM|Failed attempted abortion complicated by shock|Failed attempted abortion complicated by shock
C0156590|T046|AB|638.6|ICD9CM|Attemp abort w embolism|Attemp abort w embolism
C0156590|T046|PT|638.6|ICD9CM|Failed attempted abortion complicated by embolism|Failed attempted abortion complicated by embolism
C0156591|T046|AB|638.7|ICD9CM|Attemp abort w compl NEC|Attemp abort w compl NEC
C0156591|T046|PT|638.7|ICD9CM|Failed attempted abortion with other specified complications|Failed attempted abortion with other specified complications
C0156592|T046|AB|638.8|ICD9CM|Attemp abort w compl NOS|Attemp abort w compl NOS
C0156592|T046|PT|638.8|ICD9CM|Failed attempted abortion with unspecified complication|Failed attempted abortion with unspecified complication
C0269549|T046|AB|638.9|ICD9CM|Attempted abort uncompl|Attempted abort uncompl
C0269549|T046|PT|638.9|ICD9CM|Failed attempted abortion without mention of complication|Failed attempted abortion without mention of complication
C0477810|T046|HT|639|ICD9CM|Complications following abortion or ectopic and molar pregnancies|Complications following abortion or ectopic and molar pregnancies
C0269294|T046|PT|639.0|ICD9CM|Genital tract and pelvic infection following abortion or ectopic and molar pregnancies|Genital tract and pelvic infection following abortion or ectopic and molar pregnancies
C0269294|T046|AB|639.0|ICD9CM|Postabortion gu infect|Postabortion gu infect
C0495168|T046|PT|639.1|ICD9CM|Delayed or excessive hemorrhage following abortion or ectopic and molar pregnancies|Delayed or excessive hemorrhage following abortion or ectopic and molar pregnancies
C0495168|T046|AB|639.1|ICD9CM|Postabortion hemorrhage|Postabortion hemorrhage
C0495173|T037|PT|639.2|ICD9CM|Damage to pelvic organs and tissues following abortion or ectopic and molar pregnancies|Damage to pelvic organs and tissues following abortion or ectopic and molar pregnancies
C0495173|T037|AB|639.2|ICD9CM|Postabort pelvic damage|Postabort pelvic damage
C2712637|T046|PT|639.3|ICD9CM|Kidney failure following abortion and ectopic and molar pregnancies|Kidney failure following abortion and ectopic and molar pregnancies
C2712637|T046|AB|639.3|ICD9CM|Postabort kidney failure|Postabort kidney failure
C0495172|T046|PT|639.4|ICD9CM|Metabolic disorders following abortion or ectopic and molar pregnancies|Metabolic disorders following abortion or ectopic and molar pregnancies
C0495172|T046|AB|639.4|ICD9CM|Postabort metabolic dis|Postabort metabolic dis
C0495170|T046|AB|639.5|ICD9CM|Postabortion shock|Postabortion shock
C0495170|T046|PT|639.5|ICD9CM|Shock following abortion or ectopic and molar pregnancies|Shock following abortion or ectopic and molar pregnancies
C0495169|T046|PT|639.6|ICD9CM|Embolism following abortion or ectopic and molar pregnancies|Embolism following abortion or ectopic and molar pregnancies
C0495169|T046|AB|639.6|ICD9CM|Postabortion embolism|Postabortion embolism
C0156602|T047|PT|639.8|ICD9CM|Other specified complications following abortion or ectopic and molar pregnancy|Other specified complications following abortion or ectopic and molar pregnancy
C0156602|T047|AB|639.8|ICD9CM|Postabortion compl NEC|Postabortion compl NEC
C0477810|T046|AB|639.9|ICD9CM|Postabortion compl NOS|Postabortion compl NOS
C0477810|T046|PT|639.9|ICD9CM|Unspecified complication following abortion or ectopic and molar pregnancy|Unspecified complication following abortion or ectopic and molar pregnancy
C0156604|T046|HT|640|ICD9CM|Hemorrhage in early pregnancy|Hemorrhage in early pregnancy
C0178295|T046|HT|640-649.99|ICD9CM|COMPLICATIONS MAINLY RELATED TO PREGNANCY|COMPLICATIONS MAINLY RELATED TO PREGNANCY
C0000821|T046|HT|640.0|ICD9CM|Threatened abortion|Threatened abortion
C0156605|T047|AB|640.00|ICD9CM|Threatened abort-unspec|Threatened abort-unspec
C0156605|T047|PT|640.00|ICD9CM|Threatened abortion, unspecified as to episode of care or not applicable|Threatened abortion, unspecified as to episode of care or not applicable
C0156606|T046|AB|640.01|ICD9CM|Threatened abort-deliver|Threatened abort-deliver
C0156606|T046|PT|640.01|ICD9CM|Threatened abortion, delivered, with or without mention of antepartum condition|Threatened abortion, delivered, with or without mention of antepartum condition
C0000821|T046|AB|640.03|ICD9CM|Threaten abort-antepart|Threaten abort-antepart
C0000821|T046|PT|640.03|ICD9CM|Threatened abortion, antepartum condition or complication|Threatened abortion, antepartum condition or complication
C0156608|T046|HT|640.8|ICD9CM|Other specified hemorrhage in early pregnancy|Other specified hemorrhage in early pregnancy
C0156609|T046|AB|640.80|ICD9CM|Hem early preg NEC-unsp|Hem early preg NEC-unsp
C0156609|T046|PT|640.80|ICD9CM|Other specified hemorrhage in early pregnancy, unspecified as to episode of care or not applicable|Other specified hemorrhage in early pregnancy, unspecified as to episode of care or not applicable
C0156610|T047|AB|640.81|ICD9CM|Hem early preg NEC-deliv|Hem early preg NEC-deliv
C0269607|T046|AB|640.83|ICD9CM|Hem early pg NEC-antepar|Hem early pg NEC-antepar
C0269607|T046|PT|640.83|ICD9CM|Other specified hemorrhage in early pregnancy, antepartum condition or complication|Other specified hemorrhage in early pregnancy, antepartum condition or complication
C0156604|T046|HT|640.9|ICD9CM|Unspecified hemorrhage in early pregnancy|Unspecified hemorrhage in early pregnancy
C0156613|T046|AB|640.90|ICD9CM|Hemorr early preg-unspec|Hemorr early preg-unspec
C0156613|T046|PT|640.90|ICD9CM|Unspecified hemorrhage in early pregnancy, unspecified as to episode of care or not applicable|Unspecified hemorrhage in early pregnancy, unspecified as to episode of care or not applicable
C0156614|T047|AB|640.91|ICD9CM|Hem early preg-delivered|Hem early preg-delivered
C0269599|T046|AB|640.93|ICD9CM|Hem early preg-antepart|Hem early preg-antepart
C0269599|T046|PT|640.93|ICD9CM|Unspecified hemorrhage in early pregnancy, antepartum condition or complication|Unspecified hemorrhage in early pregnancy, antepartum condition or complication
C0156616|T046|HT|641|ICD9CM|Antepartum hemorrhage, abruptio placentae, and placenta previa|Antepartum hemorrhage, abruptio placentae, and placenta previa
C0156617|T046|HT|641.0|ICD9CM|Placenta previa without hemorrhage|Placenta previa without hemorrhage
C0156618|T047|PT|641.00|ICD9CM|Placenta previa without hemorrhage, unspecified as to episode of care or not applicable|Placenta previa without hemorrhage, unspecified as to episode of care or not applicable
C0156618|T047|AB|641.00|ICD9CM|Placenta previa-unspec|Placenta previa-unspec
C0156619|T047|PT|641.01|ICD9CM|Placenta previa without hemorrhage, delivered, with or without mention of antepartum condition|Placenta previa without hemorrhage, delivered, with or without mention of antepartum condition
C0156619|T047|AB|641.01|ICD9CM|Placenta previa-deliver|Placenta previa-deliver
C0156620|T047|PT|641.03|ICD9CM|Placenta previa without hemorrhage, antepartum condition or complication|Placenta previa without hemorrhage, antepartum condition or complication
C0156620|T047|AB|641.03|ICD9CM|Placenta previa-antepart|Placenta previa-antepart
C0156621|T046|HT|641.1|ICD9CM|Hemorrhage from placenta previa|Hemorrhage from placenta previa
C0156621|T046|PT|641.10|ICD9CM|Hemorrhage from placenta previa, unspecified as to episode of care or not applicable|Hemorrhage from placenta previa, unspecified as to episode of care or not applicable
C0156621|T046|AB|641.10|ICD9CM|Placenta prev hem-unspec|Placenta prev hem-unspec
C0156623|T047|PT|641.11|ICD9CM|Hemorrhage from placenta previa, delivered, with or without mention of antepartum condition|Hemorrhage from placenta previa, delivered, with or without mention of antepartum condition
C0156623|T047|AB|641.11|ICD9CM|Placenta prev hem-deliv|Placenta prev hem-deliv
C0156624|T047|PT|641.13|ICD9CM|Hemorrhage from placenta previa, antepartum condition or complication|Hemorrhage from placenta previa, antepartum condition or complication
C0156624|T047|AB|641.13|ICD9CM|Placen prev hem-antepart|Placen prev hem-antepart
C0000832|T046|HT|641.2|ICD9CM|Premature separation of placenta|Premature separation of placenta
C0000832|T046|AB|641.20|ICD9CM|Prem separ placen-unspec|Prem separ placen-unspec
C0000832|T046|PT|641.20|ICD9CM|Premature separation of placenta, unspecified as to episode of care or not applicable|Premature separation of placenta, unspecified as to episode of care or not applicable
C0156626|T047|AB|641.21|ICD9CM|Prem separ placen-deliv|Prem separ placen-deliv
C0156626|T047|PT|641.21|ICD9CM|Premature separation of placenta, delivered, with or without mention of antepartum condition|Premature separation of placenta, delivered, with or without mention of antepartum condition
C0156627|T047|AB|641.23|ICD9CM|Prem separ plac-antepart|Prem separ plac-antepart
C0156627|T047|PT|641.23|ICD9CM|Premature separation of placenta, antepartum condition or complication|Premature separation of placenta, antepartum condition or complication
C0156631|T046|HT|641.3|ICD9CM|Antepartum hemorrhage associated with coagulation defects|Antepartum hemorrhage associated with coagulation defects
C0156629|T047|AB|641.30|ICD9CM|Coag def hemorr-unspec|Coag def hemorr-unspec
C0156630|T047|AB|641.31|ICD9CM|Coag def hemorr-deliver|Coag def hemorr-deliver
C0156631|T046|PT|641.33|ICD9CM|Antepartum hemorrhage associated with coagulation defects, antepartum condition or complication|Antepartum hemorrhage associated with coagulation defects, antepartum condition or complication
C0156631|T046|AB|641.33|ICD9CM|Coag def hemorr-antepart|Coag def hemorr-antepart
C0156635|T046|HT|641.8|ICD9CM|Other antepartum hemorrhage|Other antepartum hemorrhage
C0156633|T046|AB|641.80|ICD9CM|Antepart hem NEC-unspec|Antepart hem NEC-unspec
C0156633|T046|PT|641.80|ICD9CM|Other antepartum hemorrhage, unspecified as to episode of care or not applicable|Other antepartum hemorrhage, unspecified as to episode of care or not applicable
C0156634|T047|AB|641.81|ICD9CM|Antepartum hem NEC-deliv|Antepartum hem NEC-deliv
C0156634|T047|PT|641.81|ICD9CM|Other antepartum hemorrhage, delivered, with or without mention of antepartum condition|Other antepartum hemorrhage, delivered, with or without mention of antepartum condition
C0156635|T046|AB|641.83|ICD9CM|Antepart hem NEC-antepar|Antepart hem NEC-antepar
C0156635|T046|PT|641.83|ICD9CM|Other antepartum hemorrhage, antepartum condition or complication|Other antepartum hemorrhage, antepartum condition or complication
C0269608|T046|HT|641.9|ICD9CM|Unspecified antepartum hemorrhage|Unspecified antepartum hemorrhage
C0156637|T046|AB|641.90|ICD9CM|Antepart hem NOS-unspec|Antepart hem NOS-unspec
C0156637|T046|PT|641.90|ICD9CM|Unspecified antepartum hemorrhage, unspecified as to episode of care or not applicable|Unspecified antepartum hemorrhage, unspecified as to episode of care or not applicable
C0156638|T047|AB|641.91|ICD9CM|Antepartum hem NOS-deliv|Antepartum hem NOS-deliv
C0156638|T047|PT|641.91|ICD9CM|Unspecified antepartum hemorrhage, delivered, with or without mention of antepartum condition|Unspecified antepartum hemorrhage, delivered, with or without mention of antepartum condition
C0269608|T046|AB|641.93|ICD9CM|Antepart hem NOS-antepar|Antepart hem NOS-antepar
C0269608|T046|PT|641.93|ICD9CM|Unspecified antepartum hemorrhage, antepartum condition or complication|Unspecified antepartum hemorrhage, antepartum condition or complication
C0341909|T047|HT|642|ICD9CM|Hypertension complicating pregnancy, childbirth, and the puerperium|Hypertension complicating pregnancy, childbirth, and the puerperium
C0341930|T047|HT|642.0|ICD9CM|Benign essential hypertension complicating pregnancy, childbirth, and the puerperium|Benign essential hypertension complicating pregnancy, childbirth, and the puerperium
C0156642|T047|AB|642.00|ICD9CM|Essen hyperten preg-unsp|Essen hyperten preg-unsp
C0156643|T047|AB|642.01|ICD9CM|Essen hyperten-delivered|Essen hyperten-delivered
C0156644|T047|AB|642.02|ICD9CM|Essen hyperten-del w p/p|Essen hyperten-del w p/p
C0156645|T047|AB|642.03|ICD9CM|Essen hyperten-antepart|Essen hyperten-antepart
C0156646|T047|AB|642.04|ICD9CM|Essen hyperten-postpart|Essen hyperten-postpart
C0156647|T047|HT|642.1|ICD9CM|Hypertension secondary to renal disease, complicating pregnancy, childbirth, and the puerperium|Hypertension secondary to renal disease, complicating pregnancy, childbirth, and the puerperium
C0156648|T047|AB|642.10|ICD9CM|Renal hyperten preg-unsp|Renal hyperten preg-unsp
C0156649|T047|AB|642.11|ICD9CM|Renal hyperten pg-deliv|Renal hyperten pg-deliv
C0156650|T047|AB|642.12|ICD9CM|Renal hyperten-del p/p|Renal hyperten-del p/p
C0156651|T047|AB|642.13|ICD9CM|Renal hyperten-antepart|Renal hyperten-antepart
C0156652|T047|AB|642.14|ICD9CM|Renal hyperten-postpart|Renal hyperten-postpart
C0156653|T047|HT|642.2|ICD9CM|Other pre-existing hypertension complicating pregnancy, childbirth, and the puerperium|Other pre-existing hypertension complicating pregnancy, childbirth, and the puerperium
C0156654|T047|AB|642.20|ICD9CM|Old hyperten preg-unspec|Old hyperten preg-unspec
C0156655|T047|AB|642.21|ICD9CM|Old hyperten NEC-deliver|Old hyperten NEC-deliver
C0156656|T047|AB|642.22|ICD9CM|Old hyperten-deliv w p/p|Old hyperten-deliv w p/p
C0156657|T047|AB|642.23|ICD9CM|Old hyperten NEC-antepar|Old hyperten NEC-antepar
C0156658|T047|AB|642.24|ICD9CM|Old hyperten NEC-postpar|Old hyperten NEC-postpar
C0341934|T046|HT|642.3|ICD9CM|Transient hypertension of pregnancy|Transient hypertension of pregnancy
C0156659|T047|AB|642.30|ICD9CM|Trans hyperten preg-unsp|Trans hyperten preg-unsp
C0156659|T047|PT|642.30|ICD9CM|Transient hypertension of pregnancy, unspecified as to episode of care or not applicable|Transient hypertension of pregnancy, unspecified as to episode of care or not applicable
C0156660|T047|AB|642.31|ICD9CM|Trans hyperten-delivered|Trans hyperten-delivered
C0156660|T047|PT|642.31|ICD9CM|Transient hypertension of pregnancy, delivered , with or without mention of antepartum condition|Transient hypertension of pregnancy, delivered , with or without mention of antepartum condition
C0156661|T047|AB|642.32|ICD9CM|Trans hyperten-del w p/p|Trans hyperten-del w p/p
C0156661|T047|PT|642.32|ICD9CM|Transient hypertension of pregnancy, delivered, with mention of postpartum complication|Transient hypertension of pregnancy, delivered, with mention of postpartum complication
C0156662|T047|AB|642.33|ICD9CM|Trans hyperten-antepart|Trans hyperten-antepart
C0156662|T047|PT|642.33|ICD9CM|Transient hypertension of pregnancy, antepartum condition or complication|Transient hypertension of pregnancy, antepartum condition or complication
C0156663|T047|AB|642.34|ICD9CM|Trans hyperten-postpart|Trans hyperten-postpart
C0156663|T047|PT|642.34|ICD9CM|Transient hypertension of pregnancy, postpartum condition or complication|Transient hypertension of pregnancy, postpartum condition or complication
C0269658|T046|HT|642.4|ICD9CM|Mild or unspecified pre-eclampsia|Mild or unspecified pre-eclampsia
C0156664|T047|PT|642.40|ICD9CM|Mild or unspecified pre-eclampsia, unspecified as to episode of care or not applicable|Mild or unspecified pre-eclampsia, unspecified as to episode of care or not applicable
C0156664|T047|AB|642.40|ICD9CM|Mild/NOS preeclamp-unsp|Mild/NOS preeclamp-unsp
C0156665|T047|PT|642.41|ICD9CM|Mild or unspecified pre-eclampsia, delivered, with or without mention of antepartum condition|Mild or unspecified pre-eclampsia, delivered, with or without mention of antepartum condition
C0156665|T047|AB|642.41|ICD9CM|Mild/NOS preeclamp-deliv|Mild/NOS preeclamp-deliv
C0156666|T047|PT|642.42|ICD9CM|Mild or unspecified pre-eclampsia, delivered, with mention of postpartum complication|Mild or unspecified pre-eclampsia, delivered, with mention of postpartum complication
C0156666|T047|AB|642.42|ICD9CM|Mild preeclamp-del w p/p|Mild preeclamp-del w p/p
C0156667|T047|PT|642.43|ICD9CM|Mild or unspecified pre-eclampsia, antepartum condition or complication|Mild or unspecified pre-eclampsia, antepartum condition or complication
C0156667|T047|AB|642.43|ICD9CM|Mild/NOS preeclamp-antep|Mild/NOS preeclamp-antep
C0156668|T047|PT|642.44|ICD9CM|Mild or unspecified pre-eclampsia, postpartum condition or complication|Mild or unspecified pre-eclampsia, postpartum condition or complication
C0156668|T047|AB|642.44|ICD9CM|Mild/NOS preeclamp-p/p|Mild/NOS preeclamp-p/p
C0341950|T046|HT|642.5|ICD9CM|Severe pre-eclampsia|Severe pre-eclampsia
C0156669|T047|PT|642.50|ICD9CM|Severe pre-eclampsia, unspecified as to episode of care or not applicable|Severe pre-eclampsia, unspecified as to episode of care or not applicable
C0156669|T047|AB|642.50|ICD9CM|Severe preeclamp-unspec|Severe preeclamp-unspec
C0156670|T047|PT|642.51|ICD9CM|Severe pre-eclampsia, delivered, with or without mention of antepartum condition|Severe pre-eclampsia, delivered, with or without mention of antepartum condition
C0156670|T047|AB|642.51|ICD9CM|Severe preeclamp-deliver|Severe preeclamp-deliver
C0156671|T047|AB|642.52|ICD9CM|Sev preeclamp-del w p/p|Sev preeclamp-del w p/p
C0156671|T047|PT|642.52|ICD9CM|Severe pre-eclampsia, delivered, with mention of postpartum complication|Severe pre-eclampsia, delivered, with mention of postpartum complication
C0156672|T047|AB|642.53|ICD9CM|Sev preeclamp-antepartum|Sev preeclamp-antepartum
C0156672|T047|PT|642.53|ICD9CM|Severe pre-eclampsia, antepartum condition or complication|Severe pre-eclampsia, antepartum condition or complication
C0156673|T047|AB|642.54|ICD9CM|Sev preeclamp-postpartum|Sev preeclamp-postpartum
C0156673|T047|PT|642.54|ICD9CM|Severe pre-eclampsia, postpartum condition or complication|Severe pre-eclampsia, postpartum condition or complication
C0260338|T047|HT|642.6|ICD9CM|Eclampsia complicating pregnancy, childbirth or the puerperium|Eclampsia complicating pregnancy, childbirth or the puerperium
C0156674|T047|AB|642.60|ICD9CM|Eclampsia-unspecified|Eclampsia-unspecified
C0156674|T047|PT|642.60|ICD9CM|Eclampsia, unspecified as to episode of care or not applicable|Eclampsia, unspecified as to episode of care or not applicable
C0156675|T047|AB|642.61|ICD9CM|Eclampsia-delivered|Eclampsia-delivered
C0156675|T047|PT|642.61|ICD9CM|Eclampsia, delivered, with or without mention of antepartum condition|Eclampsia, delivered, with or without mention of antepartum condition
C0156676|T047|AB|642.62|ICD9CM|Eclampsia-deliv w p/p|Eclampsia-deliv w p/p
C0156676|T047|PT|642.62|ICD9CM|Eclampsia, delivered, with mention of postpartum complication|Eclampsia, delivered, with mention of postpartum complication
C0156677|T046|AB|642.63|ICD9CM|Eclampsia-antepartum|Eclampsia-antepartum
C0156677|T046|PT|642.63|ICD9CM|Eclampsia, antepartum condition or complication|Eclampsia, antepartum condition or complication
C0156678|T047|AB|642.64|ICD9CM|Eclampsia-postpartum|Eclampsia-postpartum
C0156678|T047|PT|642.64|ICD9CM|Eclampsia, postpartum condition or complication|Eclampsia, postpartum condition or complication
C0156679|T047|HT|642.7|ICD9CM|Pre-eclampsia or eclampsia superimposed on pre-existing hypertension|Pre-eclampsia or eclampsia superimposed on pre-existing hypertension
C0156680|T047|AB|642.70|ICD9CM|Tox w old hyperten-unsp|Tox w old hyperten-unsp
C0156681|T047|AB|642.71|ICD9CM|Tox w old hyperten-deliv|Tox w old hyperten-deliv
C0156682|T047|AB|642.72|ICD9CM|Tox w old hyp-del w p/p|Tox w old hyp-del w p/p
C0156683|T047|AB|642.73|ICD9CM|Tox w old hyper-antepart|Tox w old hyper-antepart
C0156684|T047|AB|642.74|ICD9CM|Tox w old hyper-postpart|Tox w old hyper-postpart
C1261262|T047|HT|642.9|ICD9CM|Unspecified hypertension complicating pregnancy, childbirth, or the puerperium|Unspecified hypertension complicating pregnancy, childbirth, or the puerperium
C0156686|T047|AB|642.90|ICD9CM|Hyperten preg NOS-unspec|Hyperten preg NOS-unspec
C0156687|T047|AB|642.91|ICD9CM|Hypertens NOS-delivered|Hypertens NOS-delivered
C0156688|T047|AB|642.92|ICD9CM|Hypertens NOS-del w p/p|Hypertens NOS-del w p/p
C0156689|T047|AB|642.93|ICD9CM|Hypertens NOS-antepartum|Hypertens NOS-antepartum
C0156690|T047|AB|642.94|ICD9CM|Hypertens NOS-postpartum|Hypertens NOS-postpartum
C0020450|T184|HT|643|ICD9CM|Excessive vomiting in pregnancy|Excessive vomiting in pregnancy
C0020451|T047|HT|643.0|ICD9CM|Mild hyperemesis gravidarum|Mild hyperemesis gravidarum
C0156692|T047|AB|643.00|ICD9CM|Mild hyperem grav-unspec|Mild hyperem grav-unspec
C0156692|T047|PT|643.00|ICD9CM|Mild hyperemesis gravidarum, unspecified as to episode of care or not applicable|Mild hyperemesis gravidarum, unspecified as to episode of care or not applicable
C0156693|T047|AB|643.01|ICD9CM|Mild hyperem grav-deliv|Mild hyperem grav-deliv
C0156693|T047|PT|643.01|ICD9CM|Mild hyperemesis gravidarum, delivered, with or without mention of antepartum condition|Mild hyperemesis gravidarum, delivered, with or without mention of antepartum condition
C0156694|T047|PT|643.03|ICD9CM|Mild hyperemesis gravidarum, antepartum condition or complication|Mild hyperemesis gravidarum, antepartum condition or complication
C0156694|T047|AB|643.03|ICD9CM|Mild hyperemesis-antepar|Mild hyperemesis-antepar
C0405080|T047|HT|643.1|ICD9CM|Hyperemesis gravidarum with metabolic disturbance|Hyperemesis gravidarum with metabolic disturbance
C0156696|T047|AB|643.10|ICD9CM|Hyperem w metab dis-unsp|Hyperem w metab dis-unsp
C0156697|T047|AB|643.11|ICD9CM|Hyperem w metab dis-del|Hyperem w metab dis-del
C0156698|T047|AB|643.13|ICD9CM|Hyperem w metab-antepart|Hyperem w metab-antepart
C0156698|T047|PT|643.13|ICD9CM|Hyperemesis gravidarum with metabolic disturbance, antepartum condition or complication|Hyperemesis gravidarum with metabolic disturbance, antepartum condition or complication
C0156699|T046|HT|643.2|ICD9CM|Late vomiting of pregnancy|Late vomiting of pregnancy
C0156700|T047|AB|643.20|ICD9CM|Late vomit of preg-unsp|Late vomit of preg-unsp
C0156700|T047|PT|643.20|ICD9CM|Late vomiting of pregnancy, unspecified as to episode of care or not applicable|Late vomiting of pregnancy, unspecified as to episode of care or not applicable
C0156701|T184|AB|643.21|ICD9CM|Late vomit of preg-deliv|Late vomit of preg-deliv
C0156701|T184|PT|643.21|ICD9CM|Late vomiting of pregnancy, delivered, with or without mention of antepartum condition|Late vomiting of pregnancy, delivered, with or without mention of antepartum condition
C0156702|T047|AB|643.23|ICD9CM|Late vomit preg-antepart|Late vomit preg-antepart
C0156702|T047|PT|643.23|ICD9CM|Late vomiting of pregnancy, antepartum condition or complication|Late vomiting of pregnancy, antepartum condition or complication
C0156703|T184|HT|643.8|ICD9CM|Other vomiting complicating pregnancy|Other vomiting complicating pregnancy
C0156704|T047|PT|643.80|ICD9CM|Other vomiting complicating pregnancy, unspecified as to episode of care or not applicable|Other vomiting complicating pregnancy, unspecified as to episode of care or not applicable
C0156704|T047|AB|643.80|ICD9CM|Vomit compl preg-unspec|Vomit compl preg-unspec
C0156705|T047|PT|643.81|ICD9CM|Other vomiting complicating pregnancy, delivered, with or without mention of antepartum condition|Other vomiting complicating pregnancy, delivered, with or without mention of antepartum condition
C0156705|T047|AB|643.81|ICD9CM|Vomit compl preg-deliver|Vomit compl preg-deliver
C0156706|T047|PT|643.83|ICD9CM|Other vomiting complicating pregnancy, antepartum condition or complication|Other vomiting complicating pregnancy, antepartum condition or complication
C0156706|T047|AB|643.83|ICD9CM|Vomit compl preg-antepar|Vomit compl preg-antepar
C0269661|T046|HT|643.9|ICD9CM|Unspecified vomiting of pregnancy|Unspecified vomiting of pregnancy
C0156708|T047|PT|643.90|ICD9CM|Unspecified vomiting of pregnancy, unspecified as to episode of care or not applicable|Unspecified vomiting of pregnancy, unspecified as to episode of care or not applicable
C0156708|T047|AB|643.90|ICD9CM|Vomit of preg NOS-unspec|Vomit of preg NOS-unspec
C0156709|T184|PT|643.91|ICD9CM|Unspecified vomiting of pregnancy, delivered, with or without mention of antepartum condition|Unspecified vomiting of pregnancy, delivered, with or without mention of antepartum condition
C0156709|T184|AB|643.91|ICD9CM|Vomit of preg NOS-deliv|Vomit of preg NOS-deliv
C0156710|T047|PT|643.93|ICD9CM|Unspecified vomiting of pregnancy, antepartum condition or complication|Unspecified vomiting of pregnancy, antepartum condition or complication
C0156710|T047|AB|643.93|ICD9CM|Vomit of pg NOS-antepart|Vomit of pg NOS-antepart
C0156711|T046|HT|644|ICD9CM|Early or threatened labor|Early or threatened labor
C0473390|T046|HT|644.0|ICD9CM|Threatened premature labor|Threatened premature labor
C0156713|T047|AB|644.00|ICD9CM|Threat prem labor-unspec|Threat prem labor-unspec
C0156713|T047|PT|644.00|ICD9CM|Threatened premature labor, unspecified as to episode of care or not applicable|Threatened premature labor, unspecified as to episode of care or not applicable
C0156714|T047|PT|644.03|ICD9CM|Threatened premature labor, antepartum condition or complication|Threatened premature labor, antepartum condition or complication
C0156714|T047|AB|644.03|ICD9CM|Thrt prem labor-antepart|Thrt prem labor-antepart
C0473388|T046|HT|644.1|ICD9CM|Other threatened labor|Other threatened labor
C0156716|T046|PT|644.10|ICD9CM|Other threatened labor, unspecified as to episode of care or not applicable|Other threatened labor, unspecified as to episode of care or not applicable
C0156716|T046|AB|644.10|ICD9CM|Threat labor NEC-unspec|Threat labor NEC-unspec
C0156717|T047|PT|644.13|ICD9CM|Other threatened labor, antepartum condition or complication|Other threatened labor, antepartum condition or complication
C0156717|T047|AB|644.13|ICD9CM|Threat labor NEC-antepar|Threat labor NEC-antepar
C0151526|T046|HT|644.2|ICD9CM|Early onset of delivery|Early onset of delivery
C0156718|T047|AB|644.20|ICD9CM|Early onset deliv-unspec|Early onset deliv-unspec
C0156718|T047|PT|644.20|ICD9CM|Early onset of delivery, unspecified as to episode of care or not applicable|Early onset of delivery, unspecified as to episode of care or not applicable
C0156719|T047|AB|644.21|ICD9CM|Early onset delivery-del|Early onset delivery-del
C0156719|T047|PT|644.21|ICD9CM|Early onset of delivery, delivered, with or without mention of antepartum condition|Early onset of delivery, delivered, with or without mention of antepartum condition
C0878751|T046|HT|645|ICD9CM|Late pregnancy|Late pregnancy
C0032993|T046|HT|645.1|ICD9CM|Post term pregnancy|Post term pregnancy
C1176343|T047|AB|645.10|ICD9CM|Post term preg-unsp|Post term preg-unsp
C1176343|T047|PT|645.10|ICD9CM|Post term pregnancy, unspecified as to episode of care or not applicable|Post term pregnancy, unspecified as to episode of care or not applicable
C1176344|T047|AB|645.11|ICD9CM|Post term preg-del|Post term preg-del
C1176344|T047|PT|645.11|ICD9CM|Post term pregnancy, delivered, with or without mention of antepartum condition|Post term pregnancy, delivered, with or without mention of antepartum condition
C1176345|T047|AB|645.13|ICD9CM|Post term preg-antepar|Post term preg-antepar
C1176345|T047|PT|645.13|ICD9CM|Post term pregnancy, antepartum condition or complication|Post term pregnancy, antepartum condition or complication
C0032993|T046|HT|645.2|ICD9CM|Prolonged pregnancy|Prolonged pregnancy
C1176346|T047|AB|645.20|ICD9CM|Prolonged preg-unsp|Prolonged preg-unsp
C1176346|T047|PT|645.20|ICD9CM|Prolonged pregnancy, unspecified as to episode of care or not applicable|Prolonged pregnancy, unspecified as to episode of care or not applicable
C1176347|T047|AB|645.21|ICD9CM|Prolonged preg-del|Prolonged preg-del
C1176347|T047|PT|645.21|ICD9CM|Prolonged pregnancy, delivered, with or without mention of antepartum condition|Prolonged pregnancy, delivered, with or without mention of antepartum condition
C1176348|T047|AB|645.23|ICD9CM|Prolonged preg-antepar|Prolonged preg-antepar
C1176348|T047|PT|645.23|ICD9CM|Prolonged pregnancy, antepartum condition or complication|Prolonged pregnancy, antepartum condition or complication
C0869265|T046|HT|646|ICD9CM|Other complications of pregnancy, not elsewhere classified|Other complications of pregnancy, not elsewhere classified
C0156724|T019|HT|646.0|ICD9CM|Papyraceous fetus|Papyraceous fetus
C0156725|T047|AB|646.00|ICD9CM|Papyraceous fetus-unspec|Papyraceous fetus-unspec
C0156725|T047|PT|646.00|ICD9CM|Papyraceous fetus, unspecified as to episode of care or not applicable|Papyraceous fetus, unspecified as to episode of care or not applicable
C0156726|T047|AB|646.01|ICD9CM|Papyraceous fetus-deliv|Papyraceous fetus-deliv
C0156726|T047|PT|646.01|ICD9CM|Papyraceous fetus, delivered, with or without mention of antepartum condition|Papyraceous fetus, delivered, with or without mention of antepartum condition
C0156727|T047|AB|646.03|ICD9CM|Papyraceous fet-antepar|Papyraceous fet-antepar
C0156727|T047|PT|646.03|ICD9CM|Papyraceous fetus, antepartum condition or complication|Papyraceous fetus, antepartum condition or complication
C0156728|T046|HT|646.1|ICD9CM|Edema or excessive weight gain in pregnancy, without mention of hypertension|Edema or excessive weight gain in pregnancy, without mention of hypertension
C0156729|T047|AB|646.10|ICD9CM|Edema in preg-unspec|Edema in preg-unspec
C0156730|T047|AB|646.11|ICD9CM|Edema in preg-delivered|Edema in preg-delivered
C0473384|T184|AB|646.12|ICD9CM|Edema in preg-del w p/p|Edema in preg-del w p/p
C0815336|T184|AB|646.13|ICD9CM|Edema in preg-antepartum|Edema in preg-antepartum
C0156733|T047|AB|646.14|ICD9CM|Edema in preg-postpartum|Edema in preg-postpartum
C0269673|T047|HT|646.2|ICD9CM|Unspecified renal disease in pregnancy, without mention of hypertension|Unspecified renal disease in pregnancy, without mention of hypertension
C0156738|T047|AB|646.20|ICD9CM|Renal dis preg NOS-unsp|Renal dis preg NOS-unsp
C0156736|T047|AB|646.21|ICD9CM|Renal dis NOS-delivered|Renal dis NOS-delivered
C0156737|T047|AB|646.22|ICD9CM|Renal dis NOS-del w p/p|Renal dis NOS-del w p/p
C0156738|T047|AB|646.23|ICD9CM|Renal dis NOS-antepartum|Renal dis NOS-antepartum
C0156739|T047|AB|646.24|ICD9CM|Renal dis NOS-postpartum|Renal dis NOS-postpartum
C2921106|T046|HT|646.3|ICD9CM|Recurrent pregnancy loss|Recurrent pregnancy loss
C0156741|T047|AB|646.30|ICD9CM|Recur preg loss-unspec|Recur preg loss-unspec
C0156741|T047|PT|646.30|ICD9CM|Recurrent pregnancy loss, unspecified as to episode of care or not applicable|Recurrent pregnancy loss, unspecified as to episode of care or not applicable
C0156742|T047|AB|646.31|ICD9CM|Recurnt preg loss-deliv|Recurnt preg loss-deliv
C0156742|T047|PT|646.31|ICD9CM|Recurrent pregnancy loss, delivered, with or without mention of antepartum condition|Recurrent pregnancy loss, delivered, with or without mention of antepartum condition
C0156743|T047|AB|646.33|ICD9CM|Recurnt preg loss-antep|Recurnt preg loss-antep
C0156743|T047|PT|646.33|ICD9CM|Recurrent pregnancy loss, antepartum condition or complication|Recurrent pregnancy loss, antepartum condition or complication
C0405072|T047|HT|646.4|ICD9CM|Peripheral neuritis in pregnancy|Peripheral neuritis in pregnancy
C0156745|T047|AB|646.40|ICD9CM|Neuritis of preg-unspec|Neuritis of preg-unspec
C0156745|T047|PT|646.40|ICD9CM|Peripheral neuritis in pregnancy, unspecified as to episode of care or not applicable|Peripheral neuritis in pregnancy, unspecified as to episode of care or not applicable
C0156746|T047|AB|646.41|ICD9CM|Neuritis-delivered|Neuritis-delivered
C0156746|T047|PT|646.41|ICD9CM|Peripheral neuritis in pregnancy, delivered, with or without mention of antepartum condition|Peripheral neuritis in pregnancy, delivered, with or without mention of antepartum condition
C0156747|T047|AB|646.42|ICD9CM|Neuritis-delivered w p/p|Neuritis-delivered w p/p
C0156747|T047|PT|646.42|ICD9CM|Peripheral neuritis in pregnancy, delivered, with mention of postpartum complication|Peripheral neuritis in pregnancy, delivered, with mention of postpartum complication
C0405072|T047|AB|646.43|ICD9CM|Neuritis of preg-antepar|Neuritis of preg-antepar
C0405072|T047|PT|646.43|ICD9CM|Peripheral neuritis in pregnancy, antepartum condition or complication|Peripheral neuritis in pregnancy, antepartum condition or complication
C0156749|T047|AB|646.44|ICD9CM|Neuritis of preg-postpar|Neuritis of preg-postpar
C0156749|T047|PT|646.44|ICD9CM|Peripheral neuritis in pregnancy, postpartum condition or complication|Peripheral neuritis in pregnancy, postpartum condition or complication
C0156750|T047|HT|646.5|ICD9CM|Asymptomatic bacteriuria in pregnancy|Asymptomatic bacteriuria in pregnancy
C0156750|T047|PT|646.50|ICD9CM|Asymptomatic bacteriuria in pregnancy, unspecified as to episode of care or not applicable|Asymptomatic bacteriuria in pregnancy, unspecified as to episode of care or not applicable
C0156750|T047|AB|646.50|ICD9CM|Bacteriuria preg-unspec|Bacteriuria preg-unspec
C0156752|T047|AB|646.51|ICD9CM|Asym bacteriuria-deliver|Asym bacteriuria-deliver
C0156752|T047|PT|646.51|ICD9CM|Asymptomatic bacteriuria in pregnancy, delivered, with or without mention of antepartum condition|Asymptomatic bacteriuria in pregnancy, delivered, with or without mention of antepartum condition
C0156753|T047|AB|646.52|ICD9CM|Asy bacteruria-del w p/p|Asy bacteruria-del w p/p
C0156753|T047|PT|646.52|ICD9CM|Asymptomatic bacteriuria in pregnancy, delivered, with mention of postpartum complication|Asymptomatic bacteriuria in pregnancy, delivered, with mention of postpartum complication
C0156750|T047|AB|646.53|ICD9CM|Asy bacteriuria-antepart|Asy bacteriuria-antepart
C0156750|T047|PT|646.53|ICD9CM|Asymptomatic bacteriuria in pregnancy, antepartum condition or complication|Asymptomatic bacteriuria in pregnancy, antepartum condition or complication
C0156755|T047|AB|646.54|ICD9CM|Asy bacteriuria-postpart|Asy bacteriuria-postpart
C0156755|T047|PT|646.54|ICD9CM|Asymptomatic bacteriuria in pregnancy, postpartum condition or complication|Asymptomatic bacteriuria in pregnancy, postpartum condition or complication
C0156756|T046|HT|646.6|ICD9CM|Infections of genitourinary tract in pregnancy|Infections of genitourinary tract in pregnancy
C0156756|T046|AB|646.60|ICD9CM|Gu infect in preg-unspec|Gu infect in preg-unspec
C0156756|T046|PT|646.60|ICD9CM|Infections of genitourinary tract in pregnancy, unspecified as to episode of care or not applicable|Infections of genitourinary tract in pregnancy, unspecified as to episode of care or not applicable
C0156758|T047|AB|646.61|ICD9CM|Gu infection-delivered|Gu infection-delivered
C0156759|T047|AB|646.62|ICD9CM|Gu infection-deliv w p/p|Gu infection-deliv w p/p
C0156759|T047|PT|646.62|ICD9CM|Infections of genitourinary tract in pregnancy, delivered, with mention of postpartum complication|Infections of genitourinary tract in pregnancy, delivered, with mention of postpartum complication
C0156756|T046|AB|646.63|ICD9CM|Gu infection-antepartum|Gu infection-antepartum
C0156756|T046|PT|646.63|ICD9CM|Infections of genitourinary tract in pregnancy, antepartum condition or complication|Infections of genitourinary tract in pregnancy, antepartum condition or complication
C0156761|T047|AB|646.64|ICD9CM|Gu infection-postpartum|Gu infection-postpartum
C0156761|T047|PT|646.64|ICD9CM|Infections of genitourinary tract in pregnancy, postpartum condition or complication|Infections of genitourinary tract in pregnancy, postpartum condition or complication
C3161439|T047|HT|646.7|ICD9CM|Liver and biliary tract disorders in pregnancy|Liver and biliary tract disorders in pregnancy
C0156762|T046|PT|646.70|ICD9CM|Liver and biliary tract disorders in pregnancy, unspecified as to episode of care or not applicable|Liver and biliary tract disorders in pregnancy, unspecified as to episode of care or not applicable
C0156762|T046|AB|646.70|ICD9CM|Liver/bil trct disr-unsp|Liver/bil trct disr-unsp
C0400932|T047|AB|646.71|ICD9CM|Liver/bil trct disr-del|Liver/bil trct disr-del
C0156762|T046|PT|646.73|ICD9CM|Liver and biliary tract disorders in pregnancy, antepartum condition or complication|Liver and biliary tract disorders in pregnancy, antepartum condition or complication
C0156762|T046|AB|646.73|ICD9CM|Liver/bil trct disr-ante|Liver/bil trct disr-ante
C0156769|T046|HT|646.8|ICD9CM|Other specified complications of pregnancy|Other specified complications of pregnancy
C0156769|T046|PT|646.80|ICD9CM|Other specified complications of pregnancy, unspecified as to episode of care or not applicable|Other specified complications of pregnancy, unspecified as to episode of care or not applicable
C0156769|T046|AB|646.80|ICD9CM|Preg compl NEC-unspec|Preg compl NEC-unspec
C0156767|T047|AB|646.81|ICD9CM|Preg compl NEC-delivered|Preg compl NEC-delivered
C0156768|T047|PT|646.82|ICD9CM|Other specified complications of pregnancy, delivered, with mention of postpartum complication|Other specified complications of pregnancy, delivered, with mention of postpartum complication
C0156768|T047|AB|646.82|ICD9CM|Preg compl NEC-del w p/p|Preg compl NEC-del w p/p
C0156769|T046|PT|646.83|ICD9CM|Other specified complications of pregnancy, antepartum condition or complication|Other specified complications of pregnancy, antepartum condition or complication
C0156769|T046|AB|646.83|ICD9CM|Preg compl NEC-antepart|Preg compl NEC-antepart
C0156770|T046|PT|646.84|ICD9CM|Other specified complications of pregnancy, postpartum condition or complication|Other specified complications of pregnancy, postpartum condition or complication
C0156770|T046|AB|646.84|ICD9CM|Preg compl NEC-postpart|Preg compl NEC-postpart
C0032962|T046|HT|646.9|ICD9CM|Unspecified complication of pregnancy|Unspecified complication of pregnancy
C0156771|T047|AB|646.90|ICD9CM|Preg compl NOS-unspec|Preg compl NOS-unspec
C0156771|T047|PT|646.90|ICD9CM|Unspecified complication of pregnancy, unspecified as to episode of care or not applicable|Unspecified complication of pregnancy, unspecified as to episode of care or not applicable
C0156772|T047|AB|646.91|ICD9CM|Preg compl NOS-delivered|Preg compl NOS-delivered
C0156772|T047|PT|646.91|ICD9CM|Unspecified complication of pregnancy, delivered, with or without mention of antepartum condition|Unspecified complication of pregnancy, delivered, with or without mention of antepartum condition
C0156773|T047|AB|646.93|ICD9CM|Preg compl NOS-antepart|Preg compl NOS-antepart
C0156773|T047|PT|646.93|ICD9CM|Unspecified complication of pregnancy, antepartum condition or complication|Unspecified complication of pregnancy, antepartum condition or complication
C0275820|T047|HT|647.0|ICD9CM|Syphilis complicating pregnancy, childbirth, or the puerperium|Syphilis complicating pregnancy, childbirth, or the puerperium
C0156776|T047|AB|647.00|ICD9CM|Syphilis in preg-unspec|Syphilis in preg-unspec
C0156777|T047|AB|647.01|ICD9CM|Syphilis-delivered|Syphilis-delivered
C0156778|T047|AB|647.02|ICD9CM|Syphilis-delivered w p/p|Syphilis-delivered w p/p
C0747833|T047|AB|647.03|ICD9CM|Syphilis-antepartum|Syphilis-antepartum
C0156780|T047|AB|647.04|ICD9CM|Syphilis-postpartum|Syphilis-postpartum
C0275667|T047|HT|647.1|ICD9CM|Gonorrhea complicating pregnancy, childbirth, or the puerperium|Gonorrhea complicating pregnancy, childbirth, or the puerperium
C0156782|T047|AB|647.10|ICD9CM|Gonorrhea in preg-unspec|Gonorrhea in preg-unspec
C0156783|T047|AB|647.11|ICD9CM|Gonorrhea-delivered|Gonorrhea-delivered
C0156784|T047|AB|647.12|ICD9CM|Gonorrhea-deliver w p/p|Gonorrhea-deliver w p/p
C0747817|T047|AB|647.13|ICD9CM|Gonorrhea-antepartum|Gonorrhea-antepartum
C0473333|T033|AB|647.14|ICD9CM|Gonorrhea-postpartum|Gonorrhea-postpartum
C0495308|T047|HT|647.2|ICD9CM|Other venereal diseases in the mother complicating pregnancy, childbirth, or the puerperium|Other venereal diseases in the mother complicating pregnancy, childbirth, or the puerperium
C0156788|T047|AB|647.20|ICD9CM|Other VD in preg-unspec|Other VD in preg-unspec
C0490049|T047|AB|647.21|ICD9CM|Other vd-delivered|Other vd-delivered
C0490050|T047|AB|647.22|ICD9CM|Other vd-delivered w p/p|Other vd-delivered w p/p
C0375389|T047|AB|647.23|ICD9CM|Other vd-antepartum|Other vd-antepartum
C0375390|T047|AB|647.24|ICD9CM|Other vd-postpartum|Other vd-postpartum
C1533626|T046|HT|647.3|ICD9CM|Tuberculosis complicating pregnancy, childbirth, or the puerperium|Tuberculosis complicating pregnancy, childbirth, or the puerperium
C0156794|T047|AB|647.30|ICD9CM|TB in preg-unspecified|TB in preg-unspecified
C0156795|T047|AB|647.31|ICD9CM|Tuberculosis-delivered|Tuberculosis-delivered
C0156796|T047|AB|647.32|ICD9CM|Tuberculosis-deliv w p/p|Tuberculosis-deliv w p/p
C0156797|T047|AB|647.33|ICD9CM|Tuberculosis-antepartum|Tuberculosis-antepartum
C0156798|T047|AB|647.34|ICD9CM|Tuberculosis-postpartum|Tuberculosis-postpartum
C0156799|T047|HT|647.4|ICD9CM|Malaria complicating pregnancy, childbirth, or the puerperium|Malaria complicating pregnancy, childbirth, or the puerperium
C0156800|T047|AB|647.40|ICD9CM|Malaria in preg-unspec|Malaria in preg-unspec
C0156800|T047|PT|647.40|ICD9CM|Malaria in the mother, unspecified as to episode of care or not applicable|Malaria in the mother, unspecified as to episode of care or not applicable
C0156801|T047|PT|647.41|ICD9CM|Malaria in the mother, delivered, with or without mention of antepartum condition|Malaria in the mother, delivered, with or without mention of antepartum condition
C0156801|T047|AB|647.41|ICD9CM|Malaria-delivered|Malaria-delivered
C0156802|T047|PT|647.42|ICD9CM|Malaria in the mother, delivered, with mention of postpartum complication|Malaria in the mother, delivered, with mention of postpartum complication
C0156802|T047|AB|647.42|ICD9CM|Malaria-delivered w p/p|Malaria-delivered w p/p
C0747820|T047|PT|647.43|ICD9CM|Malaria in the mother, antepartum condition or complication|Malaria in the mother, antepartum condition or complication
C0747820|T047|AB|647.43|ICD9CM|Malaria-antepartum|Malaria-antepartum
C0156804|T047|PT|647.44|ICD9CM|Malaria in the mother, postpartum condition or complication|Malaria in the mother, postpartum condition or complication
C0156804|T047|AB|647.44|ICD9CM|Malaria-postpartum|Malaria-postpartum
C0156805|T047|HT|647.5|ICD9CM|Rubella complicating pregnancy, childbirth, or the puerperium|Rubella complicating pregnancy, childbirth, or the puerperium
C0276306|T047|AB|647.50|ICD9CM|Rubella in preg-unspec|Rubella in preg-unspec
C0276306|T047|PT|647.50|ICD9CM|Rubella in the mother, unspecified as to episode of care or not applicable|Rubella in the mother, unspecified as to episode of care or not applicable
C0156807|T047|PT|647.51|ICD9CM|Rubella in the mother, delivered, with or without mention of antepartum condition|Rubella in the mother, delivered, with or without mention of antepartum condition
C0156807|T047|AB|647.51|ICD9CM|Rubella-delivered|Rubella-delivered
C0156808|T047|PT|647.52|ICD9CM|Rubella in the mother, delivered, with mention of postpartum complication|Rubella in the mother, delivered, with mention of postpartum complication
C0156808|T047|AB|647.52|ICD9CM|Rubella-delivered w p/p|Rubella-delivered w p/p
C0156809|T047|PT|647.53|ICD9CM|Rubella in the mother, antepartum condition or complication|Rubella in the mother, antepartum condition or complication
C0156809|T047|AB|647.53|ICD9CM|Rubella-antepartum|Rubella-antepartum
C0156810|T047|PT|647.54|ICD9CM|Rubella in the mother, postpartum condition or complication|Rubella in the mother, postpartum condition or complication
C0156810|T047|AB|647.54|ICD9CM|Rubella-postpartum|Rubella-postpartum
C0477876|T047|HT|647.6|ICD9CM|Other viral diseases complicating pregnancy, childbirth, or the puerperium|Other viral diseases complicating pregnancy, childbirth, or the puerperium
C0156812|T047|AB|647.60|ICD9CM|Oth virus in preg-unspec|Oth virus in preg-unspec
C0156812|T047|PT|647.60|ICD9CM|Other viral diseases in the mother, unspecified as to episode of care or not applicable|Other viral diseases in the mother, unspecified as to episode of care or not applicable
C0156813|T047|AB|647.61|ICD9CM|Oth viral dis-delivered|Oth viral dis-delivered
C0156813|T047|PT|647.61|ICD9CM|Other viral diseases in the mother, delivered, with or without mention of antepartum condition|Other viral diseases in the mother, delivered, with or without mention of antepartum condition
C0156814|T047|AB|647.62|ICD9CM|Oth viral dis-del w p/p|Oth viral dis-del w p/p
C0156814|T047|PT|647.62|ICD9CM|Other viral diseases in the mother, delivered, with mention of postpartum complication|Other viral diseases in the mother, delivered, with mention of postpartum complication
C0156815|T047|AB|647.63|ICD9CM|Oth viral dis-antepartum|Oth viral dis-antepartum
C0156815|T047|PT|647.63|ICD9CM|Other viral diseases in the mother, antepartum condition or complication|Other viral diseases in the mother, antepartum condition or complication
C0156816|T047|AB|647.64|ICD9CM|Oth viral dis-postpartum|Oth viral dis-postpartum
C0156816|T047|PT|647.64|ICD9CM|Other viral diseases in the mother, postpartum condition or complication|Other viral diseases in the mother, postpartum condition or complication
C0156818|T047|AB|647.80|ICD9CM|Inf dis in preg NEC-unsp|Inf dis in preg NEC-unsp
C0156819|T047|AB|647.81|ICD9CM|Infect dis NEC-delivered|Infect dis NEC-delivered
C0156820|T047|AB|647.82|ICD9CM|Infect dis NEC-del w p/p|Infect dis NEC-del w p/p
C0156821|T047|AB|647.83|ICD9CM|Infect dis NEC-antepart|Infect dis NEC-antepart
C0156821|T047|PT|647.83|ICD9CM|Other specified infectious and parasitic diseases of mother, antepartum condition or complication|Other specified infectious and parasitic diseases of mother, antepartum condition or complication
C0156822|T047|AB|647.84|ICD9CM|Infect dis NEC-postpart|Infect dis NEC-postpart
C0156822|T047|PT|647.84|ICD9CM|Other specified infectious and parasitic diseases of mother, postpartum condition or complication|Other specified infectious and parasitic diseases of mother, postpartum condition or complication
C0156823|T047|HT|647.9|ICD9CM|Unspecified infection or infestation complicating pregnancy, childbirth, or the puerperium|Unspecified infection or infestation complicating pregnancy, childbirth, or the puerperium
C0156824|T047|AB|647.90|ICD9CM|Infect in preg NOS-unsp|Infect in preg NOS-unsp
C0156824|T047|PT|647.90|ICD9CM|Unspecified infection or infestation of mother, unspecified as to episode of care or not applicable|Unspecified infection or infestation of mother, unspecified as to episode of care or not applicable
C0156825|T047|AB|647.91|ICD9CM|Infect NOS-delivered|Infect NOS-delivered
C0156826|T047|AB|647.92|ICD9CM|Infect NOS-deliver w p/p|Infect NOS-deliver w p/p
C0156826|T047|PT|647.92|ICD9CM|Unspecified infection or infestation of mother, delivered, with mention of postpartum complication|Unspecified infection or infestation of mother, delivered, with mention of postpartum complication
C0156827|T047|AB|647.93|ICD9CM|Infect NOS-antepartum|Infect NOS-antepartum
C0156827|T047|PT|647.93|ICD9CM|Unspecified infection or infestation of mother, antepartum condition or complication|Unspecified infection or infestation of mother, antepartum condition or complication
C0156828|T047|AB|647.94|ICD9CM|Infect NOS-postpartum|Infect NOS-postpartum
C0156828|T047|PT|647.94|ICD9CM|Unspecified infection or infestation of mother, postpartum condition or complication|Unspecified infection or infestation of mother, postpartum condition or complication
C0341893|T047|HT|648.0|ICD9CM|Diabetes mellitus complicating pregnancy, childbirth, or the puerperium|Diabetes mellitus complicating pregnancy, childbirth, or the puerperium
C0341893|T047|AB|648.00|ICD9CM|Diabetes in preg-unspec|Diabetes in preg-unspec
C0341897|T047|AB|648.01|ICD9CM|Diabetes-delivered|Diabetes-delivered
C0341896|T047|AB|648.02|ICD9CM|Diabetes-delivered w p/p|Diabetes-delivered w p/p
C0032969|T047|AB|648.03|ICD9CM|Diabetes-antepartum|Diabetes-antepartum
C0341894|T047|AB|648.04|ICD9CM|Diabetes-postpartum|Diabetes-postpartum
C0269683|T047|HT|648.1|ICD9CM|Thyroid dysfunction complicating pregnancy, childbirth, or the puerperium|Thyroid dysfunction complicating pregnancy, childbirth, or the puerperium
C0156837|T047|AB|648.10|ICD9CM|Thyroid dysfun preg-unsp|Thyroid dysfun preg-unsp
C0156837|T047|PT|648.10|ICD9CM|Thyroid dysfunction of mother, unspecified as to episode of care or not applicable|Thyroid dysfunction of mother, unspecified as to episode of care or not applicable
C0156838|T047|AB|648.11|ICD9CM|Thyroid dysfunc-deliver|Thyroid dysfunc-deliver
C0156838|T047|PT|648.11|ICD9CM|Thyroid dysfunction of mother, delivered, with or without mention of antepartum condition|Thyroid dysfunction of mother, delivered, with or without mention of antepartum condition
C0156839|T047|AB|648.12|ICD9CM|Thyroid dysfun-del w p/p|Thyroid dysfun-del w p/p
C0156839|T047|PT|648.12|ICD9CM|Thyroid dysfunction of mother, delivered, with mention of postpartum complication|Thyroid dysfunction of mother, delivered, with mention of postpartum complication
C0747834|T047|AB|648.13|ICD9CM|Thyroid dysfunc-antepart|Thyroid dysfunc-antepart
C0747834|T047|PT|648.13|ICD9CM|Thyroid dysfunction of mother, antepartum condition or complication|Thyroid dysfunction of mother, antepartum condition or complication
C0156841|T047|AB|648.14|ICD9CM|Thyroid dysfunc-postpart|Thyroid dysfunc-postpart
C0156841|T047|PT|648.14|ICD9CM|Thyroid dysfunction of mother, postpartum condition or complication|Thyroid dysfunction of mother, postpartum condition or complication
C0269684|T047|HT|648.2|ICD9CM|Anemia complicating pregnancy, childbirth, or the puerperium|Anemia complicating pregnancy, childbirth, or the puerperium
C0269684|T047|AB|648.20|ICD9CM|Anemia in preg-unspec|Anemia in preg-unspec
C0269684|T047|PT|648.20|ICD9CM|Anemia of mother, unspecified as to episode of care or not applicable|Anemia of mother, unspecified as to episode of care or not applicable
C0156844|T047|PT|648.21|ICD9CM|Anemia of mother, delivered, with or without mention of antepartum condition|Anemia of mother, delivered, with or without mention of antepartum condition
C0156844|T047|AB|648.21|ICD9CM|Anemia-delivered|Anemia-delivered
C0156845|T047|PT|648.22|ICD9CM|Anemia of mother, delivered, with mention of postpartum complication|Anemia of mother, delivered, with mention of postpartum complication
C0156845|T047|AB|648.22|ICD9CM|Anemia-delivered w p/p|Anemia-delivered w p/p
C0271930|T047|PT|648.23|ICD9CM|Anemia of mother, antepartum condition or complication|Anemia of mother, antepartum condition or complication
C0271930|T047|AB|648.23|ICD9CM|Anemia-antepartum|Anemia-antepartum
C0156847|T047|PT|648.24|ICD9CM|Anemia of mother, postpartum condition or complication|Anemia of mother, postpartum condition or complication
C0156847|T047|AB|648.24|ICD9CM|Anemia-postpartum|Anemia-postpartum
C0269685|T048|HT|648.3|ICD9CM|Drug dependence complicating pregnancy, childbirth, or the puerperium|Drug dependence complicating pregnancy, childbirth, or the puerperium
C0269685|T048|AB|648.30|ICD9CM|Drug depend preg-unspec|Drug depend preg-unspec
C0269685|T048|PT|648.30|ICD9CM|Drug dependence of mother, unspecified as to episode of care or not applicable|Drug dependence of mother, unspecified as to episode of care or not applicable
C0156850|T048|PT|648.31|ICD9CM|Drug dependence of mother, delivered, with or without mention of antepartum condition|Drug dependence of mother, delivered, with or without mention of antepartum condition
C0156850|T048|AB|648.31|ICD9CM|Drug dependence-deliver|Drug dependence-deliver
C0156851|T048|AB|648.32|ICD9CM|Drug dependen-del w p/p|Drug dependen-del w p/p
C0156851|T048|PT|648.32|ICD9CM|Drug dependence of mother, delivered, with mention of postpartum complication|Drug dependence of mother, delivered, with mention of postpartum complication
C0156852|T048|PT|648.33|ICD9CM|Drug dependence of mother, antepartum condition or complication|Drug dependence of mother, antepartum condition or complication
C0156852|T048|AB|648.33|ICD9CM|Drug dependence-antepart|Drug dependence-antepart
C0156853|T048|PT|648.34|ICD9CM|Drug dependence of mother, postpartum condition or complication|Drug dependence of mother, postpartum condition or complication
C0156853|T048|AB|648.34|ICD9CM|Drug dependence-postpart|Drug dependence-postpart
C0156854|T048|HT|648.4|ICD9CM|Mental disorders complicating pregnancy, childbirth, or the puerperium|Mental disorders complicating pregnancy, childbirth, or the puerperium
C0156855|T048|AB|648.40|ICD9CM|Mental dis preg-unspec|Mental dis preg-unspec
C0156855|T048|PT|648.40|ICD9CM|Mental disorders of mother, unspecified as to episode of care or not applicable|Mental disorders of mother, unspecified as to episode of care or not applicable
C0156856|T048|AB|648.41|ICD9CM|Mental disorder-deliver|Mental disorder-deliver
C0156856|T048|PT|648.41|ICD9CM|Mental disorders of mother, delivered, with or without mention of antepartum condition|Mental disorders of mother, delivered, with or without mention of antepartum condition
C0156857|T048|AB|648.42|ICD9CM|Mental dis-deliv w p/p|Mental dis-deliv w p/p
C0156857|T048|PT|648.42|ICD9CM|Mental disorders of mother, delivered, with mention of postpartum complication|Mental disorders of mother, delivered, with mention of postpartum complication
C0156858|T048|AB|648.43|ICD9CM|Mental disorder-antepart|Mental disorder-antepart
C0156858|T048|PT|648.43|ICD9CM|Mental disorders of mother, antepartum condition or complication|Mental disorders of mother, antepartum condition or complication
C0156859|T048|AB|648.44|ICD9CM|Mental disorder-postpart|Mental disorder-postpart
C0156859|T048|PT|648.44|ICD9CM|Mental disorders of mother, postpartum condition or complication|Mental disorders of mother, postpartum condition or complication
C0156860|T047|HT|648.5|ICD9CM|Congenital cardiovascular disorders complicating pregnancy, childbirth, or the puerperium|Congenital cardiovascular disorders complicating pregnancy, childbirth, or the puerperium
C0156861|T047|AB|648.50|ICD9CM|Congen CV dis preg-unsp|Congen CV dis preg-unsp
C0156861|T047|PT|648.50|ICD9CM|Congenital cardiovascular disorders of mother, unspecified as to episode of care or not applicable|Congenital cardiovascular disorders of mother, unspecified as to episode of care or not applicable
C0156862|T047|AB|648.51|ICD9CM|Congen CV dis-delivered|Congen CV dis-delivered
C0156863|T047|AB|648.52|ICD9CM|Congen CV dis-del w p/p|Congen CV dis-del w p/p
C0156863|T047|PT|648.52|ICD9CM|Congenital cardiovascular disorders of mother, delivered, with mention of postpartum complication|Congenital cardiovascular disorders of mother, delivered, with mention of postpartum complication
C0156864|T047|AB|648.53|ICD9CM|Congen CV dis-antepartum|Congen CV dis-antepartum
C0156864|T047|PT|648.53|ICD9CM|Congenital cardiovascular disorders of mother, antepartum condition or complication|Congenital cardiovascular disorders of mother, antepartum condition or complication
C0156865|T047|AB|648.54|ICD9CM|Congen CV dis-postpartum|Congen CV dis-postpartum
C0156865|T047|PT|648.54|ICD9CM|Congenital cardiovascular disorders of mother, postpartum condition or complication|Congenital cardiovascular disorders of mother, postpartum condition or complication
C0156866|T047|HT|648.6|ICD9CM|Other cardiovascular diseases complicating pregnancy, childbirth, or the puerperium|Other cardiovascular diseases complicating pregnancy, childbirth, or the puerperium
C0156867|T047|AB|648.60|ICD9CM|CV dis NEC preg-unspec|CV dis NEC preg-unspec
C0156867|T047|PT|648.60|ICD9CM|Other cardiovascular diseases of mother, unspecified as to episode of care or not applicable|Other cardiovascular diseases of mother, unspecified as to episode of care or not applicable
C0156868|T047|AB|648.61|ICD9CM|CV dis NEC preg-deliver|CV dis NEC preg-deliver
C0156868|T047|PT|648.61|ICD9CM|Other cardiovascular diseases of mother, delivered, with or without mention of antepartum condition|Other cardiovascular diseases of mother, delivered, with or without mention of antepartum condition
C0156869|T047|AB|648.62|ICD9CM|CV dis NEC-deliver w p/p|CV dis NEC-deliver w p/p
C0156869|T047|PT|648.62|ICD9CM|Other cardiovascular diseases of mother, delivered, with mention of postpartum complication|Other cardiovascular diseases of mother, delivered, with mention of postpartum complication
C0156870|T047|AB|648.63|ICD9CM|CV dis NEC-antepartum|CV dis NEC-antepartum
C0156870|T047|PT|648.63|ICD9CM|Other cardiovascular diseases of mother, antepartum condition or complication|Other cardiovascular diseases of mother, antepartum condition or complication
C0156871|T047|AB|648.64|ICD9CM|CV dis NEC-postpartum|CV dis NEC-postpartum
C0156871|T047|PT|648.64|ICD9CM|Other cardiovascular diseases of mother, postpartum condition or complication|Other cardiovascular diseases of mother, postpartum condition or complication
C0156873|T047|AB|648.70|ICD9CM|Bone disord in preg-unsp|Bone disord in preg-unsp
C0156874|T047|AB|648.71|ICD9CM|Bone disorder-delivered|Bone disorder-delivered
C0156875|T047|AB|648.72|ICD9CM|Bone disorder-del w p/p|Bone disorder-del w p/p
C0156876|T047|AB|648.73|ICD9CM|Bone disorder-antepartum|Bone disorder-antepartum
C0156877|T047|AB|648.74|ICD9CM|Bone disorder-postpartum|Bone disorder-postpartum
C0156878|T047|HT|648.8|ICD9CM|Abnormal glucose tolerance of mother, complicating pregnancy, childbirth, or the puerperium|Abnormal glucose tolerance of mother, complicating pregnancy, childbirth, or the puerperium
C0156879|T047|AB|648.80|ICD9CM|Abn glucose in preg-unsp|Abn glucose in preg-unsp
C0156879|T047|PT|648.80|ICD9CM|Abnormal glucose tolerance of mother, unspecified as to episode of care or not applicable|Abnormal glucose tolerance of mother, unspecified as to episode of care or not applicable
C0156880|T047|AB|648.81|ICD9CM|Abn glucose toler-deliv|Abn glucose toler-deliv
C0156880|T047|PT|648.81|ICD9CM|Abnormal glucose tolerance of mother, delivered, with or without mention of antepartum condition|Abnormal glucose tolerance of mother, delivered, with or without mention of antepartum condition
C0156881|T046|AB|648.82|ICD9CM|Abn glucose-deliv w p/p|Abn glucose-deliv w p/p
C0156881|T046|PT|648.82|ICD9CM|Abnormal glucose tolerance of mother, delivered, with mention of postpartum complication|Abnormal glucose tolerance of mother, delivered, with mention of postpartum complication
C0156882|T047|AB|648.83|ICD9CM|Abn glucose-antepartum|Abn glucose-antepartum
C0156882|T047|PT|648.83|ICD9CM|Abnormal glucose tolerance of mother, antepartum condition or complication|Abnormal glucose tolerance of mother, antepartum condition or complication
C0156883|T047|AB|648.84|ICD9CM|Abn glucose-postpartum|Abn glucose-postpartum
C0156883|T047|PT|648.84|ICD9CM|Abnormal glucose tolerance of mother, postpartum condition or complication|Abnormal glucose tolerance of mother, postpartum condition or complication
C0156884|T047|HT|648.9|ICD9CM|Other current conditions complicating pregnancy, childbirth, or the puerperium|Other current conditions complicating pregnancy, childbirth, or the puerperium
C0156885|T047|AB|648.90|ICD9CM|Oth curr cond preg-unsp|Oth curr cond preg-unsp
C0156886|T047|AB|648.91|ICD9CM|Oth curr cond-delivered|Oth curr cond-delivered
C0156887|T047|AB|648.92|ICD9CM|Oth curr cond-del w p/p|Oth curr cond-del w p/p
C0156888|T047|AB|648.93|ICD9CM|Oth curr cond-antepartum|Oth curr cond-antepartum
C0156888|T047|PT|648.93|ICD9CM|Other current conditions classifiable elsewhere of mother, antepartum condition or complication|Other current conditions classifiable elsewhere of mother, antepartum condition or complication
C0156889|T047|AB|648.94|ICD9CM|Oth curr cond-postpartum|Oth curr cond-postpartum
C0156889|T047|PT|648.94|ICD9CM|Other current conditions classifiable elsewhere of mother, postpartum condition or complication|Other current conditions classifiable elsewhere of mother, postpartum condition or complication
C1719602|T047|HT|649|ICD9CM|Other conditions or status of the mother complicating pregnancy, childbirth, or the puerperium|Other conditions or status of the mother complicating pregnancy, childbirth, or the puerperium
C1719563|T047|HT|649.0|ICD9CM|Tobacco use disorder complicating pregnancy, childbirth, or the puerperium|Tobacco use disorder complicating pregnancy, childbirth, or the puerperium
C1719558|T047|AB|649.00|ICD9CM|Tobacco use disord-unsp|Tobacco use disord-unsp
C1719559|T047|AB|649.01|ICD9CM|Tobacco use disor-delliv|Tobacco use disor-delliv
C1719560|T047|AB|649.02|ICD9CM|Tobacco use dis-del-p/p|Tobacco use dis-del-p/p
C1719561|T047|AB|649.03|ICD9CM|Tobacco use dis-antepart|Tobacco use dis-antepart
C1719562|T047|AB|649.04|ICD9CM|Tobacco use dis-postpart|Tobacco use dis-postpart
C1719570|T047|HT|649.1|ICD9CM|Obesity complicating pregnancy, childbirth, or the puerperium|Obesity complicating pregnancy, childbirth, or the puerperium
C1719565|T047|AB|649.10|ICD9CM|Obesity-unspecified|Obesity-unspecified
C1719566|T047|AB|649.11|ICD9CM|Obesity-delivered|Obesity-delivered
C1719567|T047|AB|649.12|ICD9CM|Obesity-delivered w p/p|Obesity-delivered w p/p
C1719568|T047|PT|649.13|ICD9CM|Obesity complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication|Obesity complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C1719568|T047|AB|649.13|ICD9CM|Obesity-antepartum|Obesity-antepartum
C1719569|T047|PT|649.14|ICD9CM|Obesity complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication|Obesity complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication
C1719569|T047|AB|649.14|ICD9CM|Obesity-postpartum|Obesity-postpartum
C1719576|T046|HT|649.2|ICD9CM|Bariatric surgery status complicating pregnancy, childbirth, or the puerperium|Bariatric surgery status complicating pregnancy, childbirth, or the puerperium
C1719571|T033|AB|649.20|ICD9CM|Bariatric surg stat-unsp|Bariatric surg stat-unsp
C1719572|T033|AB|649.21|ICD9CM|Bariatric surg stat-del|Bariatric surg stat-del
C1719573|T033|AB|649.22|ICD9CM|Bariatric surg-del w p/p|Bariatric surg-del w p/p
C1719574|T033|AB|649.23|ICD9CM|Bariatrc surg stat-antep|Bariatrc surg stat-antep
C1719575|T033|AB|649.24|ICD9CM|Bariatrc surg stat w p/p|Bariatrc surg stat w p/p
C1719585|T047|HT|649.3|ICD9CM|Coagulation defects complicating pregnancy, childbirth, or the puerperium|Coagulation defects complicating pregnancy, childbirth, or the puerperium
C1719580|T047|AB|649.30|ICD9CM|Coagulation def-unspec|Coagulation def-unspec
C1719581|T047|AB|649.31|ICD9CM|Coagulation def-deliv|Coagulation def-deliv
C1719582|T047|AB|649.32|ICD9CM|Coagulatn def-del w p/p|Coagulatn def-del w p/p
C1719583|T047|AB|649.33|ICD9CM|Coagulation def-antepart|Coagulation def-antepart
C1719584|T047|AB|649.34|ICD9CM|Coagulation def-postpart|Coagulation def-postpart
C1719591|T047|HT|649.4|ICD9CM|Epilepsy complicating pregnancy, childbirth, or the puerperium|Epilepsy complicating pregnancy, childbirth, or the puerperium
C1719586|T047|AB|649.40|ICD9CM|Epilepsy-unspecified|Epilepsy-unspecified
C1719587|T047|AB|649.41|ICD9CM|Epilepsy-delivered|Epilepsy-delivered
C1719588|T047|AB|649.42|ICD9CM|Epilepsy-delivered w p/p|Epilepsy-delivered w p/p
C1719589|T047|PT|649.43|ICD9CM|Epilepsy complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication|Epilepsy complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C1719589|T047|AB|649.43|ICD9CM|Epilepsy-antepartum|Epilepsy-antepartum
C1719590|T047|PT|649.44|ICD9CM|Epilepsy complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication|Epilepsy complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication
C1719590|T047|AB|649.44|ICD9CM|Epilepsy-postpartum|Epilepsy-postpartum
C1719595|T046|HT|649.5|ICD9CM|Spotting complicating pregnancy|Spotting complicating pregnancy
C1719592|T047|PT|649.50|ICD9CM|Spotting complicating pregnancy, unspecified as to episode of care or not applicable|Spotting complicating pregnancy, unspecified as to episode of care or not applicable
C1719592|T047|AB|649.50|ICD9CM|Spotting-unspecified|Spotting-unspecified
C1719593|T047|PT|649.51|ICD9CM|Spotting complicating pregnancy, delivered, with or without mention of antepartum condition|Spotting complicating pregnancy, delivered, with or without mention of antepartum condition
C1719593|T047|AB|649.51|ICD9CM|Spotting-delivered|Spotting-delivered
C1719594|T047|PT|649.53|ICD9CM|Spotting complicating pregnancy, antepartum condition or complication|Spotting complicating pregnancy, antepartum condition or complication
C1719594|T047|AB|649.53|ICD9CM|Spotting-antepartum|Spotting-antepartum
C1719601|T033|HT|649.6|ICD9CM|Uterine size date discrepancy|Uterine size date discrepancy
C1719596|T033|PT|649.60|ICD9CM|Uterine size date discrepancy, unspecified as to episode of care or not applicable|Uterine size date discrepancy, unspecified as to episode of care or not applicable
C1719596|T033|AB|649.60|ICD9CM|Uterine size descrp-unsp|Uterine size descrp-unsp
C1719597|T033|PT|649.61|ICD9CM|Uterine size date discrepancy, delivered, with or without mention of antepartum condition|Uterine size date discrepancy, delivered, with or without mention of antepartum condition
C1719597|T033|AB|649.61|ICD9CM|Uterine size descrep-del|Uterine size descrep-del
C1719598|T033|PT|649.62|ICD9CM|Uterine size date discrepancy, delivered, with mention of postpartum complication|Uterine size date discrepancy, delivered, with mention of postpartum complication
C1719598|T033|AB|649.62|ICD9CM|Uterine size-del w p/p|Uterine size-del w p/p
C1719599|T033|PT|649.63|ICD9CM|Uterine size date discrepancy, antepartum condition or complication|Uterine size date discrepancy, antepartum condition or complication
C1719599|T033|AB|649.63|ICD9CM|Uterine size des-antepar|Uterine size des-antepar
C1719600|T033|PT|649.64|ICD9CM|Uterine size date discrepancy, postpartum condition or complication|Uterine size date discrepancy, postpartum condition or complication
C1719600|T033|AB|649.64|ICD9CM|Uterine size descrep-p/p|Uterine size descrep-p/p
C2349587|T046|HT|649.7|ICD9CM|Cervical shortening|Cervical shortening
C2349584|T046|AB|649.70|ICD9CM|Cervical shortening-unsp|Cervical shortening-unsp
C2349584|T046|PT|649.70|ICD9CM|Cervical shortening, unspecified as to episode of care or not applicable|Cervical shortening, unspecified as to episode of care or not applicable
C2349585|T046|AB|649.71|ICD9CM|Cervical shortening-del|Cervical shortening-del
C2349585|T046|PT|649.71|ICD9CM|Cervical shortening, delivered, with or without mention of antepartum condition|Cervical shortening, delivered, with or without mention of antepartum condition
C2349586|T046|AB|649.73|ICD9CM|Cervical shortening-ante|Cervical shortening-ante
C2349586|T046|PT|649.73|ICD9CM|Cervical shortening, antepartum condition or complication|Cervical shortening, antepartum condition or complication
C3161121|T033|AB|649.81|ICD9CM|Spon labr w plan C/S-del|Spon labr w plan C/S-del
C3161122|T033|AB|649.82|ICD9CM|Lbr w plan C/S-del w p/p|Lbr w plan C/S-del w p/p
C1384485|T033|AB|650|ICD9CM|Normal delivery|Normal delivery
C1384485|T033|PT|650|ICD9CM|Normal delivery|Normal delivery
C0032989|T033|HT|651|ICD9CM|Multiple gestation|Multiple gestation
C0152150|T033|HT|651.0|ICD9CM|Twin pregnancy|Twin pregnancy
C0156893|T033|AB|651.01|ICD9CM|Twin pregnancy-delivered|Twin pregnancy-delivered
C0156893|T033|PT|651.01|ICD9CM|Twin pregnancy, delivered, with or without mention of antepartum condition|Twin pregnancy, delivered, with or without mention of antepartum condition
C0156894|T047|AB|651.03|ICD9CM|Twin pregnancy-antepart|Twin pregnancy-antepart
C0156894|T047|PT|651.03|ICD9CM|Twin pregnancy, antepartum condition or complication|Twin pregnancy, antepartum condition or complication
C0152151|T046|HT|651.1|ICD9CM|Triplet pregnancy|Triplet pregnancy
C0156896|T033|AB|651.11|ICD9CM|Triplet pregnancy-deliv|Triplet pregnancy-deliv
C0156896|T033|PT|651.11|ICD9CM|Triplet pregnancy, delivered, with or without mention of antepartum condition|Triplet pregnancy, delivered, with or without mention of antepartum condition
C0156897|T047|AB|651.13|ICD9CM|Triplet preg-antepartum|Triplet preg-antepartum
C0156897|T047|PT|651.13|ICD9CM|Triplet pregnancy, antepartum condition or complication|Triplet pregnancy, antepartum condition or complication
C0152152|T046|HT|651.2|ICD9CM|Quadruplet pregnancy|Quadruplet pregnancy
C0156899|T033|AB|651.21|ICD9CM|Quadruplet preg-deliver|Quadruplet preg-deliver
C0156899|T033|PT|651.21|ICD9CM|Quadruplet pregnancy, delivered, with or without mention of antepartum condition|Quadruplet pregnancy, delivered, with or without mention of antepartum condition
C0156900|T047|AB|651.23|ICD9CM|Quadruplet preg-antepart|Quadruplet preg-antepart
C0156900|T047|PT|651.23|ICD9CM|Quadruplet pregnancy, antepartum condition or complication|Quadruplet pregnancy, antepartum condition or complication
C0156901|T046|HT|651.3|ICD9CM|Twin pregnancy with fetal loss and retention of one fetus|Twin pregnancy with fetal loss and retention of one fetus
C0156902|T047|AB|651.30|ICD9CM|Twins w fetal loss-unsp|Twins w fetal loss-unsp
C0156903|T047|AB|651.31|ICD9CM|Twins w fetal loss-del|Twins w fetal loss-del
C0156904|T047|PT|651.33|ICD9CM|Twin pregnancy with fetal loss and retention of one fetus, antepartum condition or complication|Twin pregnancy with fetal loss and retention of one fetus, antepartum condition or complication
C0156904|T047|AB|651.33|ICD9CM|Twins w fetal loss-ante|Twins w fetal loss-ante
C0156905|T046|HT|651.4|ICD9CM|Triplet pregnancy with fetal loss and retention of one or more fetus (es)|Triplet pregnancy with fetal loss and retention of one or more fetus (es)
C0156906|T047|AB|651.40|ICD9CM|Triplets w fet loss-unsp|Triplets w fet loss-unsp
C0156907|T047|AB|651.41|ICD9CM|Triplets w fet loss-del|Triplets w fet loss-del
C0156908|T047|AB|651.43|ICD9CM|Triplets w fet loss-ante|Triplets w fet loss-ante
C0156909|T046|HT|651.5|ICD9CM|Quadruplet pregnancy with fetal loss and retention of one or more fetus(es)|Quadruplet pregnancy with fetal loss and retention of one or more fetus(es)
C0156910|T047|AB|651.50|ICD9CM|Quads w fetal loss-unsp|Quads w fetal loss-unsp
C0156911|T047|AB|651.51|ICD9CM|Quads w fetal loss-del|Quads w fetal loss-del
C0156912|T047|AB|651.53|ICD9CM|Quads w fetal loss-ante|Quads w fetal loss-ante
C0156913|T047|HT|651.6|ICD9CM|Other multiple pregnancy with fetal loss and retention of one or more fetus(es)|Other multiple pregnancy with fetal loss and retention of one or more fetus(es)
C0156914|T047|AB|651.60|ICD9CM|Mult ges w fet loss-unsp|Mult ges w fet loss-unsp
C0156915|T047|AB|651.61|ICD9CM|Mult ges w fet loss-del|Mult ges w fet loss-del
C0156916|T047|AB|651.63|ICD9CM|Mult ges w fet loss-ante|Mult ges w fet loss-ante
C1561650|T033|HT|651.7|ICD9CM|Multiple gestation following (elective) fetal reduction|Multiple gestation following (elective) fetal reduction
C1561647|T033|AB|651.70|ICD9CM|Mul gest-fet reduct unsp|Mul gest-fet reduct unsp
C1561648|T033|AB|651.71|ICD9CM|Mult gest-fet reduct del|Mult gest-fet reduct del
C1561649|T033|AB|651.73|ICD9CM|Mul gest-fet reduct ante|Mul gest-fet reduct ante
C1561649|T033|PT|651.73|ICD9CM|Multiple gestation following (elective) fetal reduction, antepartum condition or complication|Multiple gestation following (elective) fetal reduction, antepartum condition or complication
C0156917|T033|HT|651.8|ICD9CM|Other specified multiple gestation|Other specified multiple gestation
C0032989|T033|HT|651.9|ICD9CM|Unspecified multiple gestation|Unspecified multiple gestation
C0032989|T033|AB|651.90|ICD9CM|Multi gestat NOS-unspec|Multi gestat NOS-unspec
C0032989|T033|PT|651.90|ICD9CM|Unspecified multiple gestation, unspecified as to episode of care or not applicable|Unspecified multiple gestation, unspecified as to episode of care or not applicable
C0156923|T046|AB|651.93|ICD9CM|Multi gest NOS-antepart|Multi gest NOS-antepart
C0156923|T046|PT|651.93|ICD9CM|Unspecified multiple gestation, antepartum condition or complication|Unspecified multiple gestation, antepartum condition or complication
C0156924|T033|HT|652|ICD9CM|Malposition and malpresentation of fetus|Malposition and malpresentation of fetus
C0426066|T033|HT|652.0|ICD9CM|Unstable lie of fetus|Unstable lie of fetus
C0156926|T047|AB|652.00|ICD9CM|Unstable lie-unspecified|Unstable lie-unspecified
C0156926|T047|PT|652.00|ICD9CM|Unstable lie, unspecified as to episode of care or not applicable|Unstable lie, unspecified as to episode of care or not applicable
C0156927|T033|AB|652.01|ICD9CM|Unstable lie-delivered|Unstable lie-delivered
C0156927|T033|PT|652.01|ICD9CM|Unstable lie, delivered, with or without mention of antepartum condition|Unstable lie, delivered, with or without mention of antepartum condition
C0156928|T047|AB|652.03|ICD9CM|Unstable lie-antepartum|Unstable lie-antepartum
C0156928|T047|PT|652.03|ICD9CM|Unstable lie, antepartum condition or complication|Unstable lie, antepartum condition or complication
C0156929|T047|HT|652.1|ICD9CM|Breech or other malpresentation successfully converted to cephalic presentation|Breech or other malpresentation successfully converted to cephalic presentation
C0156930|T047|AB|652.10|ICD9CM|Cephalic vers NOS-unspec|Cephalic vers NOS-unspec
C0156931|T047|AB|652.11|ICD9CM|Cephalic vers NOS-deliv|Cephalic vers NOS-deliv
C0156932|T047|AB|652.13|ICD9CM|Cephal vers NOS-antepart|Cephal vers NOS-antepart
C0156933|T047|AB|652.20|ICD9CM|Breech presentat-unspec|Breech presentat-unspec
C0156933|T047|PT|652.20|ICD9CM|Breech presentation without mention of version, unspecified as to episode of care or not applicable|Breech presentation without mention of version, unspecified as to episode of care or not applicable
C0156934|T047|AB|652.21|ICD9CM|Breech presentat-deliver|Breech presentat-deliver
C0156935|T047|AB|652.23|ICD9CM|Breech present-antepart|Breech present-antepart
C0156935|T047|PT|652.23|ICD9CM|Breech presentation without mention of version, antepartum condition or complication|Breech presentation without mention of version, antepartum condition or complication
C0156936|T033|HT|652.3|ICD9CM|Transverse or oblique presentation of fetus|Transverse or oblique presentation of fetus
C0375391|T033|AB|652.30|ICD9CM|Transv/obliq lie-unspec|Transv/obliq lie-unspec
C0375391|T033|PT|652.30|ICD9CM|Transverse or oblique presentation, unspecified as to episode of care or not applicable|Transverse or oblique presentation, unspecified as to episode of care or not applicable
C0375392|T033|AB|652.31|ICD9CM|Transver/obliq lie-deliv|Transver/obliq lie-deliv
C0375392|T033|PT|652.31|ICD9CM|Transverse or oblique presentation, delivered, with or without mention of antepartum condition|Transverse or oblique presentation, delivered, with or without mention of antepartum condition
C0375393|T033|AB|652.33|ICD9CM|Transv/obliq lie-antepar|Transv/obliq lie-antepar
C0375393|T033|PT|652.33|ICD9CM|Transverse or oblique presentation, antepartum condition or complication|Transverse or oblique presentation, antepartum condition or complication
C0156940|T033|HT|652.4|ICD9CM|Face or brow presentation of fetus|Face or brow presentation of fetus
C0156941|T033|PT|652.40|ICD9CM|Face or brow presentation, unspecified as to episode of care or not applicable|Face or brow presentation, unspecified as to episode of care or not applicable
C0156941|T033|AB|652.40|ICD9CM|Face/brow present-unspec|Face/brow present-unspec
C0156942|T033|PT|652.41|ICD9CM|Face or brow presentation, delivered, with or without mention of antepartum condition|Face or brow presentation, delivered, with or without mention of antepartum condition
C0156942|T033|AB|652.41|ICD9CM|Face/brow present-deliv|Face/brow present-deliv
C0156943|T033|PT|652.43|ICD9CM|Face or brow presentation, antepartum condition or complication|Face or brow presentation, antepartum condition or complication
C0156943|T033|AB|652.43|ICD9CM|Face/brow pres-antepart|Face/brow pres-antepart
C0426187|T033|HT|652.5|ICD9CM|High fetal head at term|High fetal head at term
C0156945|T047|AB|652.50|ICD9CM|High head at term-unspec|High head at term-unspec
C0156945|T047|PT|652.50|ICD9CM|High head at term, unspecified as to episode of care or not applicable|High head at term, unspecified as to episode of care or not applicable
C0156946|T033|AB|652.51|ICD9CM|High head at term-deliv|High head at term-deliv
C0156946|T033|PT|652.51|ICD9CM|High head at term, delivered, with or without mention of antepartum condition|High head at term, delivered, with or without mention of antepartum condition
C0156947|T047|PT|652.53|ICD9CM|High head at term, antepartum condition or complication|High head at term, antepartum condition or complication
C0156947|T047|AB|652.53|ICD9CM|High head term-antepart|High head term-antepart
C0156948|T047|HT|652.6|ICD9CM|Multiple gestation with malpresentation of one fetus or more|Multiple gestation with malpresentation of one fetus or more
C0156949|T047|AB|652.60|ICD9CM|Mult gest malpresen-unsp|Mult gest malpresen-unsp
C0156950|T047|AB|652.61|ICD9CM|Mult gest malpres-deliv|Mult gest malpres-deliv
C0156951|T047|AB|652.63|ICD9CM|Mult ges malpres-antepar|Mult ges malpres-antepar
C0156951|T047|PT|652.63|ICD9CM|Multiple gestation with malpresentation of one fetus or more, antepartum condtion or complication|Multiple gestation with malpresentation of one fetus or more, antepartum condtion or complication
C0269709|T046|HT|652.7|ICD9CM|Prolapsed arm of fetus|Prolapsed arm of fetus
C0156953|T047|PT|652.70|ICD9CM|Prolapsed arm of fetus, unspecified as to episode of care or not applicable|Prolapsed arm of fetus, unspecified as to episode of care or not applicable
C0156953|T047|AB|652.70|ICD9CM|Prolapsed arm-unspec|Prolapsed arm-unspec
C0156954|T047|PT|652.71|ICD9CM|Prolapsed arm of fetus, delivered, with or without mention of antepartum condition|Prolapsed arm of fetus, delivered, with or without mention of antepartum condition
C0156954|T047|AB|652.71|ICD9CM|Prolapsed arm-delivered|Prolapsed arm-delivered
C0156955|T047|PT|652.73|ICD9CM|Prolapsed arm of fetus, antepartum condition or complication|Prolapsed arm of fetus, antepartum condition or complication
C0156955|T047|AB|652.73|ICD9CM|Prolapsed arm-antepart|Prolapsed arm-antepart
C0156956|T047|HT|652.8|ICD9CM|Other specified malposition or malpresentation of fetus|Other specified malposition or malpresentation of fetus
C0156957|T047|AB|652.80|ICD9CM|Malposition NEC-unspec|Malposition NEC-unspec
C0156957|T047|PT|652.80|ICD9CM|Other specified malposition or malpresentation, unspecified as to episode of care or not applicable|Other specified malposition or malpresentation, unspecified as to episode of care or not applicable
C0156958|T047|AB|652.81|ICD9CM|Malposition NEC-deliver|Malposition NEC-deliver
C0156959|T047|AB|652.83|ICD9CM|Malposition NEC-antepart|Malposition NEC-antepart
C0156959|T047|PT|652.83|ICD9CM|Other specified malposition or malpresentation, antepartum condition or complication|Other specified malposition or malpresentation, antepartum condition or complication
C0156924|T033|HT|652.9|ICD9CM|Unspecified malposition or malpresentation of fetus|Unspecified malposition or malpresentation of fetus
C0156961|T047|AB|652.90|ICD9CM|Malposition NOS-unspec|Malposition NOS-unspec
C0156961|T047|PT|652.90|ICD9CM|Unspecified malposition or malpresentation, unspecified as to episode of care or not applicable|Unspecified malposition or malpresentation, unspecified as to episode of care or not applicable
C0156962|T047|AB|652.91|ICD9CM|Malposition NOS-deliver|Malposition NOS-deliver
C0156963|T047|AB|652.93|ICD9CM|Malposition NOS-antepart|Malposition NOS-antepart
C0156963|T047|PT|652.93|ICD9CM|Unspecified malposition or malpresentation, antepartum condition or complication|Unspecified malposition or malpresentation, antepartum condition or complication
C0156964|T046|HT|653|ICD9CM|Disproportion in pregnancy, labor, and delivery|Disproportion in pregnancy, labor, and delivery
C0269713|T046|HT|653.0|ICD9CM|Major abnormality of bony pelvis, not further specified, in pregnancy, labor, and delivery|Major abnormality of bony pelvis, not further specified, in pregnancy, labor, and delivery
C0156966|T020|AB|653.00|ICD9CM|Pelvic deform NOS-unspec|Pelvic deform NOS-unspec
C0156967|T020|AB|653.01|ICD9CM|Pelvic deform NOS-deliv|Pelvic deform NOS-deliv
C0156968|T020|PT|653.03|ICD9CM|Major abnormality of bony pelvis, not further specified, antepartum condition or complication|Major abnormality of bony pelvis, not further specified, antepartum condition or complication
C0156968|T020|AB|653.03|ICD9CM|Pelv deform NOS-antepart|Pelv deform NOS-antepart
C0156969|T020|HT|653.1|ICD9CM|Generally contracted pelvis in pregnancy, labor, and delivery|Generally contracted pelvis in pregnancy, labor, and delivery
C0156970|T020|AB|653.10|ICD9CM|Contract pelv NOS-unspec|Contract pelv NOS-unspec
C0156970|T020|PT|653.10|ICD9CM|Generally contracted pelvis, unspecified as to episode of care or not applicable|Generally contracted pelvis, unspecified as to episode of care or not applicable
C0156971|T033|AB|653.11|ICD9CM|Contract pelv NOS-deliv|Contract pelv NOS-deliv
C0156971|T033|PT|653.11|ICD9CM|Generally contracted pelvis, delivered, with or without mention of antepartum condition|Generally contracted pelvis, delivered, with or without mention of antepartum condition
C0156972|T020|AB|653.13|ICD9CM|Contrac pelv NOS-antepar|Contrac pelv NOS-antepar
C0156972|T020|PT|653.13|ICD9CM|Generally contracted pelvis, antepartum condition or complication|Generally contracted pelvis, antepartum condition or complication
C0156973|T020|HT|653.2|ICD9CM|Inlet contraction of pelvis in pregnancy, labor, and delivery|Inlet contraction of pelvis in pregnancy, labor, and delivery
C0156974|T020|PT|653.20|ICD9CM|Inlet contraction of pelvis, unspecified as to episode of care or not applicable|Inlet contraction of pelvis, unspecified as to episode of care or not applicable
C0156974|T020|AB|653.20|ICD9CM|Inlet contraction-unspec|Inlet contraction-unspec
C0156975|T190|PT|653.21|ICD9CM|Inlet contraction of pelvis, delivered, with or without mention of antepartum condition|Inlet contraction of pelvis, delivered, with or without mention of antepartum condition
C0156975|T190|AB|653.21|ICD9CM|Inlet contraction-deliv|Inlet contraction-deliv
C0156976|T020|AB|653.23|ICD9CM|Inlet contract-antepart|Inlet contract-antepart
C0156976|T020|PT|653.23|ICD9CM|Inlet contraction of pelvis, antepartum condition or complication|Inlet contraction of pelvis, antepartum condition or complication
C0156977|T046|HT|653.3|ICD9CM|Outlet contraction of pelvis in pregnancy, labor, and delivery|Outlet contraction of pelvis in pregnancy, labor, and delivery
C0156978|T020|PT|653.30|ICD9CM|Outlet contraction of pelvis, unspecified as to episode of care or not applicable|Outlet contraction of pelvis, unspecified as to episode of care or not applicable
C0156978|T020|AB|653.30|ICD9CM|Outlet contraction-unsp|Outlet contraction-unsp
C0156979|T190|PT|653.31|ICD9CM|Outlet contraction of pelvis, delivered, with or without mention of antepartum condition|Outlet contraction of pelvis, delivered, with or without mention of antepartum condition
C0156979|T190|AB|653.31|ICD9CM|Outlet contraction-deliv|Outlet contraction-deliv
C0156980|T020|AB|653.33|ICD9CM|Outlet contract-antepart|Outlet contract-antepart
C0156980|T020|PT|653.33|ICD9CM|Outlet contraction of pelvis, antepartum condition or complication|Outlet contraction of pelvis, antepartum condition or complication
C0085988|T033|HT|653.4|ICD9CM|Fetopelvic disproportion|Fetopelvic disproportion
C1142293|T047|AB|653.40|ICD9CM|Fetopelv disprop-unspec|Fetopelv disprop-unspec
C1142293|T047|PT|653.40|ICD9CM|Fetopelvic disproportion, unspecified as to episode of care or not applicable|Fetopelvic disproportion, unspecified as to episode of care or not applicable
C0156982|T047|AB|653.41|ICD9CM|Fetopelv dispropor-deliv|Fetopelv dispropor-deliv
C0156982|T047|PT|653.41|ICD9CM|Fetopelvic disproportion, delivered, with or without mention of antepartum condition|Fetopelvic disproportion, delivered, with or without mention of antepartum condition
C1142292|T046|AB|653.43|ICD9CM|Fetopel disprop-antepart|Fetopel disprop-antepart
C1142292|T046|PT|653.43|ICD9CM|Fetopelvic disproportion, antepartum condition or complication|Fetopelvic disproportion, antepartum condition or complication
C0156984|T033|HT|653.5|ICD9CM|Unusually large fetus causing disproportion|Unusually large fetus causing disproportion
C0156985|T047|AB|653.50|ICD9CM|Fetal disprop NOS-unspec|Fetal disprop NOS-unspec
C0156985|T047|PT|653.50|ICD9CM|Unusually large fetus causing disproportion, unspecified as to episode of care or not applicable|Unusually large fetus causing disproportion, unspecified as to episode of care or not applicable
C0156986|T047|AB|653.51|ICD9CM|Fetal disprop NOS-deliv|Fetal disprop NOS-deliv
C0156987|T047|AB|653.53|ICD9CM|Fetal dispro NOS-antepar|Fetal dispro NOS-antepar
C0156987|T047|PT|653.53|ICD9CM|Unusually large fetus causing disproportion, antepartum condition or complication|Unusually large fetus causing disproportion, antepartum condition or complication
C0405012|T190|HT|653.6|ICD9CM|Hydrocephalic fetus causing disproportion|Hydrocephalic fetus causing disproportion
C0156989|T047|AB|653.60|ICD9CM|Hydrocephal fetus-unspec|Hydrocephal fetus-unspec
C0156989|T047|PT|653.60|ICD9CM|Hydrocephalic fetus causing disproportion, unspecified as to episode of care or not applicable|Hydrocephalic fetus causing disproportion, unspecified as to episode of care or not applicable
C0156990|T047|AB|653.61|ICD9CM|Hydroceph fetus-deliver|Hydroceph fetus-deliver
C0156991|T047|AB|653.63|ICD9CM|Hydroceph fetus-antepart|Hydroceph fetus-antepart
C0156991|T047|PT|653.63|ICD9CM|Hydrocephalic fetus causing disproportion, antepartum condition or complication|Hydrocephalic fetus causing disproportion, antepartum condition or complication
C0405011|T190|HT|653.7|ICD9CM|Other fetal abnormality causing disproportion|Other fetal abnormality causing disproportion
C0156993|T047|AB|653.70|ICD9CM|Oth abn fet disprop-unsp|Oth abn fet disprop-unsp
C0156993|T047|PT|653.70|ICD9CM|Other fetal abnormality causing disproportion, unspecified as to episode of care or not applicable|Other fetal abnormality causing disproportion, unspecified as to episode of care or not applicable
C0156994|T019|AB|653.71|ICD9CM|Oth abn fet dispro-deliv|Oth abn fet dispro-deliv
C0156995|T047|AB|653.73|ICD9CM|Oth abn fet dispro-antep|Oth abn fet dispro-antep
C0156995|T047|PT|653.73|ICD9CM|Other fetal abnormality causing disproportion, antepartum condition or complication|Other fetal abnormality causing disproportion, antepartum condition or complication
C0156996|T046|HT|653.8|ICD9CM|Disproportion of other origin in pregnancy, labor, and delivery|Disproportion of other origin in pregnancy, labor, and delivery
C0156997|T047|AB|653.80|ICD9CM|Disproportion NEC-unspec|Disproportion NEC-unspec
C0156997|T047|PT|653.80|ICD9CM|Disproportion of other origin, unspecified as to episode of care or not applicable|Disproportion of other origin, unspecified as to episode of care or not applicable
C0156998|T047|AB|653.81|ICD9CM|Disproportion NEC-deliv|Disproportion NEC-deliv
C0156998|T047|PT|653.81|ICD9CM|Disproportion of other origin, delivered, with or without mention of antepartum condition|Disproportion of other origin, delivered, with or without mention of antepartum condition
C0156999|T047|AB|653.83|ICD9CM|Dispropor NEC-antepartum|Dispropor NEC-antepartum
C0156999|T047|PT|653.83|ICD9CM|Disproportion of other origin, antepartum condition or complication|Disproportion of other origin, antepartum condition or complication
C0157000|T046|HT|653.9|ICD9CM|Unspecified disproportion in pregnancy, labor, and delivery|Unspecified disproportion in pregnancy, labor, and delivery
C0157001|T047|AB|653.90|ICD9CM|Disproportion NOS-unspec|Disproportion NOS-unspec
C0157001|T047|PT|653.90|ICD9CM|Unspecified disproportion, unspecified as to episode of care or not applicable|Unspecified disproportion, unspecified as to episode of care or not applicable
C0157002|T047|AB|653.91|ICD9CM|Disproportion NOS-deliv|Disproportion NOS-deliv
C0157002|T047|PT|653.91|ICD9CM|Unspecified disproportion, delivered, with or without mention of antepartum condition|Unspecified disproportion, delivered, with or without mention of antepartum condition
C0157003|T047|AB|653.93|ICD9CM|Dispropor NOS-antepartum|Dispropor NOS-antepartum
C0157003|T047|PT|653.93|ICD9CM|Unspecified disproportion, antepartum condition or complication|Unspecified disproportion, antepartum condition or complication
C0157005|T047|HT|654.0|ICD9CM|Congenital abnormalities of uterus complicating pregnancy, childbirth, or the puerperium|Congenital abnormalities of uterus complicating pregnancy, childbirth, or the puerperium
C0157006|T019|AB|654.00|ICD9CM|Cong abn uter preg-unsp|Cong abn uter preg-unsp
C0157006|T019|PT|654.00|ICD9CM|Congenital abnormalities of uterus, unspecified as to episode of care or not applicable|Congenital abnormalities of uterus, unspecified as to episode of care or not applicable
C0157007|T019|AB|654.01|ICD9CM|Congen abn uterus-deliv|Congen abn uterus-deliv
C0157007|T019|PT|654.01|ICD9CM|Congenital abnormalities of uterus, delivered, with or without mention of antepartum condition|Congenital abnormalities of uterus, delivered, with or without mention of antepartum condition
C0157008|T047|AB|654.02|ICD9CM|Cong abn uter-del w p/p|Cong abn uter-del w p/p
C0157008|T047|PT|654.02|ICD9CM|Congenital abnormalities of uterus, delivered, with mention of postpartum complication|Congenital abnormalities of uterus, delivered, with mention of postpartum complication
C0157009|T019|AB|654.03|ICD9CM|Congen abn uter-antepart|Congen abn uter-antepart
C0157009|T047|AB|654.03|ICD9CM|Congen abn uter-antepart|Congen abn uter-antepart
C0157009|T019|PT|654.03|ICD9CM|Congenital abnormalities of uterus, antepartum condition or complication|Congenital abnormalities of uterus, antepartum condition or complication
C0157009|T047|PT|654.03|ICD9CM|Congenital abnormalities of uterus, antepartum condition or complication|Congenital abnormalities of uterus, antepartum condition or complication
C0157010|T047|AB|654.04|ICD9CM|Congen abn uter-postpart|Congen abn uter-postpart
C0157010|T047|PT|654.04|ICD9CM|Congenital abnormalities of uterus, postpartum condition or complication|Congenital abnormalities of uterus, postpartum condition or complication
C0157011|T191|HT|654.1|ICD9CM|Tumors of body of uterus complicating pregnancy, childbirth, or the puerperium|Tumors of body of uterus complicating pregnancy, childbirth, or the puerperium
C0157012|T191|PT|654.10|ICD9CM|Tumors of body of uterus, unspecified as to episode of care or not applicable|Tumors of body of uterus, unspecified as to episode of care or not applicable
C0157012|T191|AB|654.10|ICD9CM|Uter tumor in preg-unsp|Uter tumor in preg-unsp
C0157013|T191|PT|654.11|ICD9CM|Tumors of body of uterus, delivered, with or without mention of antepartum condition|Tumors of body of uterus, delivered, with or without mention of antepartum condition
C0157013|T191|AB|654.11|ICD9CM|Uterine tumor-delivered|Uterine tumor-delivered
C0157014|T191|PT|654.12|ICD9CM|Tumors of body of uterus, delivered, with mention of postpartum complication|Tumors of body of uterus, delivered, with mention of postpartum complication
C0157014|T191|AB|654.12|ICD9CM|Uterine tumor-del w p/p|Uterine tumor-del w p/p
C0157015|T191|PT|654.13|ICD9CM|Tumors of body of uterus, antepartum condition or complication|Tumors of body of uterus, antepartum condition or complication
C0157015|T191|AB|654.13|ICD9CM|Uterine tumor-antepartum|Uterine tumor-antepartum
C0157016|T191|PT|654.14|ICD9CM|Tumors of body of uterus, postpartum condition or complication|Tumors of body of uterus, postpartum condition or complication
C0157016|T191|AB|654.14|ICD9CM|Uterine tumor-postpartum|Uterine tumor-postpartum
C0375394|T033|HT|654.2|ICD9CM|Previous cesarean section complicating pregnancy or childbirth|Previous cesarean section complicating pregnancy or childbirth
C0157018|T033|AB|654.20|ICD9CM|Prev c-delivery unspec|Prev c-delivery unspec
C0157018|T033|PT|654.20|ICD9CM|Previous cesarean delivery, unspecified as to episode of care or not applicable|Previous cesarean delivery, unspecified as to episode of care or not applicable
C0375395|T033|AB|654.21|ICD9CM|Prev c-delivery-delivrd|Prev c-delivery-delivrd
C0375395|T033|PT|654.21|ICD9CM|Previous cesarean delivery, delivered, with or without mention of antepartum condition|Previous cesarean delivery, delivered, with or without mention of antepartum condition
C0157020|T033|AB|654.23|ICD9CM|Prev c-delivery-antepart|Prev c-delivery-antepart
C0157020|T033|PT|654.23|ICD9CM|Previous cesarean delivery, antepartum condition or complication|Previous cesarean delivery, antepartum condition or complication
C0404709|T047|HT|654.3|ICD9CM|Retroverted and incarcerated gravid uterus|Retroverted and incarcerated gravid uterus
C0157022|T047|AB|654.30|ICD9CM|Retrovert uterus-unspec|Retrovert uterus-unspec
C0157022|T047|PT|654.30|ICD9CM|Retroverted and incarcerated gravid uterus, unspecified as to episode of care or not applicable|Retroverted and incarcerated gravid uterus, unspecified as to episode of care or not applicable
C0157023|T047|AB|654.31|ICD9CM|Retrovert uterus-deliver|Retrovert uterus-deliver
C0157023|T047|PT|654.31|ICD9CM|Retroverted and incarcerated gravid uterus, delivered, with mention of antepartum condition|Retroverted and incarcerated gravid uterus, delivered, with mention of antepartum condition
C0157024|T047|AB|654.32|ICD9CM|Retrovert uter-del w p/p|Retrovert uter-del w p/p
C0157024|T047|PT|654.32|ICD9CM|Retroverted and incarcerated gravid uterus, delivered, with mention of postpartum complication|Retroverted and incarcerated gravid uterus, delivered, with mention of postpartum complication
C0157025|T047|AB|654.33|ICD9CM|Retrovert uter-antepart|Retrovert uter-antepart
C0157025|T047|PT|654.33|ICD9CM|Retroverted and incarcerated gravid uterus, antepartum condition or complication|Retroverted and incarcerated gravid uterus, antepartum condition or complication
C0157026|T047|AB|654.34|ICD9CM|Retrovert uter-postpart|Retrovert uter-postpart
C0157026|T047|PT|654.34|ICD9CM|Retroverted and incarcerated gravid uterus, postpartum condition or complication|Retroverted and incarcerated gravid uterus, postpartum condition or complication
C0859820|T047|HT|654.4|ICD9CM|Other abnormalities in shape or position of gravid uterus and of neighboring structures|Other abnormalities in shape or position of gravid uterus and of neighboring structures
C0157028|T047|AB|654.40|ICD9CM|Abn grav uterus NEC-unsp|Abn grav uterus NEC-unsp
C0157029|T047|AB|654.41|ICD9CM|Abn uterus NEC-delivered|Abn uterus NEC-delivered
C0157030|T047|AB|654.42|ICD9CM|Abn uterus NEC-del w p/p|Abn uterus NEC-del w p/p
C0157031|T047|AB|654.43|ICD9CM|Abn uterus NEC-antepart|Abn uterus NEC-antepart
C0157032|T047|AB|654.44|ICD9CM|Abn uterus NEC-postpart|Abn uterus NEC-postpart
C0157033|T020|HT|654.5|ICD9CM|Cervical incompetence complicating pregnancy, childbirth, or the puerperium|Cervical incompetence complicating pregnancy, childbirth, or the puerperium
C0157034|T047|AB|654.50|ICD9CM|Cerv incompet preg-unsp|Cerv incompet preg-unsp
C0157034|T047|PT|654.50|ICD9CM|Cervical incompetence, unspecified as to episode of care or not applicable|Cervical incompetence, unspecified as to episode of care or not applicable
C0157035|T046|AB|654.51|ICD9CM|Cervical incompet-deliv|Cervical incompet-deliv
C0157035|T046|PT|654.51|ICD9CM|Cervical incompetence, delivered, with or without mention of antepartum condition|Cervical incompetence, delivered, with or without mention of antepartum condition
C0157036|T047|AB|654.52|ICD9CM|Cerv incompet-del w p/p|Cerv incompet-del w p/p
C0157036|T047|PT|654.52|ICD9CM|Cervical incompetence, delivered, with mention of postpartum complication|Cervical incompetence, delivered, with mention of postpartum complication
C0157037|T047|AB|654.53|ICD9CM|Cerv incompet-antepartum|Cerv incompet-antepartum
C0157037|T047|PT|654.53|ICD9CM|Cervical incompetence, antepartum condition or complication|Cervical incompetence, antepartum condition or complication
C0157038|T047|AB|654.54|ICD9CM|Cerv incompet-postpartum|Cerv incompet-postpartum
C0157038|T047|PT|654.54|ICD9CM|Cervical incompetence, postpartum condition or complication|Cervical incompetence, postpartum condition or complication
C0157040|T047|AB|654.60|ICD9CM|Abn cervix NEC preg-unsp|Abn cervix NEC preg-unsp
C0157041|T047|AB|654.61|ICD9CM|Abn cervix NEC-delivered|Abn cervix NEC-delivered
C0157042|T047|AB|654.62|ICD9CM|Abn cervix NEC-del w p/p|Abn cervix NEC-del w p/p
C0157043|T047|AB|654.63|ICD9CM|Abn cervix NEC-antepart|Abn cervix NEC-antepart
C0157043|T047|PT|654.63|ICD9CM|Other congenital or acquired abnormality of cervix, antepartum condition or complication|Other congenital or acquired abnormality of cervix, antepartum condition or complication
C0157044|T047|AB|654.64|ICD9CM|Abn cervix NEC-postpart|Abn cervix NEC-postpart
C0157044|T047|PT|654.64|ICD9CM|Other congenital or acquired abnormality of cervix, postpartum condition or complication|Other congenital or acquired abnormality of cervix, postpartum condition or complication
C0157045|T047|HT|654.7|ICD9CM|Congenital or acquired abnormality of vagina complicating pregnancy, childbirth, or the puerperium|Congenital or acquired abnormality of vagina complicating pregnancy, childbirth, or the puerperium
C0157046|T047|AB|654.70|ICD9CM|Abn vagina in preg-unsp|Abn vagina in preg-unsp
C0157046|T047|PT|654.70|ICD9CM|Congenital or acquired abnormality of vagina, unspecified as to episode of care or not applicable|Congenital or acquired abnormality of vagina, unspecified as to episode of care or not applicable
C0157047|T047|AB|654.71|ICD9CM|Abnorm vagina-delivered|Abnorm vagina-delivered
C0157048|T047|AB|654.72|ICD9CM|Abnorm vagina-del w p/p|Abnorm vagina-del w p/p
C0157048|T047|PT|654.72|ICD9CM|Congenital or acquired abnormality of vagina, delivered, with mention of postpartum complication|Congenital or acquired abnormality of vagina, delivered, with mention of postpartum complication
C0157049|T047|AB|654.73|ICD9CM|Abnorm vagina-antepartum|Abnorm vagina-antepartum
C0157049|T047|PT|654.73|ICD9CM|Congenital or acquired abnormality of vagina, antepartum condition or complication|Congenital or acquired abnormality of vagina, antepartum condition or complication
C0157050|T047|AB|654.74|ICD9CM|Abnorm vagina-postpartum|Abnorm vagina-postpartum
C0157050|T047|PT|654.74|ICD9CM|Congenital or acquired abnormality of vagina, postpartum condition or complication|Congenital or acquired abnormality of vagina, postpartum condition or complication
C0157051|T047|HT|654.8|ICD9CM|Congenital or acquired abnormality of vulva complicating pregnancy, childbirth, or the puerperium|Congenital or acquired abnormality of vulva complicating pregnancy, childbirth, or the puerperium
C0157052|T047|AB|654.80|ICD9CM|Abn vulva in preg-unspec|Abn vulva in preg-unspec
C0157052|T047|PT|654.80|ICD9CM|Congenital or acquired abnormality of vulva, unspecified as to episode of care or not applicable|Congenital or acquired abnormality of vulva, unspecified as to episode of care or not applicable
C0157053|T047|AB|654.81|ICD9CM|Abnormal vulva-delivered|Abnormal vulva-delivered
C0157054|T047|AB|654.82|ICD9CM|Abnormal vulva-del w p/p|Abnormal vulva-del w p/p
C0157054|T047|PT|654.82|ICD9CM|Congenital or acquired abnormality of vulva, delivered, with mention of postpartum complication|Congenital or acquired abnormality of vulva, delivered, with mention of postpartum complication
C0157055|T047|AB|654.83|ICD9CM|Abnormal vulva-antepart|Abnormal vulva-antepart
C0157055|T047|PT|654.83|ICD9CM|Congenital or acquired abnormality of vulva, antepartum condition or complication|Congenital or acquired abnormality of vulva, antepartum condition or complication
C0157056|T047|AB|654.84|ICD9CM|Abnormal vulva-postpart|Abnormal vulva-postpart
C0157056|T047|PT|654.84|ICD9CM|Congenital or acquired abnormality of vulva, postpartum condition or complication|Congenital or acquired abnormality of vulva, postpartum condition or complication
C0157058|T190|AB|654.90|ICD9CM|Abn pel NEC in preg-unsp|Abn pel NEC in preg-unsp
C0157059|T190|AB|654.91|ICD9CM|Abn pelv org NEC-deliver|Abn pelv org NEC-deliver
C0157060|T190|AB|654.92|ICD9CM|Abn pelv NEC-deliv w p/p|Abn pelv NEC-deliv w p/p
C0157061|T190|AB|654.93|ICD9CM|Abn pelv org NEC-antepar|Abn pelv org NEC-antepar
C0157062|T190|AB|654.94|ICD9CM|Abn pelv org NEC-postpar|Abn pelv org NEC-postpar
C0157063|T046|HT|655|ICD9CM|Known or suspected fetal abnormality affecting management of mother|Known or suspected fetal abnormality affecting management of mother
C0157064|T033|HT|655.0|ICD9CM|Central nervous system malformation in fetus affecting management of mother|Central nervous system malformation in fetus affecting management of mother
C0157065|T033|PT|655.00|ICD9CM|Central nervous system malformation in fetus, unspecified as to episode of care or not applicable|Central nervous system malformation in fetus, unspecified as to episode of care or not applicable
C0157065|T033|AB|655.00|ICD9CM|Fetal cns malform-unspec|Fetal cns malform-unspec
C0157066|T019|AB|655.01|ICD9CM|Fetal cns malform-deliv|Fetal cns malform-deliv
C0157066|T047|AB|655.01|ICD9CM|Fetal cns malform-deliv|Fetal cns malform-deliv
C0157067|T033|PT|655.03|ICD9CM|Central nervous system malformation in fetus, antepartum condition or complication|Central nervous system malformation in fetus, antepartum condition or complication
C0157067|T033|AB|655.03|ICD9CM|Fetal cns malfor-antepar|Fetal cns malfor-antepar
C0157068|T047|HT|655.1|ICD9CM|Chromosomal abnormality in fetus affecting management of mother|Chromosomal abnormality in fetus affecting management of mother
C0157069|T033|AB|655.10|ICD9CM|Fetal chromos abn-unspec|Fetal chromos abn-unspec
C0157070|T033|AB|655.11|ICD9CM|Fetal chromoso abn-deliv|Fetal chromoso abn-deliv
C0157071|T033|AB|655.13|ICD9CM|Fet chromo abn-antepart|Fet chromo abn-antepart
C0157072|T047|HT|655.2|ICD9CM|Hereditary disease in family possibly affecting fetus, affecting management of mother|Hereditary disease in family possibly affecting fetus, affecting management of mother
C0157073|T047|AB|655.20|ICD9CM|Famil heredit dis-unspec|Famil heredit dis-unspec
C0157074|T047|AB|655.21|ICD9CM|Famil heredit dis-deliv|Famil heredit dis-deliv
C0157075|T047|AB|655.23|ICD9CM|Famil hered dis-antepart|Famil hered dis-antepart
C0157076|T047|HT|655.3|ICD9CM|Suspected damage to fetus from viral disease in the mother, affecting management of mother|Suspected damage to fetus from viral disease in the mother, affecting management of mother
C0157077|T047|AB|655.30|ICD9CM|Fet damg d/t virus-unsp|Fet damg d/t virus-unsp
C0157078|T047|AB|655.31|ICD9CM|Fet damg d/t virus-deliv|Fet damg d/t virus-deliv
C0157079|T047|AB|655.33|ICD9CM|Fet damg d/t virus-antep|Fet damg d/t virus-antep
C0157080|T047|HT|655.4|ICD9CM|Suspected damage to fetus from other disease in the mother, affecting management of mother|Suspected damage to fetus from other disease in the mother, affecting management of mother
C0157081|T047|AB|655.40|ICD9CM|Fet damg d/t dis-unspec|Fet damg d/t dis-unspec
C0157082|T047|AB|655.41|ICD9CM|Fet damg d/t dis-deliver|Fet damg d/t dis-deliver
C0157083|T047|AB|655.43|ICD9CM|Fet damg d/t dis-antepar|Fet damg d/t dis-antepar
C0157084|T037|HT|655.5|ICD9CM|Suspected damage to fetus from drugs, affecting management of mother|Suspected damage to fetus from drugs, affecting management of mother
C0157085|T047|AB|655.50|ICD9CM|Fetal damg d/t drug-unsp|Fetal damg d/t drug-unsp
C0157086|T047|AB|655.51|ICD9CM|Fet damag d/t drug-deliv|Fet damag d/t drug-deliv
C0157087|T047|AB|655.53|ICD9CM|Fet damg d/t drug-antepa|Fet damg d/t drug-antepa
C0157088|T037|HT|655.6|ICD9CM|Suspected damage to fetus from radiation, affecting management of mother|Suspected damage to fetus from radiation, affecting management of mother
C0157089|T037|AB|655.60|ICD9CM|Radiat fetal damag-unsp|Radiat fetal damag-unsp
C0157090|T047|AB|655.61|ICD9CM|Radiat fetal damag-deliv|Radiat fetal damag-deliv
C0157090|T047|PT|655.61|ICD9CM|Suspected damage to fetus from radiation, affecting management of mother, delivered,|Suspected damage to fetus from radiation, affecting management of mother, delivered,
C0157091|T037|AB|655.63|ICD9CM|Radiat fet damag-antepar|Radiat fet damag-antepar
C0490008|T046|HT|655.7|ICD9CM|Decreased fetal movements, affecting management of mother|Decreased fetal movements, affecting management of mother
C0695214|T046|AB|655.70|ICD9CM|Decrease fetl movmt unsp|Decrease fetl movmt unsp
C0695214|T046|PT|655.70|ICD9CM|Decreased fetal movements, affecting management of mother, unspecified as to episode of care|Decreased fetal movements, affecting management of mother, unspecified as to episode of care
C0695215|T046|AB|655.71|ICD9CM|Decrease fetal movmt del|Decrease fetal movmt del
C0695216|T046|AB|655.73|ICD9CM|Dec fetal movmt antepart|Dec fetal movmt antepart
C0695216|T046|PT|655.73|ICD9CM|Decreased fetal movements, affecting management of mother, antepartum condition or complication|Decreased fetal movements, affecting management of mother, antepartum condition or complication
C0869483|T047|HT|655.8|ICD9CM|Other known or suspected fetal abnormality, not elsewhere classified, affecting management of mother|Other known or suspected fetal abnormality, not elsewhere classified, affecting management of mother
C0157093|T047|AB|655.80|ICD9CM|Fetal abnorm NEC-unspec|Fetal abnorm NEC-unspec
C0157094|T047|AB|655.81|ICD9CM|Fetal abnorm NEC-deliver|Fetal abnorm NEC-deliver
C0157095|T047|AB|655.83|ICD9CM|Fetal abnorm NEC-antepar|Fetal abnorm NEC-antepar
C0157063|T046|HT|655.9|ICD9CM|Unspecified, known or suspected fetal abnormality affecting management of mother|Unspecified, known or suspected fetal abnormality affecting management of mother
C0157097|T047|AB|655.90|ICD9CM|Fetal abnorm NOS-unspec|Fetal abnorm NOS-unspec
C0157098|T047|AB|655.91|ICD9CM|Fetal abnorm NOS-deliver|Fetal abnorm NOS-deliver
C0157099|T047|AB|655.93|ICD9CM|Fetal abnorm NOS-antepar|Fetal abnorm NOS-antepar
C2349589|T047|HT|656|ICD9CM|Other known or suspected fetal and placental problems affecting management of mother|Other known or suspected fetal and placental problems affecting management of mother
C0157101|T046|HT|656.0|ICD9CM|Fetal-maternal hemorrhage affecting management of mother|Fetal-maternal hemorrhage affecting management of mother
C0015959|T046|AB|656.00|ICD9CM|Fetal-maternal hem-unsp|Fetal-maternal hem-unsp
C0015959|T046|PT|656.00|ICD9CM|Fetal-maternal hemorrhage, unspecified as to episode of care or not applicable|Fetal-maternal hemorrhage, unspecified as to episode of care or not applicable
C0157103|T047|AB|656.01|ICD9CM|Fetal-maternal hem-deliv|Fetal-maternal hem-deliv
C0157103|T047|PT|656.01|ICD9CM|Fetal-maternal hemorrhage, delivered, with or without mention of antepartum condition|Fetal-maternal hemorrhage, delivered, with or without mention of antepartum condition
C0157104|T047|AB|656.03|ICD9CM|Fetal-matern hem-antepar|Fetal-matern hem-antepar
C0157104|T047|PT|656.03|ICD9CM|Fetal-maternal hemorrhage, antepartum condition or complication|Fetal-maternal hemorrhage, antepartum condition or complication
C0035428|T033|HT|656.1|ICD9CM|Rhesus isoimmunization affecting management of mother|Rhesus isoimmunization affecting management of mother
C0157105|T047|AB|656.10|ICD9CM|Rh isoimmunization-unsp|Rh isoimmunization-unsp
C0157105|T047|PT|656.10|ICD9CM|Rhesus isoimmunization, unspecified as to episode of care or not applicable|Rhesus isoimmunization, unspecified as to episode of care or not applicable
C0157106|T047|AB|656.11|ICD9CM|Rh isoimmunizat-deliver|Rh isoimmunizat-deliver
C0157106|T047|PT|656.11|ICD9CM|Rhesus isoimmunization, delivered, with or without mention of antepartum condition|Rhesus isoimmunization, delivered, with or without mention of antepartum condition
C0157107|T047|AB|656.13|ICD9CM|Rh isoimmunizat-antepart|Rh isoimmunizat-antepart
C0157107|T047|PT|656.13|ICD9CM|Rhesus isoimmunization, antepartum condition or complication|Rhesus isoimmunization, antepartum condition or complication
C0157109|T047|AB|656.20|ICD9CM|Abo isoimmunization-unsp|Abo isoimmunization-unsp
C0157110|T047|AB|656.21|ICD9CM|Abo isoimmunizat-deliver|Abo isoimmunizat-deliver
C0157111|T047|AB|656.23|ICD9CM|Abo isoimmunizat-antepar|Abo isoimmunizat-antepar
C0015931|T047|HT|656.3|ICD9CM|Fetal distress affecting management of mother|Fetal distress affecting management of mother
C0157112|T033|AB|656.30|ICD9CM|Fetal distress-unspec|Fetal distress-unspec
C0157112|T033|PT|656.30|ICD9CM|Fetal distress, affecting management of mother, unspecified as to episode of care or not applicable|Fetal distress, affecting management of mother, unspecified as to episode of care or not applicable
C0157113|T047|AB|656.31|ICD9CM|Fetal distress-delivered|Fetal distress-delivered
C0157114|T047|AB|656.33|ICD9CM|Fetal distress-antepart|Fetal distress-antepart
C0157114|T047|PT|656.33|ICD9CM|Fetal distress, affecting management of mother, antepartum condition or complication|Fetal distress, affecting management of mother, antepartum condition or complication
C0269792|T033|HT|656.4|ICD9CM|Intrauterine death affecting management of mother|Intrauterine death affecting management of mother
C0157116|T047|AB|656.40|ICD9CM|Intrauterine death-unsp|Intrauterine death-unsp
C0157117|T047|AB|656.41|ICD9CM|Intrauter death-deliver|Intrauter death-deliver
C0157118|T047|AB|656.43|ICD9CM|Intrauter death-antepart|Intrauter death-antepart
C0157118|T047|PT|656.43|ICD9CM|Intrauterine death, affecting management of mother, antepartum condition or complication|Intrauterine death, affecting management of mother, antepartum condition or complication
C0157119|T033|HT|656.5|ICD9CM|Poor fetal growth affecting management of mother|Poor fetal growth affecting management of mother
C0157120|T033|AB|656.50|ICD9CM|Poor fetal growth-unspec|Poor fetal growth-unspec
C0157121|T033|AB|656.51|ICD9CM|Poor fetal growth-deliv|Poor fetal growth-deliv
C0157122|T047|PT|656.53|ICD9CM|Poor fetal growth, affecting management of mother, antepartum condition or complication|Poor fetal growth, affecting management of mother, antepartum condition or complication
C0157122|T047|AB|656.53|ICD9CM|Poor fetal grth-antepart|Poor fetal grth-antepart
C0157123|T046|HT|656.6|ICD9CM|Excessive fetal growth affecting management of mother|Excessive fetal growth affecting management of mother
C0157124|T046|AB|656.60|ICD9CM|Excess fetal grth-unspec|Excess fetal grth-unspec
C0157125|T046|AB|656.61|ICD9CM|Excess fetal grth-deliv|Excess fetal grth-deliv
C0157126|T046|AB|656.63|ICD9CM|Excess fet grth-antepart|Excess fet grth-antepart
C0157126|T046|PT|656.63|ICD9CM|Excessive fetal growth, affecting management of mother, antepartum condition or complication|Excessive fetal growth, affecting management of mother, antepartum condition or complication
C0477835|T046|HT|656.7|ICD9CM|Other placental conditions affecting management of mother|Other placental conditions affecting management of mother
C0157127|T047|AB|656.70|ICD9CM|Oth placent cond-unspec|Oth placent cond-unspec
C0157128|T047|AB|656.71|ICD9CM|Oth placent cond-deliver|Oth placent cond-deliver
C0157129|T047|AB|656.73|ICD9CM|Oth placent cond-antepar|Oth placent cond-antepar
C0157129|T047|PT|656.73|ICD9CM|Other placental conditions, affecting management of mother, antepartum condition or complication|Other placental conditions, affecting management of mother, antepartum condition or complication
C0157130|T047|HT|656.8|ICD9CM|Other specified fetal and placental problems affecting management of mother|Other specified fetal and placental problems affecting management of mother
C0157131|T047|AB|656.80|ICD9CM|Fet/plac prob NEC-unspec|Fet/plac prob NEC-unspec
C0157132|T047|AB|656.81|ICD9CM|Fet/plac prob NEC-deliv|Fet/plac prob NEC-deliv
C0157133|T047|AB|656.83|ICD9CM|Fet/plac prob NEC-antepa|Fet/plac prob NEC-antepa
C0157134|T047|HT|656.9|ICD9CM|Unspecified fetal and placental problem affecting management of mother|Unspecified fetal and placental problem affecting management of mother
C0157135|T047|AB|656.90|ICD9CM|Fet/plac prob NOS-unspec|Fet/plac prob NOS-unspec
C0157136|T047|AB|656.91|ICD9CM|Fet/plac prob NOS-deliv|Fet/plac prob NOS-deliv
C0157137|T047|AB|656.93|ICD9CM|Fet/plac prob NOS-antepa|Fet/plac prob NOS-antepa
C0020224|T046|HT|657|ICD9CM|Polyhydramnios|Polyhydramnios
C0020224|T046|HT|657.0|ICD9CM|Polyhydramnios|Polyhydramnios
C1812620|T047|AB|657.00|ICD9CM|Polyhydramnios-unspec|Polyhydramnios-unspec
C1812620|T047|PT|657.00|ICD9CM|Polyhydramnios, unspecified as to episode of care or not applicable|Polyhydramnios, unspecified as to episode of care or not applicable
C0375434|T047|AB|657.01|ICD9CM|Polyhydramnios-delivered|Polyhydramnios-delivered
C0375434|T047|PT|657.01|ICD9CM|Polyhydramnios, delivered, with or without mention of antepartum condition|Polyhydramnios, delivered, with or without mention of antepartum condition
C0375436|T046|AB|657.03|ICD9CM|Polyhydramnios-antepart|Polyhydramnios-antepart
C0375436|T046|PT|657.03|ICD9CM|Polyhydramnios, antepartum condition or complication|Polyhydramnios, antepartum condition or complication
C0029715|T047|HT|658|ICD9CM|Other problems associated with amniotic cavity and membranes|Other problems associated with amniotic cavity and membranes
C0079924|T046|HT|658.0|ICD9CM|Oligohydramnios|Oligohydramnios
C0157141|T047|AB|658.00|ICD9CM|Oligohydramnios-unspec|Oligohydramnios-unspec
C0157141|T047|PT|658.00|ICD9CM|Oligohydramnios, unspecified as to episode of care or not applicable|Oligohydramnios, unspecified as to episode of care or not applicable
C0157142|T046|AB|658.01|ICD9CM|Oligohydramnios-deliver|Oligohydramnios-deliver
C0157142|T046|PT|658.01|ICD9CM|Oligohydramnios, delivered, with or without mention of antepartum condition|Oligohydramnios, delivered, with or without mention of antepartum condition
C0157143|T047|AB|658.03|ICD9CM|Oligohydramnios-antepar|Oligohydramnios-antepar
C0157143|T047|PT|658.03|ICD9CM|Oligohydramnios, antepartum condition or complication|Oligohydramnios, antepartum condition or complication
C0015944|T046|HT|658.1|ICD9CM|Premature rupture of membranes|Premature rupture of membranes
C0157145|T047|AB|658.10|ICD9CM|Prem rupt membran-unspec|Prem rupt membran-unspec
C0157145|T047|PT|658.10|ICD9CM|Premature rupture of membranes, unspecified as to episode of care or not applicable|Premature rupture of membranes, unspecified as to episode of care or not applicable
C0157146|T046|AB|658.11|ICD9CM|Prem rupt membran-deliv|Prem rupt membran-deliv
C0157146|T046|PT|658.11|ICD9CM|Premature rupture of membranes, delivered, with or without mention of antepartum condition|Premature rupture of membranes, delivered, with or without mention of antepartum condition
C0157147|T046|AB|658.13|ICD9CM|Prem rupt memb-antepart|Prem rupt memb-antepart
C0157147|T046|PT|658.13|ICD9CM|Premature rupture of membranes, antepartum condition or complication|Premature rupture of membranes, antepartum condition or complication
C0495246|T046|HT|658.2|ICD9CM|Delayed delivery after spontaneous or unspecified rupture of membranes|Delayed delivery after spontaneous or unspecified rupture of membranes
C0157149|T047|AB|658.20|ICD9CM|Prolong rupt memb-unspec|Prolong rupt memb-unspec
C0157150|T047|AB|658.21|ICD9CM|Prolong rupt memb-deliv|Prolong rupt memb-deliv
C0157151|T047|AB|658.23|ICD9CM|Prolong rup memb-antepar|Prolong rup memb-antepar
C0157152|T046|HT|658.3|ICD9CM|Delayed delivery after artificial rupture of membranes|Delayed delivery after artificial rupture of membranes
C0157153|T047|AB|658.30|ICD9CM|Artific rupt membr-unsp|Artific rupt membr-unsp
C0157154|T047|AB|658.31|ICD9CM|Artific rupt membr-deliv|Artific rupt membr-deliv
C0157155|T047|AB|658.33|ICD9CM|Artif rupt memb-antepart|Artif rupt memb-antepart
C0157155|T047|PT|658.33|ICD9CM|Delayed delivery after artificial rupture of membranes, antepartum condition or complication|Delayed delivery after artificial rupture of membranes, antepartum condition or complication
C0002631|T047|HT|658.4|ICD9CM|Infection of amniotic cavity|Infection of amniotic cavity
C0002631|T047|AB|658.40|ICD9CM|Amniotic infection-unsp|Amniotic infection-unsp
C0002631|T047|PT|658.40|ICD9CM|Infection of amniotic cavity, unspecified as to episode of care or not applicable|Infection of amniotic cavity, unspecified as to episode of care or not applicable
C0157157|T046|AB|658.41|ICD9CM|Amniotic infection-deliv|Amniotic infection-deliv
C0157157|T046|PT|658.41|ICD9CM|Infection of amniotic cavity, delivered, with or without mention of antepartum condition|Infection of amniotic cavity, delivered, with or without mention of antepartum condition
C0157158|T047|AB|658.43|ICD9CM|Amniotic infect-antepart|Amniotic infect-antepart
C0157158|T047|PT|658.43|ICD9CM|Infection of amniotic cavity, antepartum condition or complication|Infection of amniotic cavity, antepartum condition or complication
C0029715|T047|HT|658.8|ICD9CM|Other problems associated with amniotic cavity and membranes|Other problems associated with amniotic cavity and membranes
C0157159|T047|AB|658.80|ICD9CM|Amniotic prob NEC-unspec|Amniotic prob NEC-unspec
C0157160|T047|AB|658.81|ICD9CM|Amniotic prob NEC-deliv|Amniotic prob NEC-deliv
C0157161|T047|AB|658.83|ICD9CM|Amnion prob NEC-antepart|Amnion prob NEC-antepart
C0157161|T047|PT|658.83|ICD9CM|Other problems associated with amniotic cavity and membranes, antepartum|Other problems associated with amniotic cavity and membranes, antepartum
C0405034|T047|HT|658.9|ICD9CM|Unspecified problem associated with amniotic cavity and membranes|Unspecified problem associated with amniotic cavity and membranes
C0405037|T033|AB|658.90|ICD9CM|Amniotic prob NOS-unspec|Amniotic prob NOS-unspec
C2114658|T047|AB|658.91|ICD9CM|Amniotic prob NOS-deliv|Amniotic prob NOS-deliv
C0157165|T047|AB|658.93|ICD9CM|Amnion prob NOS-antepart|Amnion prob NOS-antepart
C0302388|T047|HT|659|ICD9CM|Other indications for care or intervention related to labor and delivery, not elsewhere classified|Other indications for care or intervention related to labor and delivery, not elsewhere classified
C0269807|T046|HT|659.0|ICD9CM|Failed mechanical induction of labor|Failed mechanical induction of labor
C0157168|T047|AB|659.00|ICD9CM|Fail mechan induct-unsp|Fail mechan induct-unsp
C0157168|T047|PT|659.00|ICD9CM|Failed mechanical induction of labor, unspecified as to episode of care or not applicable|Failed mechanical induction of labor, unspecified as to episode of care or not applicable
C0157169|T033|AB|659.01|ICD9CM|Fail mech induct-deliver|Fail mech induct-deliver
C0157169|T033|PT|659.01|ICD9CM|Failed mechanical induction of labor, delivered, with or without mention of antepartum condition|Failed mechanical induction of labor, delivered, with or without mention of antepartum condition
C0157170|T047|AB|659.03|ICD9CM|Fail mech induct-antepar|Fail mech induct-antepar
C0157170|T047|PT|659.03|ICD9CM|Failed mechanical induction of labor, antepartum condition or complication|Failed mechanical induction of labor, antepartum condition or complication
C0405189|T046|HT|659.1|ICD9CM|Failed medical or unspecified induction of labor|Failed medical or unspecified induction of labor
C0157172|T047|AB|659.10|ICD9CM|Fail induction NOS-unsp|Fail induction NOS-unsp
C0157173|T047|AB|659.11|ICD9CM|Fail induction NOS-deliv|Fail induction NOS-deliv
C0157174|T047|AB|659.13|ICD9CM|Fail induct NOS-antepart|Fail induct NOS-antepart
C0157174|T047|PT|659.13|ICD9CM|Failed medical or unspecified induction of labor, antepartum condition or complication|Failed medical or unspecified induction of labor, antepartum condition or complication
C0341973|T046|HT|659.2|ICD9CM|Maternal pyrexia during labor, unspecified|Maternal pyrexia during labor, unspecified
C0157176|T047|PT|659.20|ICD9CM|Maternal pyrexia during labor, unspecified, unspecified as to episode of care or not applicable|Maternal pyrexia during labor, unspecified, unspecified as to episode of care or not applicable
C0157176|T047|AB|659.20|ICD9CM|Pyrexia in labor-unspec|Pyrexia in labor-unspec
C0157177|T047|AB|659.21|ICD9CM|Pyrexia in labor-deliver|Pyrexia in labor-deliver
C0157178|T047|PT|659.23|ICD9CM|Maternal pyrexia during labor, unspecified, antepartum condition or complication|Maternal pyrexia during labor, unspecified, antepartum condition or complication
C0157178|T047|AB|659.23|ICD9CM|Pyrexia in labor-antepar|Pyrexia in labor-antepar
C0157179|T046|HT|659.3|ICD9CM|Generalized infection during labor|Generalized infection during labor
C0157180|T047|PT|659.30|ICD9CM|Generalized infection during labor, unspecified as to episode of care or not applicable|Generalized infection during labor, unspecified as to episode of care or not applicable
C0157180|T047|AB|659.30|ICD9CM|Septicemia in labor-unsp|Septicemia in labor-unsp
C0157181|T047|PT|659.31|ICD9CM|Generalized infection during labor, delivered, with or without mention of antepartum condition|Generalized infection during labor, delivered, with or without mention of antepartum condition
C0157181|T047|AB|659.31|ICD9CM|Septicem in labor-deliv|Septicem in labor-deliv
C0157182|T047|PT|659.33|ICD9CM|Generalized infection during labor, antepartum condition or complication|Generalized infection during labor, antepartum condition or complication
C0157182|T047|AB|659.33|ICD9CM|Septicem in labor-antepa|Septicem in labor-antepa
C0157183|T033|HT|659.4|ICD9CM|Grand multiparity, with current pregnancy|Grand multiparity, with current pregnancy
C0157184|T033|AB|659.40|ICD9CM|Grand multiparity-unspec|Grand multiparity-unspec
C0157184|T033|PT|659.40|ICD9CM|Grand multiparity, unspecified as to episode of care or not applicable|Grand multiparity, unspecified as to episode of care or not applicable
C0157185|T033|AB|659.41|ICD9CM|Grand multiparity-deliv|Grand multiparity-deliv
C0157185|T033|PT|659.41|ICD9CM|Grand multiparity, delivered, with or without mention of antepartum condition|Grand multiparity, delivered, with or without mention of antepartum condition
C0157186|T033|AB|659.43|ICD9CM|Grand multiparity-antepa|Grand multiparity-antepa
C0157186|T033|PT|659.43|ICD9CM|Grand multiparity, antepartum condition or complication|Grand multiparity, antepartum condition or complication
C0157187|T033|HT|659.5|ICD9CM|Elderly primigravida|Elderly primigravida
C0157189|T033|AB|659.51|ICD9CM|Elderly primigravida-del|Elderly primigravida-del
C0157189|T033|PT|659.51|ICD9CM|Elderly primigravida, delivered, with or without mention of antepartum condition|Elderly primigravida, delivered, with or without mention of antepartum condition
C0695245|T046|HT|659.7|ICD9CM|Abnormality in fetal heart rate or rhythm|Abnormality in fetal heart rate or rhythm
C0695246|T046|AB|659.70|ICD9CM|Abn ftl hrt rate/rhy-uns|Abn ftl hrt rate/rhy-uns
C0695246|T046|PT|659.70|ICD9CM|Abnormality in fetal heart rate or rhythm, unspecified as to episode of care or not applicable|Abnormality in fetal heart rate or rhythm, unspecified as to episode of care or not applicable
C0695247|T046|AB|659.71|ICD9CM|Abn ftl hrt rate/rhy-del|Abn ftl hrt rate/rhy-del
C0695248|T046|AB|659.73|ICD9CM|Abn ftl hrt rate/rhy-ant|Abn ftl hrt rate/rhy-ant
C0695248|T046|PT|659.73|ICD9CM|Abnormality in fetal heart rate or rhythm, antepartum condition or complication|Abnormality in fetal heart rate or rhythm, antepartum condition or complication
C0157191|T033|HT|659.8|ICD9CM|Other specified indications for care or intervention related to labor and delivery|Other specified indications for care or intervention related to labor and delivery
C0157192|T033|AB|659.80|ICD9CM|Complic labor NEC-unsp|Complic labor NEC-unsp
C0157193|T047|AB|659.81|ICD9CM|Complic labor NEC-deliv|Complic labor NEC-deliv
C0157194|T047|AB|659.83|ICD9CM|Compl labor NEC-antepart|Compl labor NEC-antepart
C0157195|T033|HT|659.9|ICD9CM|Unspecified indication for care or intervention related to labor and delivery|Unspecified indication for care or intervention related to labor and delivery
C0157196|T033|AB|659.90|ICD9CM|Complic labor NOS-unsp|Complic labor NOS-unsp
C0157197|T047|AB|659.91|ICD9CM|Complic labor NOS-deliv|Complic labor NOS-deliv
C0157198|T047|AB|659.93|ICD9CM|Compl labor NOS-antepart|Compl labor NOS-antepart
C0152156|T046|HT|660|ICD9CM|Obstructed labor|Obstructed labor
C0178297|T047|HT|660-669.99|ICD9CM|COMPLICATIONS OCCURRING MAINLY IN THE COURSE OF LABOR AND DELIVERY|COMPLICATIONS OCCURRING MAINLY IN THE COURSE OF LABOR AND DELIVERY
C0157199|T046|HT|660.0|ICD9CM|Obstruction caused by malposition of fetus at onset of labor|Obstruction caused by malposition of fetus at onset of labor
C0157200|T046|AB|660.00|ICD9CM|Obstruct/fet malpos-unsp|Obstruct/fet malpos-unsp
C0157201|T046|AB|660.01|ICD9CM|Obstruc/fet malpos-deliv|Obstruc/fet malpos-deliv
C0157202|T046|AB|660.03|ICD9CM|Obstruc/fet malpos-antep|Obstruc/fet malpos-antep
C0157202|T046|PT|660.03|ICD9CM|Obstruction caused by malposition of fetus at onset of labor, antepartum condition or complication|Obstruction caused by malposition of fetus at onset of labor, antepartum condition or complication
C0157203|T033|HT|660.1|ICD9CM|Obstruction by bony pelvis during labor|Obstruction by bony pelvis during labor
C0157204|T047|AB|660.10|ICD9CM|Bony pelv obstruc-unspec|Bony pelv obstruc-unspec
C0157204|T047|PT|660.10|ICD9CM|Obstruction by bony pelvis during labor, unspecified as to episode of care or not applicable|Obstruction by bony pelvis during labor, unspecified as to episode of care or not applicable
C0157205|T047|AB|660.11|ICD9CM|Bony pelv obstruct-deliv|Bony pelv obstruct-deliv
C0157205|T047|PT|660.11|ICD9CM|Obstruction by bony pelvis during labor, delivered, with or without mention of antepartum condition|Obstruction by bony pelvis during labor, delivered, with or without mention of antepartum condition
C0157206|T047|AB|660.13|ICD9CM|Bony pelv obstruc-antepa|Bony pelv obstruc-antepa
C0157206|T047|PT|660.13|ICD9CM|Obstruction by bony pelvis during labor, antepartum condition or complication|Obstruction by bony pelvis during labor, antepartum condition or complication
C0157207|T033|HT|660.2|ICD9CM|Obstruction by abnormal pelvic soft tissues during labor|Obstruction by abnormal pelvic soft tissues during labor
C0157208|T046|AB|660.20|ICD9CM|Abn pelv tiss obstr-unsp|Abn pelv tiss obstr-unsp
C0157209|T047|AB|660.21|ICD9CM|Abn pelv tis obstr-deliv|Abn pelv tis obstr-deliv
C0157210|T047|AB|660.23|ICD9CM|Abn pelv tis obstr-antep|Abn pelv tis obstr-antep
C0157210|T047|PT|660.23|ICD9CM|Obstruction by abnormal pelvic soft tissues during labor, antepartum condition or complication|Obstruction by abnormal pelvic soft tissues during labor, antepartum condition or complication
C0157211|T047|HT|660.3|ICD9CM|Deep transverse arrest and persistent occipitoposterior position during labor and delivery|Deep transverse arrest and persistent occipitoposterior position during labor and delivery
C0157212|T033|AB|660.30|ICD9CM|Persist occipitpost-unsp|Persist occipitpost-unsp
C0157213|T047|AB|660.31|ICD9CM|Persist occiptpost-deliv|Persist occiptpost-deliv
C0157214|T047|AB|660.33|ICD9CM|Persist occiptpost-antep|Persist occiptpost-antep
C0269825|T046|HT|660.4|ICD9CM|Shoulder (girdle) dystocia during labor and delivery|Shoulder (girdle) dystocia during labor and delivery
C0157216|T033|PT|660.40|ICD9CM|Shoulder (girdle) dystocia, unspecified as to episode of care or not applicable|Shoulder (girdle) dystocia, unspecified as to episode of care or not applicable
C0157216|T033|AB|660.40|ICD9CM|Shoulder dystocia-unspec|Shoulder dystocia-unspec
C0748659|T047|PT|660.41|ICD9CM|Shoulder (girdle) dystocia, delivered, with or without mention of antepartum condition|Shoulder (girdle) dystocia, delivered, with or without mention of antepartum condition
C0748659|T047|AB|660.41|ICD9CM|Shoulder dystocia-deliv|Shoulder dystocia-deliv
C0157218|T033|PT|660.43|ICD9CM|Shoulder (girdle) dystocia, antepartum condition or complication|Shoulder (girdle) dystocia, antepartum condition or complication
C0157218|T033|AB|660.43|ICD9CM|Shoulder dystocia-antepa|Shoulder dystocia-antepa
C0405185|T033|HT|660.5|ICD9CM|Locked twins|Locked twins
C0157220|T047|AB|660.50|ICD9CM|Locked twins-unspecified|Locked twins-unspecified
C0157220|T047|PT|660.50|ICD9CM|Locked twins, unspecified as to episode of care or not applicable|Locked twins, unspecified as to episode of care or not applicable
C0157221|T047|AB|660.51|ICD9CM|Locked twins-delivered|Locked twins-delivered
C0157221|T047|PT|660.51|ICD9CM|Locked twins, delivered, with or without mention of antepartum condition|Locked twins, delivered, with or without mention of antepartum condition
C0157222|T047|AB|660.53|ICD9CM|Locked twins-antepartum|Locked twins-antepartum
C0157222|T047|PT|660.53|ICD9CM|Locked twins, antepartum condition or complication|Locked twins, antepartum condition or complication
C0157223|T046|HT|660.6|ICD9CM|Failed trial of labor, unspecified|Failed trial of labor, unspecified
C0157224|T033|AB|660.60|ICD9CM|Fail trial lab NOS-unsp|Fail trial lab NOS-unsp
C0157224|T033|PT|660.60|ICD9CM|Unspecified failed trial of labor, unspecified as to episode of care or not applicable|Unspecified failed trial of labor, unspecified as to episode of care or not applicable
C0157225|T047|AB|660.61|ICD9CM|Fail trial lab NOS-deliv|Fail trial lab NOS-deliv
C0157225|T047|PT|660.61|ICD9CM|Unspecified failed trial of labor, delivered, with or without mention of antepartum condition|Unspecified failed trial of labor, delivered, with or without mention of antepartum condition
C0157226|T047|AB|660.63|ICD9CM|Fail trial lab NOS-antep|Fail trial lab NOS-antep
C0157226|T047|PT|660.63|ICD9CM|Unspecified failed trial of labor, antepartum condition or complication|Unspecified failed trial of labor, antepartum condition or complication
C0495263|T046|HT|660.7|ICD9CM|Failed forceps or vacuum extractor, unspecified|Failed forceps or vacuum extractor, unspecified
C0157228|T047|AB|660.70|ICD9CM|Failed forcep NOS-unspec|Failed forcep NOS-unspec
C0157228|T047|PT|660.70|ICD9CM|Failed forceps or vacuum extractor, unspecified, unspecified as to episode of care or not applicable|Failed forceps or vacuum extractor, unspecified, unspecified as to episode of care or not applicable
C0157229|T047|AB|660.71|ICD9CM|Failed forceps NOS-deliv|Failed forceps NOS-deliv
C0157230|T047|AB|660.73|ICD9CM|Fail forceps NOS-antepar|Fail forceps NOS-antepar
C0157230|T047|PT|660.73|ICD9CM|Failed forceps or vacuum extractor, unspecified, antepartum condition or complication|Failed forceps or vacuum extractor, unspecified, antepartum condition or complication
C0157231|T033|HT|660.8|ICD9CM|Other causes of obstructed labor|Other causes of obstructed labor
C0157232|T047|AB|660.80|ICD9CM|Obstruc labor NEC-unspec|Obstruc labor NEC-unspec
C0157232|T047|PT|660.80|ICD9CM|Other causes of obstructed labor, unspecified as to episode of care or not applicable|Other causes of obstructed labor, unspecified as to episode of care or not applicable
C0157233|T047|AB|660.81|ICD9CM|Obstruct labor NEC-deliv|Obstruct labor NEC-deliv
C0157233|T047|PT|660.81|ICD9CM|Other causes of obstructed labor, delivered, with or without mention of antepartum condition|Other causes of obstructed labor, delivered, with or without mention of antepartum condition
C0157234|T047|AB|660.83|ICD9CM|Obstruc labor NEC-antepa|Obstruc labor NEC-antepa
C0157234|T047|PT|660.83|ICD9CM|Other causes of obstructed labor, antepartum condition or complication|Other causes of obstructed labor, antepartum condition or complication
C0152156|T046|HT|660.9|ICD9CM|Unspecified obstructed labor|Unspecified obstructed labor
C0157235|T047|AB|660.90|ICD9CM|Obstruc labor NOS-unspec|Obstruc labor NOS-unspec
C0157235|T047|PT|660.90|ICD9CM|Unspecified obstructed labor, unspecified as to episode of care or not applicable|Unspecified obstructed labor, unspecified as to episode of care or not applicable
C0157236|T047|AB|660.91|ICD9CM|Obstruct labor NOS-deliv|Obstruct labor NOS-deliv
C0157236|T047|PT|660.91|ICD9CM|Unspecified obstructed labor, delivered, with or without mention of antepartum condition|Unspecified obstructed labor, delivered, with or without mention of antepartum condition
C0157237|T047|AB|660.93|ICD9CM|Obstruc labor NOS-antepa|Obstruc labor NOS-antepa
C0157237|T047|PT|660.93|ICD9CM|Unspecified obstructed labor, antepartum condition or complication|Unspecified obstructed labor, antepartum condition or complication
C0473462|T046|HT|661|ICD9CM|Abnormality of forces of labor|Abnormality of forces of labor
C0152159|T047|HT|661.0|ICD9CM|Primary uterine inertia|Primary uterine inertia
C0157239|T047|AB|661.00|ICD9CM|Prim uterine inert-unsp|Prim uterine inert-unsp
C0157239|T047|PT|661.00|ICD9CM|Primary uterine inertia, unspecified as to episode of care or not applicable|Primary uterine inertia, unspecified as to episode of care or not applicable
C0157240|T046|AB|661.01|ICD9CM|Prim uterine inert-deliv|Prim uterine inert-deliv
C0157240|T046|PT|661.01|ICD9CM|Primary uterine inertia, delivered, with or without mention of antepartum condition|Primary uterine inertia, delivered, with or without mention of antepartum condition
C0157241|T047|AB|661.03|ICD9CM|Prim uter inert-antepart|Prim uter inert-antepart
C0157241|T047|PT|661.03|ICD9CM|Primary uterine inertia, antepartum condition or complication|Primary uterine inertia, antepartum condition or complication
C0405169|T046|HT|661.1|ICD9CM|Secondary uterine inertia|Secondary uterine inertia
C0157242|T047|AB|661.10|ICD9CM|Sec uterine inert-unspec|Sec uterine inert-unspec
C0157242|T047|PT|661.10|ICD9CM|Secondary uterine inertia, unspecified as to episode of care or not applicable|Secondary uterine inertia, unspecified as to episode of care or not applicable
C0157243|T047|AB|661.11|ICD9CM|Sec uterine inert-deliv|Sec uterine inert-deliv
C0157243|T047|PT|661.11|ICD9CM|Secondary uterine inertia, delivered, with or without mention of antepartum condition|Secondary uterine inertia, delivered, with or without mention of antepartum condition
C0157244|T047|AB|661.13|ICD9CM|Sec uterine inert-antepa|Sec uterine inert-antepa
C0157244|T047|PT|661.13|ICD9CM|Secondary uterine inertia, antepartum condition or complication|Secondary uterine inertia, antepartum condition or complication
C0477838|T046|HT|661.2|ICD9CM|Other and unspecified uterine inertia|Other and unspecified uterine inertia
C0477838|T046|PT|661.20|ICD9CM|Other and unspecified uterine inertia, unspecified as to episode of care or not applicable|Other and unspecified uterine inertia, unspecified as to episode of care or not applicable
C0477838|T046|AB|661.20|ICD9CM|Uterine inertia NEC-unsp|Uterine inertia NEC-unsp
C0157246|T047|PT|661.21|ICD9CM|Other and unspecified uterine inertia, delivered, with or without mention of antepartum condition|Other and unspecified uterine inertia, delivered, with or without mention of antepartum condition
C0157246|T047|AB|661.21|ICD9CM|Uterine inert NEC-deliv|Uterine inert NEC-deliv
C0157247|T047|PT|661.23|ICD9CM|Other and unspecified uterine inertia, antepartum condition or complication|Other and unspecified uterine inertia, antepartum condition or complication
C0157247|T047|AB|661.23|ICD9CM|Uterine inert NEC-antepa|Uterine inert NEC-antepa
C0473472|T046|HT|661.3|ICD9CM|Precipitate labor|Precipitate labor
C0157248|T047|AB|661.30|ICD9CM|Precipitate labor-unspec|Precipitate labor-unspec
C0157248|T047|PT|661.30|ICD9CM|Precipitate labor, unspecified as to episode of care or not applicable|Precipitate labor, unspecified as to episode of care or not applicable
C0157249|T047|AB|661.31|ICD9CM|Precipitate labor-deliv|Precipitate labor-deliv
C0157249|T047|PT|661.31|ICD9CM|Precipitate labor, delivered, with or without mention of antepartum condition|Precipitate labor, delivered, with or without mention of antepartum condition
C0157250|T047|AB|661.33|ICD9CM|Precipitate labor-antepa|Precipitate labor-antepa
C0157250|T047|PT|661.33|ICD9CM|Precipitate labor, antepartum condition or complication|Precipitate labor, antepartum condition or complication
C0495255|T046|HT|661.4|ICD9CM|Hypertonic, incoordinate, or prolonged uterine contractions|Hypertonic, incoordinate, or prolonged uterine contractions
C0157252|T047|AB|661.40|ICD9CM|Uter dystocia NOS-unspec|Uter dystocia NOS-unspec
C0157253|T047|AB|661.41|ICD9CM|Uter dystocia NOS-deliv|Uter dystocia NOS-deliv
C0157254|T047|PT|661.43|ICD9CM|Hypertonic, incoordinate, or prolonged uterine contractions, antepartum condition or complication|Hypertonic, incoordinate, or prolonged uterine contractions, antepartum condition or complication
C0157254|T047|AB|661.43|ICD9CM|Uter dystocia NOS-antepa|Uter dystocia NOS-antepa
C0013418|T046|HT|661.9|ICD9CM|Unspecified abnormality of labor|Unspecified abnormality of labor
C0157256|T047|AB|661.90|ICD9CM|Abnormal labor NOS-unsp|Abnormal labor NOS-unsp
C0157256|T047|PT|661.90|ICD9CM|Unspecified abnormality of labor, unspecified as to episode of care or not applicable|Unspecified abnormality of labor, unspecified as to episode of care or not applicable
C0473461|T046|AB|661.91|ICD9CM|Abnormal labor NOS-deliv|Abnormal labor NOS-deliv
C0473461|T046|PT|661.91|ICD9CM|Unspecified abnormality of labor, delivered, with or without mention of antepartum condition|Unspecified abnormality of labor, delivered, with or without mention of antepartum condition
C0157258|T047|AB|661.93|ICD9CM|Abnorm labor NOS-antepar|Abnorm labor NOS-antepar
C0157258|T047|PT|661.93|ICD9CM|Unspecified abnormality of labor, antepartum condition or complication|Unspecified abnormality of labor, antepartum condition or complication
C0152154|T046|HT|662|ICD9CM|Long labor|Long labor
C0157259|T046|HT|662.0|ICD9CM|Prolonged first stage of labor|Prolonged first stage of labor
C0157260|T047|AB|662.00|ICD9CM|Prolonged 1st stage-unsp|Prolonged 1st stage-unsp
C0157260|T047|PT|662.00|ICD9CM|Prolonged first stage of labor, unspecified as to episode of care or not applicable|Prolonged first stage of labor, unspecified as to episode of care or not applicable
C0157261|T047|AB|662.01|ICD9CM|Prolong 1st stage-deliv|Prolong 1st stage-deliv
C0157261|T047|PT|662.01|ICD9CM|Prolonged first stage of labor, delivered, with or without mention of antepartum condition|Prolonged first stage of labor, delivered, with or without mention of antepartum condition
C0157262|T047|AB|662.03|ICD9CM|Prolong 1st stage-antepa|Prolong 1st stage-antepa
C0157262|T047|PT|662.03|ICD9CM|Prolonged first stage of labor, antepartum condition or complication|Prolonged first stage of labor, antepartum condition or complication
C0152154|T046|HT|662.1|ICD9CM|Prolonged labor, unspecified|Prolonged labor, unspecified
C0157263|T047|AB|662.10|ICD9CM|Prolonged labor NOS-unsp|Prolonged labor NOS-unsp
C0157263|T047|PT|662.10|ICD9CM|Unspecified prolonged labor, unspecified as to episode of care or not applicable|Unspecified prolonged labor, unspecified as to episode of care or not applicable
C0157264|T047|AB|662.11|ICD9CM|Prolong labor NOS-deliv|Prolong labor NOS-deliv
C0157264|T047|PT|662.11|ICD9CM|Unspecified prolonged labor, delivered, with or without mention of antepartum condition|Unspecified prolonged labor, delivered, with or without mention of antepartum condition
C0157265|T047|AB|662.13|ICD9CM|Prolong labor NOS-antepa|Prolong labor NOS-antepa
C0157265|T047|PT|662.13|ICD9CM|Unspecified prolonged labor, antepartum condition or complication|Unspecified prolonged labor, antepartum condition or complication
C0157266|T046|HT|662.2|ICD9CM|Prolonged second stage of labor|Prolonged second stage of labor
C0157267|T047|AB|662.20|ICD9CM|Prolonged 2nd stage-unsp|Prolonged 2nd stage-unsp
C0157267|T047|PT|662.20|ICD9CM|Prolonged second stage of labor, unspecified as to episode of care or not applicable|Prolonged second stage of labor, unspecified as to episode of care or not applicable
C0157268|T047|AB|662.21|ICD9CM|Prolong 2nd stage-deliv|Prolong 2nd stage-deliv
C0157268|T047|PT|662.21|ICD9CM|Prolonged second stage of labor, delivered, with or without mention of antepartum condition|Prolonged second stage of labor, delivered, with or without mention of antepartum condition
C0157269|T047|AB|662.23|ICD9CM|Prolong 2nd stage-antepa|Prolong 2nd stage-antepa
C0157269|T047|PT|662.23|ICD9CM|Prolonged second stage of labor, antepartum condition or complication|Prolonged second stage of labor, antepartum condition or complication
C0157270|T046|HT|662.3|ICD9CM|Delayed delivery of second twin, triplet, etc.|Delayed delivery of second twin, triplet, etc.
C0157271|T047|AB|662.30|ICD9CM|Delay del 2nd twin-unsp|Delay del 2nd twin-unsp
C0157271|T047|PT|662.30|ICD9CM|Delayed delivery of second twin, triplet, etc., unspecified as to episode of care or not applicable|Delayed delivery of second twin, triplet, etc., unspecified as to episode of care or not applicable
C0157272|T047|AB|662.31|ICD9CM|Delay del 2nd twin-deliv|Delay del 2nd twin-deliv
C0157270|T046|AB|662.33|ICD9CM|Delay del 2 twin-antepar|Delay del 2 twin-antepar
C0157270|T046|PT|662.33|ICD9CM|Delayed delivery of second twin, triplet, etc., antepartum condition or complication|Delayed delivery of second twin, triplet, etc., antepartum condition or complication
C0157307|T046|HT|663|ICD9CM|Umbilical cord complications during labor and delivery|Umbilical cord complications during labor and delivery
C0157275|T046|HT|663.0|ICD9CM|Prolapse of cord complicating labor and delivery|Prolapse of cord complicating labor and delivery
C0157275|T046|AB|663.00|ICD9CM|Cord prolapse-unspec|Cord prolapse-unspec
C0157277|T047|AB|663.01|ICD9CM|Cord prolapse-delivered|Cord prolapse-delivered
C0157278|T047|AB|663.03|ICD9CM|Cord prolapse-antepartum|Cord prolapse-antepartum
C0157278|T047|PT|663.03|ICD9CM|Prolapse of cord complicating labor and delivery, antepartum condition or complication|Prolapse of cord complicating labor and delivery, antepartum condition or complication
C0566742|T046|HT|663.1|ICD9CM|Cord around neck, with compression, complicating labor and delivery|Cord around neck, with compression, complicating labor and delivery
C0157280|T047|AB|663.10|ICD9CM|Cord around neck-unspec|Cord around neck-unspec
C0157281|T046|AB|663.11|ICD9CM|Cord around neck-deliver|Cord around neck-deliver
C0157282|T046|AB|663.13|ICD9CM|Cord around neck-antepar|Cord around neck-antepar
C0157283|T046|HT|663.2|ICD9CM|Other and unspecified cord entanglement, with compression, complicating labor and delivery|Other and unspecified cord entanglement, with compression, complicating labor and delivery
C0157284|T047|AB|663.20|ICD9CM|Cord compress NEC-unspec|Cord compress NEC-unspec
C0157285|T047|AB|663.21|ICD9CM|Cord compress NEC-deliv|Cord compress NEC-deliv
C0157286|T047|AB|663.23|ICD9CM|Cord compres NEC-antepar|Cord compres NEC-antepar
C0157288|T047|AB|663.30|ICD9CM|Cord entangle NEC-unspec|Cord entangle NEC-unspec
C0157289|T047|AB|663.31|ICD9CM|Cord entangle NEC-deliv|Cord entangle NEC-deliv
C0157290|T047|AB|663.33|ICD9CM|Cord entangl NEC-antepar|Cord entangl NEC-antepar
C0157291|T047|HT|663.4|ICD9CM|Short cord complicating labor and delivery|Short cord complicating labor and delivery
C0157292|T047|PT|663.40|ICD9CM|Short cord complicating labor and delivery, unspecified as to episode of care or not applicable|Short cord complicating labor and delivery, unspecified as to episode of care or not applicable
C0157292|T047|AB|663.40|ICD9CM|Short cord-unspecified|Short cord-unspecified
C0157293|T047|AB|663.41|ICD9CM|Short cord-delivered|Short cord-delivered
C0157294|T047|PT|663.43|ICD9CM|Short cord complicating labor and delivery, antepartum condition or complication|Short cord complicating labor and delivery, antepartum condition or complication
C0157294|T047|AB|663.43|ICD9CM|Short cord-antepartum|Short cord-antepartum
C0495270|T047|HT|663.5|ICD9CM|Vasa previa complicating labor and delivery|Vasa previa complicating labor and delivery
C0495270|T047|PT|663.50|ICD9CM|Vasa previa complicating labor and delivery, unspecified as to episode of care or not applicable|Vasa previa complicating labor and delivery, unspecified as to episode of care or not applicable
C0495270|T047|AB|663.50|ICD9CM|Vasa previa-unspecified|Vasa previa-unspecified
C0157297|T047|AB|663.51|ICD9CM|Vasa previa-delivered|Vasa previa-delivered
C0269852|T190|PT|663.53|ICD9CM|Vasa previa complicating labor and delivery, antepartum condition or complication|Vasa previa complicating labor and delivery, antepartum condition or complication
C0269852|T190|AB|663.53|ICD9CM|Vasa previa-antepartum|Vasa previa-antepartum
C0157299|T047|HT|663.6|ICD9CM|Vascular lesions of cord complicating labor and delivery|Vascular lesions of cord complicating labor and delivery
C0157300|T047|AB|663.60|ICD9CM|Vasc lesion cord-unspec|Vasc lesion cord-unspec
C0157301|T047|AB|663.61|ICD9CM|Vasc lesion cord-deliver|Vasc lesion cord-deliver
C0157302|T047|AB|663.63|ICD9CM|Vasc lesion cord-antepar|Vasc lesion cord-antepar
C0157302|T047|PT|663.63|ICD9CM|Vascular lesions of cord complicating labor and delivery, antepartum condition or complication|Vascular lesions of cord complicating labor and delivery, antepartum condition or complication
C0157303|T046|HT|663.8|ICD9CM|Other umbilical cord complications during labor and delivery|Other umbilical cord complications during labor and delivery
C0157304|T047|AB|663.80|ICD9CM|Cord complicat NEC-unsp|Cord complicat NEC-unsp
C0157305|T047|AB|663.81|ICD9CM|Cord complicat NEC-deliv|Cord complicat NEC-deliv
C0157306|T047|AB|663.83|ICD9CM|Cord compl NEC-antepart|Cord compl NEC-antepart
C0157307|T046|HT|663.9|ICD9CM|Unspecified umbilical cord complication during labor and delivery|Unspecified umbilical cord complication during labor and delivery
C0157308|T047|AB|663.90|ICD9CM|Cord complicat NOS-unsp|Cord complicat NOS-unsp
C0157309|T047|AB|663.91|ICD9CM|Cord complicat NOS-deliv|Cord complicat NOS-deliv
C0157310|T046|AB|663.93|ICD9CM|Cord compl NOS-antepart|Cord compl NOS-antepart
C0157311|T037|HT|664|ICD9CM|Trauma to perineum and vulva during delivery|Trauma to perineum and vulva during delivery
C0269863|T037|HT|664.0|ICD9CM|First-degree perineal laceration during delivery|First-degree perineal laceration during delivery
C0157313|T037|AB|664.00|ICD9CM|Del w 1 deg lacerat-unsp|Del w 1 deg lacerat-unsp
C0157313|T037|PT|664.00|ICD9CM|First-degree perineal laceration, unspecified as to episode of care or not applicable|First-degree perineal laceration, unspecified as to episode of care or not applicable
C1812626|T037|AB|664.01|ICD9CM|Del w 1 deg lacerat-del|Del w 1 deg lacerat-del
C1812626|T037|PT|664.01|ICD9CM|First-degree perineal laceration, delivered, with or without mention of antepartum condition|First-degree perineal laceration, delivered, with or without mention of antepartum condition
C0157315|T037|AB|664.04|ICD9CM|Del w 1 deg lac-postpart|Del w 1 deg lac-postpart
C0157315|T037|PT|664.04|ICD9CM|First-degree perineal laceration, postpartum condition or complication|First-degree perineal laceration, postpartum condition or complication
C0269870|T037|HT|664.1|ICD9CM|Second-degree perineal laceration during delivery|Second-degree perineal laceration during delivery
C0157317|T037|AB|664.10|ICD9CM|Del w 2 deg lacerat-unsp|Del w 2 deg lacerat-unsp
C0157317|T037|PT|664.10|ICD9CM|Second-degree perineal laceration, unspecified as to episode of care or not applicable|Second-degree perineal laceration, unspecified as to episode of care or not applicable
C0269870|T037|AB|664.11|ICD9CM|Del w 2 deg lacerat-del|Del w 2 deg lacerat-del
C0269870|T037|PT|664.11|ICD9CM|Second-degree perineal laceration, delivered, with or without mention of antepartum condition|Second-degree perineal laceration, delivered, with or without mention of antepartum condition
C0490051|T037|AB|664.14|ICD9CM|Del w 2 deg lac-postpart|Del w 2 deg lac-postpart
C0490051|T037|PT|664.14|ICD9CM|Second-degree perineal laceration, postpartum condition or complication|Second-degree perineal laceration, postpartum condition or complication
C0269874|T037|HT|664.2|ICD9CM|Third-degree perineal laceration during delivery|Third-degree perineal laceration during delivery
C0157321|T037|AB|664.20|ICD9CM|Del w 3 deg lacerat-unsp|Del w 3 deg lacerat-unsp
C0157321|T037|PT|664.20|ICD9CM|Third-degree perineal laceration, unspecified as to episode of care or not applicable|Third-degree perineal laceration, unspecified as to episode of care or not applicable
C0269874|T037|AB|664.21|ICD9CM|Del w 3 deg lacerat-del|Del w 3 deg lacerat-del
C0269874|T037|PT|664.21|ICD9CM|Third-degree perineal laceration, delivered, with or without mention of antepartum condition|Third-degree perineal laceration, delivered, with or without mention of antepartum condition
C0157323|T037|AB|664.24|ICD9CM|Del w 3 deg lac-postpart|Del w 3 deg lac-postpart
C0157323|T037|PT|664.24|ICD9CM|Third-degree perineal laceration, postpartum condition or complication|Third-degree perineal laceration, postpartum condition or complication
C1275806|T033|HT|664.3|ICD9CM|Fourth-degree perineal laceration during delivery|Fourth-degree perineal laceration during delivery
C0157325|T037|AB|664.30|ICD9CM|Del w 4 deg lacerat-unsp|Del w 4 deg lacerat-unsp
C0157325|T037|PT|664.30|ICD9CM|Fourth-degree perineal laceration, unspecified as to episode of care or not applicable|Fourth-degree perineal laceration, unspecified as to episode of care or not applicable
C1275806|T033|AB|664.31|ICD9CM|Del w 4 deg lacerat-del|Del w 4 deg lacerat-del
C1275806|T033|PT|664.31|ICD9CM|Fourth-degree perineal laceration, delivered, with or without mention of antepartum condition|Fourth-degree perineal laceration, delivered, with or without mention of antepartum condition
C0157327|T037|AB|664.34|ICD9CM|Del w 4 deg lac-postpart|Del w 4 deg lac-postpart
C0157327|T037|PT|664.34|ICD9CM|Fourth-degree perineal laceration, postpartum condition or complication|Fourth-degree perineal laceration, postpartum condition or complication
C0269859|T037|HT|664.4|ICD9CM|Unspecified perineal laceration during delivery|Unspecified perineal laceration during delivery
C0157329|T047|AB|664.40|ICD9CM|Ob perineal lac NOS-unsp|Ob perineal lac NOS-unsp
C0157329|T047|PT|664.40|ICD9CM|Unspecified perineal laceration, unspecified as to episode of care or not applicable|Unspecified perineal laceration, unspecified as to episode of care or not applicable
C0269859|T037|AB|664.41|ICD9CM|Ob perineal lac NOS-del|Ob perineal lac NOS-del
C0269859|T037|PT|664.41|ICD9CM|Unspecified perineal laceration, delivered, with or without mention of antepartum condition|Unspecified perineal laceration, delivered, with or without mention of antepartum condition
C0157331|T037|AB|664.44|ICD9CM|Perineal lac NOS-postpar|Perineal lac NOS-postpar
C0157331|T037|PT|664.44|ICD9CM|Unspecified perineal laceration, postpartum condition or complication|Unspecified perineal laceration, postpartum condition or complication
C0157332|T037|HT|664.5|ICD9CM|Vulvar and perineal hematoma during delivery|Vulvar and perineal hematoma during delivery
C0157333|T047|AB|664.50|ICD9CM|Ob perineal hematom-unsp|Ob perineal hematom-unsp
C0157333|T047|PT|664.50|ICD9CM|Vulvar and perineal hematoma, unspecified as to episode of care or not applicable|Vulvar and perineal hematoma, unspecified as to episode of care or not applicable
C0157334|T047|AB|664.51|ICD9CM|Ob perineal hematoma-del|Ob perineal hematoma-del
C0157334|T047|PT|664.51|ICD9CM|Vulvar and perineal hematoma, delivered, with or without mention of antepartum condition|Vulvar and perineal hematoma, delivered, with or without mention of antepartum condition
C0157335|T047|AB|664.54|ICD9CM|Perin hematoma-postpart|Perin hematoma-postpart
C0157335|T047|PT|664.54|ICD9CM|Vulvar and perineal hematoma, postpartum condition or complication|Vulvar and perineal hematoma, postpartum condition or complication
C1955493|T047|HT|664.6|ICD9CM|Anal sphincter tear complicating delivery, not associated with third-degree perineal laceration|Anal sphincter tear complicating delivery, not associated with third-degree perineal laceration
C1955490|T047|AB|664.60|ICD9CM|Anal sphincter tear NOS|Anal sphincter tear NOS
C1955491|T047|AB|664.61|ICD9CM|Anal sphincter tear-del|Anal sphincter tear-del
C1955492|T047|AB|664.64|ICD9CM|Anal sphinctr tear w p/p|Anal sphinctr tear w p/p
C0157336|T037|HT|664.8|ICD9CM|Other specified trauma to perineum and vulva during delivery|Other specified trauma to perineum and vulva during delivery
C0157337|T037|AB|664.80|ICD9CM|Ob perin traum NEC-unsp|Ob perin traum NEC-unsp
C0157337|T037|PT|664.80|ICD9CM|Other specified trauma to perineum and vulva, unspecified as to episode of care or not applicable|Other specified trauma to perineum and vulva, unspecified as to episode of care or not applicable
C0157338|T037|AB|664.81|ICD9CM|Ob perineal trau NEC-del|Ob perineal trau NEC-del
C0157339|T037|PT|664.84|ICD9CM|Other specified trauma to perineum and vulva, postpartum condition or complication|Other specified trauma to perineum and vulva, postpartum condition or complication
C0157339|T037|AB|664.84|ICD9CM|Perin traum NEC-postpart|Perin traum NEC-postpart
C0157340|T037|HT|664.9|ICD9CM|Unspecified trauma to perineum and vulva during delivery|Unspecified trauma to perineum and vulva during delivery
C0157341|T037|AB|664.90|ICD9CM|Ob perin traum NOS-unsp|Ob perin traum NOS-unsp
C0157341|T037|PT|664.90|ICD9CM|Unspecified trauma to perineum and vulva, unspecified as to episode of care or not applicable|Unspecified trauma to perineum and vulva, unspecified as to episode of care or not applicable
C0157342|T037|AB|664.91|ICD9CM|Ob perineal trau NOS-del|Ob perineal trau NOS-del
C0157342|T037|PT|664.91|ICD9CM|Unspecified trauma to perineum and vulva, delivered, with or without mention of antepartum condition|Unspecified trauma to perineum and vulva, delivered, with or without mention of antepartum condition
C0157343|T037|AB|664.94|ICD9CM|Perin traum NOS-postpart|Perin traum NOS-postpart
C0157343|T037|PT|664.94|ICD9CM|Unspecified trauma to perineum and vulva, postpartum condition or complication|Unspecified trauma to perineum and vulva, postpartum condition or complication
C0157344|T037|HT|665|ICD9CM|Other obstetrical trauma|Other obstetrical trauma
C0157345|T037|HT|665.0|ICD9CM|Rupture of uterus before onset of labor|Rupture of uterus before onset of labor
C0157346|T047|AB|665.00|ICD9CM|Prelabor rupt uter-unsp|Prelabor rupt uter-unsp
C0157346|T047|PT|665.00|ICD9CM|Rupture of uterus before onset of labor, unspecified as to episode of care or not applicable|Rupture of uterus before onset of labor, unspecified as to episode of care or not applicable
C0157347|T046|AB|665.01|ICD9CM|Prelabor rupt uterus-del|Prelabor rupt uterus-del
C0157347|T046|PT|665.01|ICD9CM|Rupture of uterus before onset of labor, delivered, with or without mention of antepartum condition|Rupture of uterus before onset of labor, delivered, with or without mention of antepartum condition
C1812625|T047|AB|665.03|ICD9CM|Prelab rupt uter-antepar|Prelab rupt uter-antepar
C1812625|T047|PT|665.03|ICD9CM|Rupture of uterus before onset of labor, antepartum condition or complication|Rupture of uterus before onset of labor, antepartum condition or complication
C3812903|T046|HT|665.1|ICD9CM|Rupture of uterus during labor|Rupture of uterus during labor
C0157350|T037|PT|665.10|ICD9CM|Rupture of uterus during labor, unspecified as to episode of care or not applicable|Rupture of uterus during labor, unspecified as to episode of care or not applicable
C0157350|T037|AB|665.10|ICD9CM|Rupture uterus NOS-unsp|Rupture uterus NOS-unsp
C0157351|T037|PT|665.11|ICD9CM|Rupture of uterus during labor, delivered, with or without mention of antepartum condition|Rupture of uterus during labor, delivered, with or without mention of antepartum condition
C0157351|T037|AB|665.11|ICD9CM|Rupture uterus NOS-deliv|Rupture uterus NOS-deliv
C0162482|T046|HT|665.2|ICD9CM|Obstetrical inversion of uterus|Obstetrical inversion of uterus
C0157355|T047|AB|665.20|ICD9CM|Inversion of uterus-unsp|Inversion of uterus-unsp
C0157355|T047|PT|665.20|ICD9CM|Inversion of uterus, unspecified as to episode of care or not applicable|Inversion of uterus, unspecified as to episode of care or not applicable
C0157356|T047|AB|665.22|ICD9CM|Invers uterus-del w p/p|Invers uterus-del w p/p
C0157356|T047|PT|665.22|ICD9CM|Inversion of uterus, delivered, with mention of postpartum complication|Inversion of uterus, delivered, with mention of postpartum complication
C0157357|T046|AB|665.24|ICD9CM|Invers uterus-postpart|Invers uterus-postpart
C0157357|T046|PT|665.24|ICD9CM|Inversion of uterus, postpartum condition or complication|Inversion of uterus, postpartum condition or complication
C0157358|T037|HT|665.3|ICD9CM|Obstetrical laceration of cervix|Obstetrical laceration of cervix
C0157359|T047|AB|665.30|ICD9CM|Lacerat of cervix-unspec|Lacerat of cervix-unspec
C0157359|T047|PT|665.30|ICD9CM|Laceration of cervix, unspecified as to episode of care or not applicable|Laceration of cervix, unspecified as to episode of care or not applicable
C0157358|T037|AB|665.31|ICD9CM|Lacerat of cervix-deliv|Lacerat of cervix-deliv
C0157358|T037|PT|665.31|ICD9CM|Laceration of cervix, delivered, with or without mention of antepartum condition|Laceration of cervix, delivered, with or without mention of antepartum condition
C0157361|T047|AB|665.34|ICD9CM|Lacer of cervix-postpart|Lacer of cervix-postpart
C0157361|T047|PT|665.34|ICD9CM|Laceration of cervix, postpartum condition or complication|Laceration of cervix, postpartum condition or complication
C0157362|T037|HT|665.4|ICD9CM|High vaginal laceration during and after labor|High vaginal laceration during and after labor
C0157363|T047|AB|665.40|ICD9CM|High vaginal lacer-unsp|High vaginal lacer-unsp
C0157363|T047|PT|665.40|ICD9CM|High vaginal laceration, unspecified as to episode of care or not applicable|High vaginal laceration, unspecified as to episode of care or not applicable
C0157364|T037|AB|665.41|ICD9CM|High vaginal lacer-deliv|High vaginal lacer-deliv
C0157364|T037|PT|665.41|ICD9CM|High vaginal laceration, delivered, with or without mention of antepartum condition|High vaginal laceration, delivered, with or without mention of antepartum condition
C0157365|T037|AB|665.44|ICD9CM|High vaginal lac-postpar|High vaginal lac-postpar
C0157365|T037|PT|665.44|ICD9CM|High vaginal laceration, postpartum condition or complication|High vaginal laceration, postpartum condition or complication
C0157366|T037|HT|665.5|ICD9CM|Other obstetrical injury to pelvic organs|Other obstetrical injury to pelvic organs
C0157367|T037|AB|665.50|ICD9CM|Ob inj pelv org NEC-unsp|Ob inj pelv org NEC-unsp
C0157367|T037|PT|665.50|ICD9CM|Other injury to pelvic organs, unspecified as to episode of care or not applicable|Other injury to pelvic organs, unspecified as to episode of care or not applicable
C0157368|T037|AB|665.51|ICD9CM|Ob inj pelv org NEC-del|Ob inj pelv org NEC-del
C0157368|T037|PT|665.51|ICD9CM|Other injury to pelvic organs, delivered, with or without mention of antepartum condition|Other injury to pelvic organs, delivered, with or without mention of antepartum condition
C0157369|T037|AB|665.54|ICD9CM|Inj pelv org NEC-postpar|Inj pelv org NEC-postpar
C0157369|T037|PT|665.54|ICD9CM|Other injury to pelvic organs, postpartum condition or complication|Other injury to pelvic organs, postpartum condition or complication
C0269891|T037|HT|665.6|ICD9CM|Obstetrical damage to pelvic joints and ligaments|Obstetrical damage to pelvic joints and ligaments
C0157371|T037|PT|665.60|ICD9CM|Damage to pelvic joints and ligaments, unspecified as to episode of care or not applicable|Damage to pelvic joints and ligaments, unspecified as to episode of care or not applicable
C0157371|T037|AB|665.60|ICD9CM|Damage to pelvic jt-unsp|Damage to pelvic jt-unsp
C0269891|T037|PT|665.61|ICD9CM|Damage to pelvic joints and ligaments, delivered, with or without mention of antepartum condition|Damage to pelvic joints and ligaments, delivered, with or without mention of antepartum condition
C0269891|T037|AB|665.61|ICD9CM|Damage to pelvic jt-del|Damage to pelvic jt-del
C0157373|T037|AB|665.64|ICD9CM|Damage pelvic jt-postpar|Damage pelvic jt-postpar
C0157373|T037|PT|665.64|ICD9CM|Damage to pelvic joints and ligaments, postpartum condition or complication|Damage to pelvic joints and ligaments, postpartum condition or complication
C0269895|T046|HT|665.7|ICD9CM|Obstetrical pelvic hematoma|Obstetrical pelvic hematoma
C0157375|T047|AB|665.70|ICD9CM|Ob pelvic hematoma-unsp|Ob pelvic hematoma-unsp
C0157375|T047|PT|665.70|ICD9CM|Pelvic hematoma, unspecified as to episode of care or not applicable|Pelvic hematoma, unspecified as to episode of care or not applicable
C0269895|T046|AB|665.71|ICD9CM|Ob pelvic hematoma-deliv|Ob pelvic hematoma-deliv
C0269895|T046|PT|665.71|ICD9CM|Pelvic hematoma, delivered, with or without mention of antepartum condition|Pelvic hematoma, delivered, with or without mention of antepartum condition
C0157377|T047|AB|665.72|ICD9CM|Pelvic hematom-del w pp|Pelvic hematom-del w pp
C0157377|T047|PT|665.72|ICD9CM|Pelvic hematoma, delivered with mention of postpartum complication|Pelvic hematoma, delivered with mention of postpartum complication
C0157378|T047|AB|665.74|ICD9CM|Pelvic hematoma-postpart|Pelvic hematoma-postpart
C0157378|T047|PT|665.74|ICD9CM|Pelvic hematoma, postpartum condition or complication|Pelvic hematoma, postpartum condition or complication
C0157379|T037|HT|665.8|ICD9CM|Other specified obstetrical trauma|Other specified obstetrical trauma
C0157380|T037|AB|665.80|ICD9CM|Ob trauma NEC-unspec|Ob trauma NEC-unspec
C0157380|T037|PT|665.80|ICD9CM|Other specified obstetrical trauma, unspecified as to episode of care or not applicable|Other specified obstetrical trauma, unspecified as to episode of care or not applicable
C0157381|T037|AB|665.81|ICD9CM|Ob trauma NEC-delivered|Ob trauma NEC-delivered
C0157381|T037|PT|665.81|ICD9CM|Other specified obstetrical trauma, delivered, with or without mention of antepartum condition|Other specified obstetrical trauma, delivered, with or without mention of antepartum condition
C0157382|T037|AB|665.82|ICD9CM|Ob trauma NEC-del w p/p|Ob trauma NEC-del w p/p
C0157382|T037|PT|665.82|ICD9CM|Other specified obstetrical trauma, delivered, with mention of postpartum complication|Other specified obstetrical trauma, delivered, with mention of postpartum complication
C0157383|T037|AB|665.83|ICD9CM|Ob trauma NEC-antepartum|Ob trauma NEC-antepartum
C0157383|T037|PT|665.83|ICD9CM|Other specified obstetrical trauma, antepartum condition or complication|Other specified obstetrical trauma, antepartum condition or complication
C0157384|T037|AB|665.84|ICD9CM|Ob trauma NEC-postpartum|Ob trauma NEC-postpartum
C0157384|T037|PT|665.84|ICD9CM|Other specified obstetrical trauma, postpartum condition or complication|Other specified obstetrical trauma, postpartum condition or complication
C0269858|T037|HT|665.9|ICD9CM|Unspecified obstetrical trauma|Unspecified obstetrical trauma
C0157386|T037|AB|665.90|ICD9CM|Ob trauma NOS-unspec|Ob trauma NOS-unspec
C0157386|T037|PT|665.90|ICD9CM|Unspecified obstetrical trauma, unspecified as to episode of care or not applicable|Unspecified obstetrical trauma, unspecified as to episode of care or not applicable
C0157387|T037|AB|665.91|ICD9CM|Ob trauma NOS-delivered|Ob trauma NOS-delivered
C0157387|T037|PT|665.91|ICD9CM|Unspecified obstetrical trauma, delivered, with or without mention of antepartum condition|Unspecified obstetrical trauma, delivered, with or without mention of antepartum condition
C0157388|T037|AB|665.92|ICD9CM|Ob trauma NOS-del w p/p|Ob trauma NOS-del w p/p
C0157388|T037|PT|665.92|ICD9CM|Unspecified obstetrical trauma, delivered, with mention of postpartum complication|Unspecified obstetrical trauma, delivered, with mention of postpartum complication
C0157389|T037|AB|665.93|ICD9CM|Ob trauma NOS-antepartum|Ob trauma NOS-antepartum
C0157389|T037|PT|665.93|ICD9CM|Unspecified obstetrical trauma, antepartum condition or complication|Unspecified obstetrical trauma, antepartum condition or complication
C0157390|T037|AB|665.94|ICD9CM|Ob trauma NOS-postpartum|Ob trauma NOS-postpartum
C0157390|T037|PT|665.94|ICD9CM|Unspecified obstetrical trauma, postpartum condition or complication|Unspecified obstetrical trauma, postpartum condition or complication
C0032797|T046|HT|666|ICD9CM|Postpartum hemorrhage|Postpartum hemorrhage
C0269898|T046|HT|666.0|ICD9CM|Third-stage postpartum hemorrhage|Third-stage postpartum hemorrhage
C0157392|T037|AB|666.00|ICD9CM|Third-stage hem-unspec|Third-stage hem-unspec
C0157392|T037|PT|666.00|ICD9CM|Third-stage postpartum hemorrhage, unspecified as to episode of care or not applicable|Third-stage postpartum hemorrhage, unspecified as to episode of care or not applicable
C0157393|T046|PT|666.02|ICD9CM|Third-stage postpartum hemorrhage, delivered, with mention of postpartum complication|Third-stage postpartum hemorrhage, delivered, with mention of postpartum complication
C0157393|T046|AB|666.02|ICD9CM|Thrd-stage hem-del w p/p|Thrd-stage hem-del w p/p
C0269898|T046|AB|666.04|ICD9CM|Third-stage hem-postpart|Third-stage hem-postpart
C0269898|T046|PT|666.04|ICD9CM|Third-stage postpartum hemorrhage, postpartum condition or complication|Third-stage postpartum hemorrhage, postpartum condition or complication
C0220887|T046|HT|666.1|ICD9CM|Other immediate postpartum hemorrhage|Other immediate postpartum hemorrhage
C0157394|T046|PT|666.10|ICD9CM|Other immediate postpartum hemorrhage, unspecified as to episode of care or not applicable|Other immediate postpartum hemorrhage, unspecified as to episode of care or not applicable
C0157394|T046|AB|666.10|ICD9CM|Postpartum hem NEC-unsp|Postpartum hem NEC-unsp
C0157395|T046|PT|666.12|ICD9CM|Other immediate postpartum hemorrhage, delivered, with mention of postpartum complication|Other immediate postpartum hemorrhage, delivered, with mention of postpartum complication
C0157395|T046|AB|666.12|ICD9CM|Postpa hem NEC-del w p/p|Postpa hem NEC-del w p/p
C0220887|T046|PT|666.14|ICD9CM|Other immediate postpartum hemorrhage, postpartum condition or complication|Other immediate postpartum hemorrhage, postpartum condition or complication
C0220887|T046|AB|666.14|ICD9CM|Postpart hem NEC-postpar|Postpart hem NEC-postpar
C0473508|T046|HT|666.2|ICD9CM|Delayed and secondary postpartum hemorrhage|Delayed and secondary postpartum hemorrhage
C0473508|T046|AB|666.20|ICD9CM|Delay p/part hem-unspec|Delay p/part hem-unspec
C0473508|T046|PT|666.20|ICD9CM|Delayed and secondary postpartum hemorrhage, unspecified as to episode of care or not applicable|Delayed and secondary postpartum hemorrhage, unspecified as to episode of care or not applicable
C0157398|T047|AB|666.22|ICD9CM|Delay p/p hem-del w p/p|Delay p/p hem-del w p/p
C0157398|T047|PT|666.22|ICD9CM|Delayed and secondary postpartum hemorrhage, delivered, with mention of postpartum complication|Delayed and secondary postpartum hemorrhage, delivered, with mention of postpartum complication
C0473508|T046|AB|666.24|ICD9CM|Delay p/part hem-postpar|Delay p/part hem-postpar
C0473508|T046|PT|666.24|ICD9CM|Delayed and secondary postpartum hemorrhage, postpartum condition or complication|Delayed and secondary postpartum hemorrhage, postpartum condition or complication
C0157403|T047|HT|666.3|ICD9CM|Postpartum coagulation defects|Postpartum coagulation defects
C0157401|T047|AB|666.30|ICD9CM|Postpart coagul def-unsp|Postpart coagul def-unsp
C0157401|T047|PT|666.30|ICD9CM|Postpartum coagulation defects, unspecified as to episode of care or not applicable|Postpartum coagulation defects, unspecified as to episode of care or not applicable
C0157402|T047|AB|666.32|ICD9CM|P/p coag def-del w p/p|P/p coag def-del w p/p
C0157402|T047|PT|666.32|ICD9CM|Postpartum coagulation defects, delivered, with mention of postpartum complication|Postpartum coagulation defects, delivered, with mention of postpartum complication
C0157403|T047|AB|666.34|ICD9CM|Postpart coag def-postpa|Postpart coag def-postpa
C0157403|T047|PT|666.34|ICD9CM|Postpartum coagulation defects, postpartum condition or complication|Postpartum coagulation defects, postpartum condition or complication
C0157404|T046|HT|667|ICD9CM|Retained placenta or membranes, without hemorrhage|Retained placenta or membranes, without hemorrhage
C0269905|T046|HT|667.0|ICD9CM|Retained placenta without hemorrhage|Retained placenta without hemorrhage
C0157405|T047|AB|667.00|ICD9CM|Retain placenta NOS-unsp|Retain placenta NOS-unsp
C0157405|T047|PT|667.00|ICD9CM|Retained placenta without hemorrhage, unspecified as to episode of care or not applicable|Retained placenta without hemorrhage, unspecified as to episode of care or not applicable
C0157406|T047|PT|667.02|ICD9CM|Retained placenta without hemorrhage, delivered, with mention of postpartum complication|Retained placenta without hemorrhage, delivered, with mention of postpartum complication
C0157406|T047|AB|667.02|ICD9CM|Retnd plac NOS-del w p/p|Retnd plac NOS-del w p/p
C0157407|T047|AB|667.04|ICD9CM|Retain plac NOS-postpart|Retain plac NOS-postpart
C0157407|T047|PT|667.04|ICD9CM|Retained placenta without hemorrhage, postpartum condition or complication|Retained placenta without hemorrhage, postpartum condition or complication
C0157408|T046|HT|667.1|ICD9CM|Retained portions of placenta or membranes, without hemorrhage|Retained portions of placenta or membranes, without hemorrhage
C0157409|T047|AB|667.10|ICD9CM|Retain prod concept-unsp|Retain prod concept-unsp
C0157410|T047|AB|667.12|ICD9CM|Ret prod conc-del w p/p|Ret prod conc-del w p/p
C0157411|T047|AB|667.14|ICD9CM|Ret prod concept-postpar|Ret prod concept-postpar
C0157411|T047|PT|667.14|ICD9CM|Retained portions of placenta or membranes, without hemorrhage, postpartum condition or complication|Retained portions of placenta or membranes, without hemorrhage, postpartum condition or complication
C0157412|T046|HT|668|ICD9CM|Complications of the administration of anesthetic or other sedation in labor and delivery|Complications of the administration of anesthetic or other sedation in labor and delivery
C0157413|T037|HT|668.0|ICD9CM|Pulmonary complications of anesthesia or other sedation in labor and delivery|Pulmonary complications of anesthesia or other sedation in labor and delivery
C0157414|T047|AB|668.00|ICD9CM|Pulm compl in del-unspec|Pulm compl in del-unspec
C0157415|T047|AB|668.01|ICD9CM|Pulm compl in del-deliv|Pulm compl in del-deliv
C0157416|T047|AB|668.02|ICD9CM|Pulm complic-del w p/p|Pulm complic-del w p/p
C0157417|T047|AB|668.03|ICD9CM|Pulm complicat-antepart|Pulm complicat-antepart
C0157418|T047|AB|668.04|ICD9CM|Pulm complicat-postpart|Pulm complicat-postpart
C0269916|T046|HT|668.1|ICD9CM|Cardiac complications of anesthesia or other sedation in labor and delivery|Cardiac complications of anesthesia or other sedation in labor and delivery
C0157420|T047|AB|668.10|ICD9CM|Heart compl in del-unsp|Heart compl in del-unsp
C0157421|T047|AB|668.11|ICD9CM|Heart compl in del-deliv|Heart compl in del-deliv
C0157422|T047|AB|668.12|ICD9CM|Heart compl-del w p/p|Heart compl-del w p/p
C0157423|T047|AB|668.13|ICD9CM|Heart complic-antepart|Heart complic-antepart
C0157424|T047|AB|668.14|ICD9CM|Heart complic-postpart|Heart complic-postpart
C0157425|T046|HT|668.2|ICD9CM|Central nervous system complications of anesthesia or other sedation in labor and delivery|Central nervous system complications of anesthesia or other sedation in labor and delivery
C0157426|T037|AB|668.20|ICD9CM|Cns compl labor/del-unsp|Cns compl labor/del-unsp
C0157427|T047|AB|668.21|ICD9CM|Cns compl lab/del-deliv|Cns compl lab/del-deliv
C0157428|T037|AB|668.22|ICD9CM|Cns complic-del w p/p|Cns complic-del w p/p
C0157429|T047|AB|668.23|ICD9CM|Cns compl in del-antepar|Cns compl in del-antepar
C0157430|T047|AB|668.24|ICD9CM|Cns compl in del-postpar|Cns compl in del-postpar
C0157431|T046|HT|668.8|ICD9CM|Other complications of anesthesia or other sedation in labor and delivery|Other complications of anesthesia or other sedation in labor and delivery
C0157432|T037|AB|668.80|ICD9CM|Anesth comp del NEC-unsp|Anesth comp del NEC-unsp
C0157436|T037|AB|668.81|ICD9CM|Anesth compl NEC-deliver|Anesth compl NEC-deliver
C0157434|T037|AB|668.82|ICD9CM|Anesth compl NEC-del p/p|Anesth compl NEC-del p/p
C0157435|T037|AB|668.83|ICD9CM|Anesth compl antepartum|Anesth compl antepartum
C0157436|T037|AB|668.84|ICD9CM|Anesth compl-postpartum|Anesth compl-postpartum
C0157437|T033|HT|668.9|ICD9CM|Unspecified complication of anesthesia or other sedation in labor and delivery|Unspecified complication of anesthesia or other sedation in labor and delivery
C0157438|T037|AB|668.90|ICD9CM|Anesth comp del NOS-unsp|Anesth comp del NOS-unsp
C0157439|T037|AB|668.91|ICD9CM|Anesth compl NOS-deliver|Anesth compl NOS-deliver
C0157440|T037|AB|668.92|ICD9CM|Anesth compl NOS-del p/p|Anesth compl NOS-del p/p
C0157441|T037|AB|668.93|ICD9CM|Anesth compl-antepartum|Anesth compl-antepartum
C0157442|T037|AB|668.94|ICD9CM|Anesth compl-postpartum|Anesth compl-postpartum
C0868755|T046|HT|669|ICD9CM|Other complications of labor and delivery, not elsewhere classified|Other complications of labor and delivery, not elsewhere classified
C0473485|T046|HT|669.0|ICD9CM|Maternal distress|Maternal distress
C0157445|T047|AB|669.00|ICD9CM|Maternal distress-unspec|Maternal distress-unspec
C0157446|T047|AB|669.01|ICD9CM|Maternal distress-deliv|Maternal distress-deliv
C0157447|T047|AB|669.02|ICD9CM|Matern distres-del w p/p|Matern distres-del w p/p
C0157448|T047|AB|669.03|ICD9CM|Matern distress-antepar|Matern distress-antepar
C0157448|T047|PT|669.03|ICD9CM|Maternal distress complicating labor and delivery, antepartum condition or complication|Maternal distress complicating labor and delivery, antepartum condition or complication
C0157449|T047|AB|669.04|ICD9CM|Matern distress-postpart|Matern distress-postpart
C0157449|T047|PT|669.04|ICD9CM|Maternal distress complicating labor and delivery, postpartum condition or complication|Maternal distress complicating labor and delivery, postpartum condition or complication
C0157450|T046|HT|669.1|ICD9CM|Shock during or following labor and delivery|Shock during or following labor and delivery
C0157451|T047|AB|669.10|ICD9CM|Obstetric shock-unspec|Obstetric shock-unspec
C0157451|T047|PT|669.10|ICD9CM|Shock during or following labor and delivery, unspecified as to episode of care or not applicable|Shock during or following labor and delivery, unspecified as to episode of care or not applicable
C0157452|T047|AB|669.11|ICD9CM|Obstetric shock-deliver|Obstetric shock-deliver
C0157453|T047|AB|669.12|ICD9CM|Obstet shock-deliv w p/p|Obstet shock-deliv w p/p
C0157453|T047|PT|669.12|ICD9CM|Shock during or following labor and delivery, delivered, with mention of postpartum complication|Shock during or following labor and delivery, delivered, with mention of postpartum complication
C0157454|T047|AB|669.13|ICD9CM|Obstetric shock-antepar|Obstetric shock-antepar
C0157454|T047|PT|669.13|ICD9CM|Shock during or following labor and delivery, antepartum condition or complication|Shock during or following labor and delivery, antepartum condition or complication
C0157455|T047|AB|669.14|ICD9CM|Obstetric shock-postpart|Obstetric shock-postpart
C0157455|T047|PT|669.14|ICD9CM|Shock during or following labor and delivery, postpartum condition or complication|Shock during or following labor and delivery, postpartum condition or complication
C0341966|T046|HT|669.2|ICD9CM|Maternal hypotension syndrome|Maternal hypotension syndrome
C0157456|T047|AB|669.20|ICD9CM|Matern hypotens syn-unsp|Matern hypotens syn-unsp
C0157456|T047|PT|669.20|ICD9CM|Maternal hypotension syndrome, unspecified as to episode of care or not applicable|Maternal hypotension syndrome, unspecified as to episode of care or not applicable
C0157457|T047|AB|669.21|ICD9CM|Matern hypoten syn-deliv|Matern hypoten syn-deliv
C0157457|T047|PT|669.21|ICD9CM|Maternal hypotension syndrome, delivered, with or without mention of antepartum condition|Maternal hypotension syndrome, delivered, with or without mention of antepartum condition
C0157458|T047|AB|669.22|ICD9CM|Matern hypoten-del w p/p|Matern hypoten-del w p/p
C0157458|T047|PT|669.22|ICD9CM|Maternal hypotension syndrome, delivered, with mention of postpartum complication|Maternal hypotension syndrome, delivered, with mention of postpartum complication
C0157459|T047|AB|669.23|ICD9CM|Matern hypotens-antepar|Matern hypotens-antepar
C0157459|T047|PT|669.23|ICD9CM|Maternal hypotension syndrome, antepartum condition or complication|Maternal hypotension syndrome, antepartum condition or complication
C0157460|T047|AB|669.24|ICD9CM|Matern hypotens-postpart|Matern hypotens-postpart
C0157460|T047|PT|669.24|ICD9CM|Maternal hypotension syndrome, postpartum condition or complication|Maternal hypotension syndrome, postpartum condition or complication
C2712851|T046|HT|669.3|ICD9CM|Acute kidney failure following labor and delivery|Acute kidney failure following labor and delivery
C0157462|T047|AB|669.30|ICD9CM|Ac kidny fail w del-unsp|Ac kidny fail w del-unsp
C0157463|T047|AB|669.32|ICD9CM|Ac kidney fail-del w p/p|Ac kidney fail-del w p/p
C0157464|T047|AB|669.34|ICD9CM|Ac kidney fail-postpart|Ac kidney fail-postpart
C0157464|T047|PT|669.34|ICD9CM|Acute kidney failure following labor and delivery, postpartum condition or complication|Acute kidney failure following labor and delivery, postpartum condition or complication
C0157465|T046|HT|669.4|ICD9CM|Other complications of obstetrical surgery and procedures|Other complications of obstetrical surgery and procedures
C0157466|T047|AB|669.40|ICD9CM|Oth ob surg compl-unspec|Oth ob surg compl-unspec
C0157467|T037|AB|669.41|ICD9CM|Oth ob compl-delivered|Oth ob compl-delivered
C0157468|T037|AB|669.42|ICD9CM|Oth ob compl-deliv w p/p|Oth ob compl-deliv w p/p
C0375475|T047|AB|669.43|ICD9CM|Complc ob surg anteprtm|Complc ob surg anteprtm
C0375475|T047|PT|669.43|ICD9CM|Other complications of obstetrical surgery and procedures, antepartum condition or complication|Other complications of obstetrical surgery and procedures, antepartum condition or complication
C0157469|T047|AB|669.44|ICD9CM|Oth ob surg compl-postpa|Oth ob surg compl-postpa
C0157469|T047|PT|669.44|ICD9CM|Other complications of obstetrical surgery and procedures, postpartum condition or complication|Other complications of obstetrical surgery and procedures, postpartum condition or complication
C0157443|T046|HT|669.8|ICD9CM|Other complications of labor and delivery|Other complications of labor and delivery
C0157479|T047|AB|669.80|ICD9CM|Compl lab/deliv NEC-unsp|Compl lab/deliv NEC-unsp
C0157479|T047|PT|669.80|ICD9CM|Other complications of labor and delivery, unspecified as to episode of care or not applicable|Other complications of labor and delivery, unspecified as to episode of care or not applicable
C0157480|T033|AB|669.81|ICD9CM|Comp lab/deliv NEC-deliv|Comp lab/deliv NEC-deliv
C0157481|T047|AB|669.82|ICD9CM|Compl del NEC-del w p/p|Compl del NEC-del w p/p
C0157481|T047|PT|669.82|ICD9CM|Other complications of labor and delivery, delivered, with mention of postpartum complication|Other complications of labor and delivery, delivered, with mention of postpartum complication
C0157482|T047|AB|669.83|ICD9CM|Compl deliv NEC-antepar|Compl deliv NEC-antepar
C0157482|T047|PT|669.83|ICD9CM|Other complications of labor and delivery, antepartum condition or complication|Other complications of labor and delivery, antepartum condition or complication
C0157483|T047|AB|669.84|ICD9CM|Compl deliv NEC-postpart|Compl deliv NEC-postpart
C0157483|T047|PT|669.84|ICD9CM|Other complications of labor and delivery, postpartum condition or complication|Other complications of labor and delivery, postpartum condition or complication
C0269815|T046|HT|669.9|ICD9CM|Unspecified complication of labor and delivery|Unspecified complication of labor and delivery
C0157484|T047|AB|669.90|ICD9CM|Compl lab/deliv NOS-unsp|Compl lab/deliv NOS-unsp
C0157484|T047|PT|669.90|ICD9CM|Unspecified complication of labor and delivery, unspecified as to episode of care or not applicable|Unspecified complication of labor and delivery, unspecified as to episode of care or not applicable
C0157485|T033|AB|669.91|ICD9CM|Comp lab/deliv NOS-deliv|Comp lab/deliv NOS-deliv
C0157486|T033|AB|669.92|ICD9CM|Compl del NOS-del w p/p|Compl del NOS-del w p/p
C0157486|T033|PT|669.92|ICD9CM|Unspecified complication of labor and delivery, delivered, with mention of postpartum complication|Unspecified complication of labor and delivery, delivered, with mention of postpartum complication
C0157487|T047|AB|669.93|ICD9CM|Compl deliv NOS-antepar|Compl deliv NOS-antepar
C0157487|T047|PT|669.93|ICD9CM|Unspecified complication of labor and delivery, antepartum condition or complication|Unspecified complication of labor and delivery, antepartum condition or complication
C0157488|T047|AB|669.94|ICD9CM|Compl deliv NOS-postpart|Compl deliv NOS-postpart
C0157488|T047|PT|669.94|ICD9CM|Unspecified complication of labor and delivery, postpartum condition or complication|Unspecified complication of labor and delivery, postpartum condition or complication
C0157489|T046|HT|670|ICD9CM|Major puerperal infection|Major puerperal infection
C0161972|T046|HT|670-677.99|ICD9CM|COMPLICATIONS OF THE PUERPERIUM|COMPLICATIONS OF THE PUERPERIUM
C0157489|T046|HT|670.0|ICD9CM|Major puerperal infection, unspecified|Major puerperal infection, unspecified
C0375476|T047|AB|670.00|ICD9CM|Maj puerp inf NOS-unsp|Maj puerp inf NOS-unsp
C0375476|T047|PT|670.00|ICD9CM|Major puerperal infection, unspecified as to episode of care or not applicable|Major puerperal infection, unspecified as to episode of care or not applicable
C0157491|T047|AB|670.02|ICD9CM|Maj puer inf NOS-del p/p|Maj puer inf NOS-del p/p
C0157491|T047|PT|670.02|ICD9CM|Major puerperal infection, delivered, with mention of postpartum complication|Major puerperal infection, delivered, with mention of postpartum complication
C0375477|T046|AB|670.04|ICD9CM|Major puerp inf NOS-p/p|Major puerp inf NOS-p/p
C0375477|T046|PT|670.04|ICD9CM|Major puerperal infection, postpartum condition or complication|Major puerperal infection, postpartum condition or complication
C0269932|T047|HT|670.1|ICD9CM|Puerperal endometritis|Puerperal endometritis
C2712345|T046|AB|670.10|ICD9CM|Puerp endometritis-unsp|Puerp endometritis-unsp
C2712345|T046|PT|670.10|ICD9CM|Puerperal endometritis, unspecified as to episode of care or not applicable|Puerperal endometritis, unspecified as to episode of care or not applicable
C2712346|T046|AB|670.12|ICD9CM|Puerp endomet del w p/p|Puerp endomet del w p/p
C2712346|T046|PT|670.12|ICD9CM|Puerperal endometritis, delivered, with mention of postpartum complication|Puerperal endometritis, delivered, with mention of postpartum complication
C2712347|T046|AB|670.14|ICD9CM|Puerp endomet-postpart|Puerp endomet-postpart
C2712347|T046|PT|670.14|ICD9CM|Puerperal endometritis, postpartum condition or complication|Puerperal endometritis, postpartum condition or complication
C0269936|T047|HT|670.2|ICD9CM|Puerperal sepsis|Puerperal sepsis
C2712348|T046|AB|670.20|ICD9CM|Puerperal sepsis-unsp|Puerperal sepsis-unsp
C2712348|T046|PT|670.20|ICD9CM|Puerperal sepsis, unspecified as to episode of care or not applicable|Puerperal sepsis, unspecified as to episode of care or not applicable
C2712349|T046|PT|670.22|ICD9CM|Puerperal sepsis, delivered, with mention of postpartum complication|Puerperal sepsis, delivered, with mention of postpartum complication
C2712349|T046|AB|670.22|ICD9CM|Puerprl sepsis-del w p/p|Puerprl sepsis-del w p/p
C2712350|T046|PT|670.24|ICD9CM|Puerperal sepsis, postpartum condition or complication|Puerperal sepsis, postpartum condition or complication
C2712350|T046|AB|670.24|ICD9CM|Puerperl sepsis-postpart|Puerperl sepsis-postpart
C2712615|T047|HT|670.3|ICD9CM|Puerperal septic thrombophlebitis|Puerperal septic thrombophlebitis
C2712351|T046|AB|670.30|ICD9CM|Puerp septc thromb-unsp|Puerp septc thromb-unsp
C2712351|T046|PT|670.30|ICD9CM|Puerperal septic thrombophlebitis, unspecified as to episode of care or not applicable|Puerperal septic thrombophlebitis, unspecified as to episode of care or not applicable
C2712352|T046|AB|670.32|ICD9CM|Prp sptc thrmb-del w p/p|Prp sptc thrmb-del w p/p
C2712352|T046|PT|670.32|ICD9CM|Puerperal septic thrombophlebitis, delivered, with mention of postpartum complication|Puerperal septic thrombophlebitis, delivered, with mention of postpartum complication
C2712353|T046|AB|670.34|ICD9CM|Prp septc thrmb-postpart|Prp septc thrmb-postpart
C2712353|T046|PT|670.34|ICD9CM|Puerperal septic thrombophlebitis, postpartum condition or complication|Puerperal septic thrombophlebitis, postpartum condition or complication
C2712902|T046|HT|670.8|ICD9CM|Other major puerperal infection|Other major puerperal infection
C2712354|T046|AB|670.80|ICD9CM|Maj prp infec NEC-unspec|Maj prp infec NEC-unspec
C2712354|T046|PT|670.80|ICD9CM|Other major puerperal infection, unspecified as to episode of care or not applicable|Other major puerperal infection, unspecified as to episode of care or not applicable
C2712355|T046|AB|670.82|ICD9CM|Maj prp inf NEC-dl w p/p|Maj prp inf NEC-dl w p/p
C2712355|T046|PT|670.82|ICD9CM|Other major puerperal infection, delivered, with mention of postpartum complication|Other major puerperal infection, delivered, with mention of postpartum complication
C2712356|T046|AB|670.84|ICD9CM|Maj puerp infec NEC-p/p|Maj puerp infec NEC-p/p
C2712356|T046|PT|670.84|ICD9CM|Other major puerperal infection, postpartum condition or complication|Other major puerperal infection, postpartum condition or complication
C0269945|T046|HT|671|ICD9CM|Venous complications in pregnancy and the puerperium|Venous complications in pregnancy and the puerperium
C0342068|T046|HT|671.0|ICD9CM|Varicose veins of legs in pregnancy and the puerperium|Varicose veins of legs in pregnancy and the puerperium
C0157495|T020|AB|671.00|ICD9CM|Varic vein leg preg-unsp|Varic vein leg preg-unsp
C0157496|T020|AB|671.01|ICD9CM|Varicose vein leg-deliv|Varicose vein leg-deliv
C0157497|T047|AB|671.02|ICD9CM|Varic vein leg-del w p/p|Varic vein leg-del w p/p
C0157498|T047|AB|671.03|ICD9CM|Varic vein leg-antepart|Varic vein leg-antepart
C0157499|T047|AB|671.04|ICD9CM|Varic vein leg-postpart|Varic vein leg-postpart
C2004479|T047|HT|671.1|ICD9CM|Varicose veins of vulva and perineum in pregnancy and the puerperium|Varicose veins of vulva and perineum in pregnancy and the puerperium
C0157501|T047|AB|671.10|ICD9CM|Varic vulva preg-unspec|Varic vulva preg-unspec
C0157502|T020|AB|671.11|ICD9CM|Varicose vulva-delivered|Varicose vulva-delivered
C0157503|T020|AB|671.12|ICD9CM|Varicose vulva-del w p/p|Varicose vulva-del w p/p
C0157504|T020|AB|671.13|ICD9CM|Varicose vulva-antepart|Varicose vulva-antepart
C0157505|T020|AB|671.14|ICD9CM|Varicose vulva-postpart|Varicose vulva-postpart
C0269951|T046|HT|671.2|ICD9CM|Superficial thrombophlebitis in pregnancy and the puerperium|Superficial thrombophlebitis in pregnancy and the puerperium
C0269951|T046|AB|671.20|ICD9CM|Thrombophleb preg-unspec|Thrombophleb preg-unspec
C0157508|T047|AB|671.21|ICD9CM|Thrombophlebitis-deliver|Thrombophlebitis-deliver
C0157509|T047|AB|671.22|ICD9CM|Thrombophleb-deliv w p/p|Thrombophleb-deliv w p/p
C0342054|T046|AB|671.23|ICD9CM|Thrombophlebit-antepart|Thrombophlebit-antepart
C0495289|T047|AB|671.24|ICD9CM|Thrombophlebit-postpart|Thrombophlebit-postpart
C0342044|T046|HT|671.3|ICD9CM|Deep phlebothrombosis, antepartum|Deep phlebothrombosis, antepartum
C0342044|T046|PT|671.30|ICD9CM|Deep phlebothrombosis, antepartum, unspecified as to episode of care or not applicable|Deep phlebothrombosis, antepartum, unspecified as to episode of care or not applicable
C0342044|T046|AB|671.30|ICD9CM|Deep thromb antepar-unsp|Deep thromb antepar-unsp
C0157514|T047|PT|671.31|ICD9CM|Deep phlebothrombosis, antepartum, delivered, with or without mention of antepartum condition|Deep phlebothrombosis, antepartum, delivered, with or without mention of antepartum condition
C0157514|T047|AB|671.31|ICD9CM|Deep throm antepar-deliv|Deep throm antepar-deliv
C0342044|T046|PT|671.33|ICD9CM|Deep phlebothrombosis, antepartum, antepartum condition or complication|Deep phlebothrombosis, antepartum, antepartum condition or complication
C0342044|T046|AB|671.33|ICD9CM|Deep vein thromb-antepar|Deep vein thromb-antepar
C0342039|T047|HT|671.4|ICD9CM|Deep phlebothrombosis, postpartum|Deep phlebothrombosis, postpartum
C0157516|T047|PT|671.40|ICD9CM|Deep phlebothrombosis, postpartum, unspecified as to episode of care or not applicable|Deep phlebothrombosis, postpartum, unspecified as to episode of care or not applicable
C0157516|T047|AB|671.40|ICD9CM|Deep thromb postpar-unsp|Deep thromb postpar-unsp
C0157517|T047|PT|671.42|ICD9CM|Deep phlebothrombosis, postpartum, delivered, with mention of postpartum complication|Deep phlebothrombosis, postpartum, delivered, with mention of postpartum complication
C0157517|T047|AB|671.42|ICD9CM|Thromb postpar-del w p/p|Thromb postpar-del w p/p
C0342039|T047|PT|671.44|ICD9CM|Deep phlebothrombosis, postpartum, postpartum condition or complication|Deep phlebothrombosis, postpartum, postpartum condition or complication
C0342039|T047|AB|671.44|ICD9CM|Deep vein thromb-postpar|Deep vein thromb-postpar
C0342038|T047|HT|671.5|ICD9CM|Other phlebitis and thrombosis in pregnancy and the puerperium|Other phlebitis and thrombosis in pregnancy and the puerperium
C0157519|T047|AB|671.50|ICD9CM|Thrombosis NEC preg-unsp|Thrombosis NEC preg-unsp
C0157520|T047|AB|671.51|ICD9CM|Thrombosis NEC-delivered|Thrombosis NEC-delivered
C0157521|T047|AB|671.52|ICD9CM|Thromb NEC-deliv w p/p|Thromb NEC-deliv w p/p
C0157522|T047|AB|671.53|ICD9CM|Thrombosis NEC-antepart|Thrombosis NEC-antepart
C0157523|T047|AB|671.54|ICD9CM|Thrombosis NEC-postpart|Thrombosis NEC-postpart
C0157524|T046|HT|671.8|ICD9CM|Other venous complications in pregnancy and the puerperium|Other venous complications in pregnancy and the puerperium
C0157525|T047|AB|671.80|ICD9CM|Ven compl preg NEC-unsp|Ven compl preg NEC-unsp
C0157526|T047|AB|671.81|ICD9CM|Venous compl NEC-deliver|Venous compl NEC-deliver
C0157527|T047|AB|671.82|ICD9CM|Ven comp NEC-deliv w p/p|Ven comp NEC-deliv w p/p
C0477814|T046|PT|671.83|ICD9CM|Other venous complications of pregnancy and the puerperium, antepartum condition or complication|Other venous complications of pregnancy and the puerperium, antepartum condition or complication
C0477814|T046|AB|671.83|ICD9CM|Venous compl NEC-antepar|Venous compl NEC-antepar
C0477869|T047|PT|671.84|ICD9CM|Other venous complications of pregnancy and the puerperium, postpartum condition or complication|Other venous complications of pregnancy and the puerperium, postpartum condition or complication
C0477869|T047|AB|671.84|ICD9CM|Venous compl NEC-postpar|Venous compl NEC-postpar
C0269945|T046|HT|671.9|ICD9CM|Unspecified venous complication in pregnancy and the puerperium|Unspecified venous complication in pregnancy and the puerperium
C0269945|T046|AB|671.90|ICD9CM|Ven compl preg NOS-unsp|Ven compl preg NOS-unsp
C0157532|T047|AB|671.91|ICD9CM|Venous compl NOS-deliver|Venous compl NOS-deliver
C0157533|T047|AB|671.92|ICD9CM|Ven comp NOS-deliv w p/p|Ven comp NOS-deliv w p/p
C0495184|T046|AB|671.93|ICD9CM|Venous compl NOS-antepar|Venous compl NOS-antepar
C0157535|T046|AB|671.94|ICD9CM|Venous compl NOS-postpar|Venous compl NOS-postpar
C0157536|T184|HT|672|ICD9CM|Pyrexia of unknown origin during the puerperium|Pyrexia of unknown origin during the puerperium
C0157536|T184|HT|672.0|ICD9CM|Pyrexia of unknown origin during the puerperium|Pyrexia of unknown origin during the puerperium
C1812621|T047|AB|672.00|ICD9CM|Puerperal pyrexia-unspec|Puerperal pyrexia-unspec
C1812621|T047|PT|672.00|ICD9CM|Pyrexia of unknown origin during the puerperium, unspecified as to episode of care or not applicable|Pyrexia of unknown origin during the puerperium, unspecified as to episode of care or not applicable
C0375478|T184|AB|672.02|ICD9CM|Puerp pyrexia-del w p/p|Puerp pyrexia-del w p/p
C0375478|T184|PT|672.02|ICD9CM|Pyrexia of unknown origin during the puerperium, delivered, with mention of postpartum complication|Pyrexia of unknown origin during the puerperium, delivered, with mention of postpartum complication
C0375479|T184|AB|672.04|ICD9CM|Puerp pyrexia-postpartum|Puerp pyrexia-postpartum
C0375479|T184|PT|672.04|ICD9CM|Pyrexia of unknown origin during the puerperium, postpartum condition or complication|Pyrexia of unknown origin during the puerperium, postpartum condition or complication
C0157540|T046|HT|673|ICD9CM|Obstetrical pulmonary embolism|Obstetrical pulmonary embolism
C0157541|T046|HT|673.0|ICD9CM|Obstetrical air embolism|Obstetrical air embolism
C0157542|T047|AB|673.00|ICD9CM|Ob air embolism-unspec|Ob air embolism-unspec
C0157542|T047|PT|673.00|ICD9CM|Obstetrical air embolism, unspecified as to episode of care or not applicable|Obstetrical air embolism, unspecified as to episode of care or not applicable
C0157543|T047|AB|673.01|ICD9CM|Ob air embolism-deliver|Ob air embolism-deliver
C0157543|T047|PT|673.01|ICD9CM|Obstetrical air embolism, delivered, with or without mention of antepartum condition|Obstetrical air embolism, delivered, with or without mention of antepartum condition
C0157544|T047|AB|673.02|ICD9CM|Ob air embol-deliv w p/p|Ob air embol-deliv w p/p
C0157544|T047|PT|673.02|ICD9CM|Obstetrical air embolism, delivered, with mention of postpartum complication|Obstetrical air embolism, delivered, with mention of postpartum complication
C0157545|T047|AB|673.03|ICD9CM|Ob air embolism-antepart|Ob air embolism-antepart
C0157545|T047|PT|673.03|ICD9CM|Obstetrical air embolism, antepartum condition or complication|Obstetrical air embolism, antepartum condition or complication
C0157546|T047|AB|673.04|ICD9CM|Ob air embolism-postpart|Ob air embolism-postpart
C0157546|T047|PT|673.04|ICD9CM|Obstetrical air embolism, postpartum condition or complication|Obstetrical air embolism, postpartum condition or complication
C0013927|T047|HT|673.1|ICD9CM|Amniotic fluid embolism|Amniotic fluid embolism
C0013927|T047|AB|673.10|ICD9CM|Amniotic embolism-unspec|Amniotic embolism-unspec
C0013927|T047|PT|673.10|ICD9CM|Amniotic fluid embolism, unspecified as to episode of care or not applicable|Amniotic fluid embolism, unspecified as to episode of care or not applicable
C0157548|T020|AB|673.11|ICD9CM|Amniotic embolism-deliv|Amniotic embolism-deliv
C0157548|T020|PT|673.11|ICD9CM|Amniotic fluid embolism, delivered, with or without mention of antepartum condition|Amniotic fluid embolism, delivered, with or without mention of antepartum condition
C0157549|T047|AB|673.12|ICD9CM|Amniot embol-deliv w p/p|Amniot embol-deliv w p/p
C0157549|T047|PT|673.12|ICD9CM|Amniotic fluid embolism, delivered, with mention of postpartum complication|Amniotic fluid embolism, delivered, with mention of postpartum complication
C0157550|T047|AB|673.13|ICD9CM|Amniotic embol-antepart|Amniotic embol-antepart
C0157550|T047|PT|673.13|ICD9CM|Amniotic fluid embolism, antepartum condition or complication|Amniotic fluid embolism, antepartum condition or complication
C0157551|T047|AB|673.14|ICD9CM|Amniotic embol-postpart|Amniotic embol-postpart
C0157551|T047|PT|673.14|ICD9CM|Amniotic fluid embolism, postpartum condition or complication|Amniotic fluid embolism, postpartum condition or complication
C0157552|T046|HT|673.2|ICD9CM|Obstetrical blood-clot embolism|Obstetrical blood-clot embolism
C0157552|T046|AB|673.20|ICD9CM|Ob pulm embol NOS-unspec|Ob pulm embol NOS-unspec
C0157552|T046|PT|673.20|ICD9CM|Obstetrical blood-clot embolism, unspecified as to episode of care or not applicable|Obstetrical blood-clot embolism, unspecified as to episode of care or not applicable
C0157554|T047|PT|673.21|ICD9CM|Obstetrical blood-clot embolism, delivered, with or without mention of antepartum condition|Obstetrical blood-clot embolism, delivered, with or without mention of antepartum condition
C0157554|T047|AB|673.21|ICD9CM|Pulm embol NOS-delivered|Pulm embol NOS-delivered
C0157555|T047|PT|673.22|ICD9CM|Obstetrical blood-clot embolism, delivered, with mention of postpartum complication|Obstetrical blood-clot embolism, delivered, with mention of postpartum complication
C0157555|T047|AB|673.22|ICD9CM|Pulm embol NOS-del w p/p|Pulm embol NOS-del w p/p
C0157556|T047|PT|673.23|ICD9CM|Obstetrical blood-clot embolism, antepartum condition or complication|Obstetrical blood-clot embolism, antepartum condition or complication
C0157556|T047|AB|673.23|ICD9CM|Pulm embol NOS-antepart|Pulm embol NOS-antepart
C0157557|T047|PT|673.24|ICD9CM|Obstetrical blood-clot embolism, postpartum condition or complication|Obstetrical blood-clot embolism, postpartum condition or complication
C0157557|T047|AB|673.24|ICD9CM|Pulm embol NOS-postpart|Pulm embol NOS-postpart
C0269959|T046|HT|673.3|ICD9CM|Obstetrical pyemic and septic embolism|Obstetrical pyemic and septic embolism
C0269959|T046|AB|673.30|ICD9CM|Ob pyemic embol-unspec|Ob pyemic embol-unspec
C0269959|T046|PT|673.30|ICD9CM|Obstetrical pyemic and septic embolism, unspecified as to episode of care or not applicable|Obstetrical pyemic and septic embolism, unspecified as to episode of care or not applicable
C0157560|T047|AB|673.31|ICD9CM|Ob pyemic embol-deliver|Ob pyemic embol-deliver
C0157560|T047|PT|673.31|ICD9CM|Obstetrical pyemic and septic embolism, delivered, with or without mention of antepartum condition|Obstetrical pyemic and septic embolism, delivered, with or without mention of antepartum condition
C0157561|T047|AB|673.32|ICD9CM|Ob pyem embol-del w p/p|Ob pyem embol-del w p/p
C0157561|T047|PT|673.32|ICD9CM|Obstetrical pyemic and septic embolism, delivered, with mention of postpartum complication|Obstetrical pyemic and septic embolism, delivered, with mention of postpartum complication
C0157562|T047|AB|673.33|ICD9CM|Ob pyemic embol-antepart|Ob pyemic embol-antepart
C0157562|T047|PT|673.33|ICD9CM|Obstetrical pyemic and septic embolism, antepartum condition or complication|Obstetrical pyemic and septic embolism, antepartum condition or complication
C0157563|T047|AB|673.34|ICD9CM|Ob pyemic embol-postpart|Ob pyemic embol-postpart
C0157563|T047|PT|673.34|ICD9CM|Obstetrical pyemic and septic embolism, postpartum condition or complication|Obstetrical pyemic and septic embolism, postpartum condition or complication
C0157564|T047|HT|673.8|ICD9CM|Other obstetrical pulmonary embolism|Other obstetrical pulmonary embolism
C0157565|T047|AB|673.80|ICD9CM|Ob pulmon embol NEC-unsp|Ob pulmon embol NEC-unsp
C0157565|T047|PT|673.80|ICD9CM|Other obstetrical pulmonary embolism, unspecified as to episode of care or not applicable|Other obstetrical pulmonary embolism, unspecified as to episode of care or not applicable
C0157566|T047|PT|673.81|ICD9CM|Other obstetrical pulmonary embolism, delivered, with or without mention of antepartum condition|Other obstetrical pulmonary embolism, delivered, with or without mention of antepartum condition
C0157566|T047|AB|673.81|ICD9CM|Pulmon embol NEC-deliver|Pulmon embol NEC-deliver
C0157567|T047|PT|673.82|ICD9CM|Other obstetrical pulmonary embolism, delivered, with mention of postpartum complication|Other obstetrical pulmonary embolism, delivered, with mention of postpartum complication
C0157567|T047|AB|673.82|ICD9CM|Pulm embol NEC-del w p/p|Pulm embol NEC-del w p/p
C0157568|T047|PT|673.83|ICD9CM|Other obstetrical pulmonary embolism, antepartum condition or complication|Other obstetrical pulmonary embolism, antepartum condition or complication
C0157568|T047|AB|673.83|ICD9CM|Pulmon embol NEC-antepar|Pulmon embol NEC-antepar
C0157569|T047|PT|673.84|ICD9CM|Other obstetrical pulmonary embolism, postpartum condition or complication|Other obstetrical pulmonary embolism, postpartum condition or complication
C0157569|T047|AB|673.84|ICD9CM|Pulmon embol NEC-postpar|Pulmon embol NEC-postpar
C0868855|T046|HT|674|ICD9CM|Other and unspecified complications of the puerperium, not elsewhere classified|Other and unspecified complications of the puerperium, not elsewhere classified
C0157571|T046|HT|674.0|ICD9CM|Cerebrovascular disorders in the puerperium|Cerebrovascular disorders in the puerperium
C0157572|T047|PT|674.00|ICD9CM|Cerebrovascular disorders in the puerperium, unspecified as to episode of care or not applicable|Cerebrovascular disorders in the puerperium, unspecified as to episode of care or not applicable
C0157572|T047|AB|674.00|ICD9CM|Puerp cerebvasc dis-unsp|Puerp cerebvasc dis-unsp
C0157573|T047|AB|674.01|ICD9CM|Puerp cerebvas dis-deliv|Puerp cerebvas dis-deliv
C0157574|T047|PT|674.02|ICD9CM|Cerebrovascular disorders in the puerperium, delivered, with mention of postpartum complication|Cerebrovascular disorders in the puerperium, delivered, with mention of postpartum complication
C0157574|T047|AB|674.02|ICD9CM|Cerebvas dis-deliv w p/p|Cerebvas dis-deliv w p/p
C0157575|T047|AB|674.03|ICD9CM|Cerebrovasc dis-antepart|Cerebrovasc dis-antepart
C0157575|T047|PT|674.03|ICD9CM|Cerebrovascular disorders in the puerperium, antepartum condition or complication|Cerebrovascular disorders in the puerperium, antepartum condition or complication
C1812627|T047|AB|674.04|ICD9CM|Cerebrovasc dis-postpart|Cerebrovasc dis-postpart
C1812627|T047|PT|674.04|ICD9CM|Cerebrovascular disorders in the puerperium, postpartum condition or complication|Cerebrovascular disorders in the puerperium, postpartum condition or complication
C3665608|T046|HT|674.1|ICD9CM|Disruption of cesarean wound|Disruption of cesarean wound
C0157578|T037|AB|674.10|ICD9CM|Disrupt c-sect wnd-unsp|Disrupt c-sect wnd-unsp
C0157578|T037|PT|674.10|ICD9CM|Disruption of cesarean wound, unspecified as to episode of care or not applicable|Disruption of cesarean wound, unspecified as to episode of care or not applicable
C0157579|T037|AB|674.12|ICD9CM|Disrupt c-sect-del w p/p|Disrupt c-sect-del w p/p
C0157579|T037|PT|674.12|ICD9CM|Disruption of cesarean wound, delivered, with mention of postpartum complication|Disruption of cesarean wound, delivered, with mention of postpartum complication
C1318514|T046|AB|674.14|ICD9CM|Disrupt c-sect-postpart|Disrupt c-sect-postpart
C1318514|T046|PT|674.14|ICD9CM|Disruption of cesarean wound, postpartum condition or complication|Disruption of cesarean wound, postpartum condition or complication
C3537063|T037|HT|674.2|ICD9CM|Disruption of obstetrical perineal wound|Disruption of obstetrical perineal wound
C0157582|T037|AB|674.20|ICD9CM|Disrupt perineum-unspec|Disrupt perineum-unspec
C0157582|T037|PT|674.20|ICD9CM|Disruption of perineal wound, unspecified as to episode of care or not applicable|Disruption of perineal wound, unspecified as to episode of care or not applicable
C0157583|T037|AB|674.22|ICD9CM|Disrupt perin-del w p/p|Disrupt perin-del w p/p
C0157583|T037|PT|674.22|ICD9CM|Disruption of perineal wound, delivered, with mention of postpartum complication|Disruption of perineal wound, delivered, with mention of postpartum complication
C3537063|T037|AB|674.24|ICD9CM|Disrupt perineum-postpar|Disrupt perineum-postpar
C3537063|T037|PT|674.24|ICD9CM|Disruption of perineal wound, postpartum condition or complication|Disruption of perineal wound, postpartum condition or complication
C0157585|T046|HT|674.3|ICD9CM|Other complications of obstetrical surgical wounds|Other complications of obstetrical surgical wounds
C0157586|T037|AB|674.30|ICD9CM|Ob surg compl NEC-unspec|Ob surg compl NEC-unspec
C0157587|T037|AB|674.32|ICD9CM|Ob surg compl-del w p/p|Ob surg compl-del w p/p
C0157588|T037|AB|674.34|ICD9CM|Ob surg comp NEC-postpar|Ob surg comp NEC-postpar
C0157588|T037|PT|674.34|ICD9CM|Other complications of obstetrical surgical wounds, postpartum condition or complication|Other complications of obstetrical surgical wounds, postpartum condition or complication
C0152437|T047|HT|674.4|ICD9CM|Placental polyp|Placental polyp
C0157589|T191|AB|674.40|ICD9CM|Placental polyp-unspec|Placental polyp-unspec
C0157589|T191|PT|674.40|ICD9CM|Placental polyp, unspecified as to episode of care or not applicable|Placental polyp, unspecified as to episode of care or not applicable
C0157590|T191|AB|674.42|ICD9CM|Placent polyp-del w p/p|Placent polyp-del w p/p
C0157590|T191|PT|674.42|ICD9CM|Placental polyp, delivered, with mention of postpartum complication|Placental polyp, delivered, with mention of postpartum complication
C0157591|T191|AB|674.44|ICD9CM|Placental polyp-postpart|Placental polyp-postpart
C0157591|T191|PT|674.44|ICD9CM|Placental polyp, postpartum condition or complication|Placental polyp, postpartum condition or complication
C0877208|T046|HT|674.5|ICD9CM|Peripartum cardiomyopathy|Peripartum cardiomyopathy
C1260427|T047|AB|674.50|ICD9CM|Peripart cardiomy-unspec|Peripart cardiomy-unspec
C1260427|T047|PT|674.50|ICD9CM|Peripartum cardiomyopathy, unspecified as to episode of care or not applicable|Peripartum cardiomyopathy, unspecified as to episode of care or not applicable
C1260428|T047|AB|674.51|ICD9CM|Peripartum cardiomy-del|Peripartum cardiomy-del
C1260428|T047|PT|674.51|ICD9CM|Peripartum cardiomyopathy, delivered, with or without mention of antepartum condition|Peripartum cardiomyopathy, delivered, with or without mention of antepartum condition
C1260429|T047|AB|674.52|ICD9CM|Peripart card del w p/p|Peripart card del w p/p
C1260429|T047|PT|674.52|ICD9CM|Peripartum cardiomyopathy, delivered, with mention of postpartum condition|Peripartum cardiomyopathy, delivered, with mention of postpartum condition
C1260430|T047|AB|674.53|ICD9CM|Peripartum card-antepart|Peripartum card-antepart
C1260430|T047|PT|674.53|ICD9CM|Peripartum cardiomyopathy, antepartum condition or complication|Peripartum cardiomyopathy, antepartum condition or complication
C1260431|T047|AB|674.54|ICD9CM|Peripartum card-postpart|Peripartum card-postpart
C1260431|T047|PT|674.54|ICD9CM|Peripartum cardiomyopathy, postpartum condition or complication|Peripartum cardiomyopathy, postpartum condition or complication
C0157592|T046|HT|674.8|ICD9CM|Other complications of the puerperium|Other complications of the puerperium
C2733633|T046|PT|674.80|ICD9CM|Other complications of puerperium, unspecified as to episode of care or not applicable|Other complications of puerperium, unspecified as to episode of care or not applicable
C2733633|T046|AB|674.80|ICD9CM|Puerp compl NEC-unspec|Puerp compl NEC-unspec
C0157594|T047|PT|674.82|ICD9CM|Other complications of puerperium, delivered, with mention of postpartum complication|Other complications of puerperium, delivered, with mention of postpartum complication
C0157594|T047|AB|674.82|ICD9CM|Puerp comp NEC-del w p/p|Puerp comp NEC-del w p/p
C2733634|T046|PT|674.84|ICD9CM|Other complications of puerperium, postpartum condition or complication|Other complications of puerperium, postpartum condition or complication
C2733634|T046|AB|674.84|ICD9CM|Puerp compl NEC-postpart|Puerp compl NEC-postpart
C0161972|T046|HT|674.9|ICD9CM|Unspecified complications of the puerperium|Unspecified complications of the puerperium
C0161972|T046|AB|674.90|ICD9CM|Puerp compl NOS-unspec|Puerp compl NOS-unspec
C0161972|T046|PT|674.90|ICD9CM|Unspecified complications of puerperium, unspecified as to episode of care or not applicable|Unspecified complications of puerperium, unspecified as to episode of care or not applicable
C0157597|T047|AB|674.92|ICD9CM|Puerp comp NOS-del w p/p|Puerp comp NOS-del w p/p
C0157597|T047|PT|674.92|ICD9CM|Unspecified complications of puerperium, delivered, with mention of postpartum complication|Unspecified complications of puerperium, delivered, with mention of postpartum complication
C0161972|T046|AB|674.94|ICD9CM|Puerp compl NOS-postpart|Puerp compl NOS-postpart
C0161972|T046|PT|674.94|ICD9CM|Unspecified complications of puerperium, postpartum condition or complication|Unspecified complications of puerperium, postpartum condition or complication
C0157623|T047|HT|675|ICD9CM|Infections of the breast and nipple associated with childbirth|Infections of the breast and nipple associated with childbirth
C0269979|T047|HT|675.0|ICD9CM|Infections of nipple associated with childbirth|Infections of nipple associated with childbirth
C0157600|T047|AB|675.00|ICD9CM|Infect nipple preg-unsp|Infect nipple preg-unsp
C0157600|T047|PT|675.00|ICD9CM|Infections of nipple associated with childbirth, unspecified as to episode of care or not applicable|Infections of nipple associated with childbirth, unspecified as to episode of care or not applicable
C0157601|T047|AB|675.01|ICD9CM|Infect nipple-delivered|Infect nipple-delivered
C0157602|T047|AB|675.02|ICD9CM|Infect nipple-del w p/p|Infect nipple-del w p/p
C0157602|T047|PT|675.02|ICD9CM|Infections of nipple associated with childbirth, delivered, with mention of postpartum complication|Infections of nipple associated with childbirth, delivered, with mention of postpartum complication
C0157603|T047|AB|675.03|ICD9CM|Infect nipple-antepartum|Infect nipple-antepartum
C0157603|T047|PT|675.03|ICD9CM|Infections of nipple associated with childbirth, antepartum condition or complication|Infections of nipple associated with childbirth, antepartum condition or complication
C0157604|T047|AB|675.04|ICD9CM|Infect nipple-postpartum|Infect nipple-postpartum
C0157604|T047|PT|675.04|ICD9CM|Infections of nipple associated with childbirth, postpartum condition or complication|Infections of nipple associated with childbirth, postpartum condition or complication
C0269981|T047|HT|675.1|ICD9CM|Abscess of breast associated with childbirth|Abscess of breast associated with childbirth
C0157606|T047|PT|675.10|ICD9CM|Abscess of breast associated with childbirth, unspecified as to episode of care or not applicable|Abscess of breast associated with childbirth, unspecified as to episode of care or not applicable
C0157606|T047|AB|675.10|ICD9CM|Breast abscess preg-unsp|Breast abscess preg-unsp
C0157607|T047|AB|675.11|ICD9CM|Breast abscess-delivered|Breast abscess-delivered
C0157608|T046|PT|675.12|ICD9CM|Abscess of breast associated with childbirth, delivered, with mention of postpartum complication|Abscess of breast associated with childbirth, delivered, with mention of postpartum complication
C0157608|T046|AB|675.12|ICD9CM|Breast abscess-del w p/p|Breast abscess-del w p/p
C0741646|T047|PT|675.13|ICD9CM|Abscess of breast associated with childbirth, antepartum condition or complication|Abscess of breast associated with childbirth, antepartum condition or complication
C0741646|T047|AB|675.13|ICD9CM|Breast abscess-antepart|Breast abscess-antepart
C0405309|T047|PT|675.14|ICD9CM|Abscess of breast associated with childbirth, postpartum condition or complication|Abscess of breast associated with childbirth, postpartum condition or complication
C0405309|T047|AB|675.14|ICD9CM|Breast abscess-postpart|Breast abscess-postpart
C0157611|T047|HT|675.2|ICD9CM|Nonpurulent mastitis associated with childbirth|Nonpurulent mastitis associated with childbirth
C0157612|T047|AB|675.20|ICD9CM|Mastitis in preg-unspec|Mastitis in preg-unspec
C0157612|T047|PT|675.20|ICD9CM|Nonpurulent mastitis associated with childbirth, unspecified as to episode of care or not applicable|Nonpurulent mastitis associated with childbirth, unspecified as to episode of care or not applicable
C0157613|T047|AB|675.21|ICD9CM|Mastitis-delivered|Mastitis-delivered
C0157614|T047|AB|675.22|ICD9CM|Mastitis-deliv w p/p|Mastitis-deliv w p/p
C0157614|T047|PT|675.22|ICD9CM|Nonpurulent mastitis associated with childbirth, delivered, with mention of postpartum complication|Nonpurulent mastitis associated with childbirth, delivered, with mention of postpartum complication
C1112795|T047|AB|675.23|ICD9CM|Mastitis-antepartum|Mastitis-antepartum
C1112795|T047|PT|675.23|ICD9CM|Nonpurulent mastitis associated with childbirth, antepartum condition or complication|Nonpurulent mastitis associated with childbirth, antepartum condition or complication
C1112702|T047|AB|675.24|ICD9CM|Mastitis-postpartum|Mastitis-postpartum
C1112702|T047|PT|675.24|ICD9CM|Nonpurulent mastitis associated with childbirth, postpartum condition or complication|Nonpurulent mastitis associated with childbirth, postpartum condition or complication
C0157617|T047|HT|675.8|ICD9CM|Other specified infections of the breast and nipple associated with childbirth|Other specified infections of the breast and nipple associated with childbirth
C0157618|T047|AB|675.80|ICD9CM|Breast inf preg NEC-unsp|Breast inf preg NEC-unsp
C0157619|T047|AB|675.81|ICD9CM|Breast infect NEC-deliv|Breast infect NEC-deliv
C0157620|T047|AB|675.82|ICD9CM|Breast inf NEC-del w p/p|Breast inf NEC-del w p/p
C0157621|T047|AB|675.83|ICD9CM|Breast inf NEC-antepart|Breast inf NEC-antepart
C0157622|T047|AB|675.84|ICD9CM|Breast inf NEC-postpart|Breast inf NEC-postpart
C0157623|T047|HT|675.9|ICD9CM|Unspecified infection of the breast and nipple associated with childbirth|Unspecified infection of the breast and nipple associated with childbirth
C0157624|T047|AB|675.90|ICD9CM|Breast inf preg NOS-unsp|Breast inf preg NOS-unsp
C0157625|T047|AB|675.91|ICD9CM|Breast infect NOS-deliv|Breast infect NOS-deliv
C0157626|T047|AB|675.92|ICD9CM|Breast inf NOS-del w p/p|Breast inf NOS-del w p/p
C0157627|T047|AB|675.93|ICD9CM|Breast inf NOS-antepart|Breast inf NOS-antepart
C0157628|T047|AB|675.94|ICD9CM|Breast inf NOS-postpart|Breast inf NOS-postpart
C0157629|T047|HT|676|ICD9CM|Other disorders of the breast associated with childbirth and disorders of lactation|Other disorders of the breast associated with childbirth and disorders of lactation
C0157630|T020|HT|676.0|ICD9CM|Retracted nipple associated with childbirth|Retracted nipple associated with childbirth
C0157631|T020|AB|676.00|ICD9CM|Retract nipple preg-unsp|Retract nipple preg-unsp
C0157631|T020|PT|676.00|ICD9CM|Retracted nipple associated with childbirth, unspecified as to episode of care or not applicable|Retracted nipple associated with childbirth, unspecified as to episode of care or not applicable
C0157632|T020|AB|676.01|ICD9CM|Retracted nipple-deliver|Retracted nipple-deliver
C0157633|T020|AB|676.02|ICD9CM|Retract nipple-del w p/p|Retract nipple-del w p/p
C0157633|T020|PT|676.02|ICD9CM|Retracted nipple associated with childbirth, delivered, with mention of postpartum complication|Retracted nipple associated with childbirth, delivered, with mention of postpartum complication
C0157634|T020|AB|676.03|ICD9CM|Retract nipple-antepart|Retract nipple-antepart
C0157634|T020|PT|676.03|ICD9CM|Retracted nipple associated with childbirth, antepartum condition or complication|Retracted nipple associated with childbirth, antepartum condition or complication
C0157635|T020|AB|676.04|ICD9CM|Retract nipple-postpart|Retract nipple-postpart
C0157635|T020|PT|676.04|ICD9CM|Retracted nipple associated with childbirth, postpartum condition or complication|Retracted nipple associated with childbirth, postpartum condition or complication
C0157636|T046|HT|676.1|ICD9CM|Cracked nipple associated with childbirth|Cracked nipple associated with childbirth
C0157637|T047|PT|676.10|ICD9CM|Cracked nipple associated with childbirth, unspecified as to episode of care or not applicable|Cracked nipple associated with childbirth, unspecified as to episode of care or not applicable
C0157637|T047|AB|676.10|ICD9CM|Cracked nipple preg-unsp|Cracked nipple preg-unsp
C0157638|T047|AB|676.11|ICD9CM|Cracked nipple-delivered|Cracked nipple-delivered
C0157639|T047|PT|676.12|ICD9CM|Cracked nipple associated with childbirth, delivered, with mention of postpartum complication|Cracked nipple associated with childbirth, delivered, with mention of postpartum complication
C0157639|T047|AB|676.12|ICD9CM|Cracked nipple-del w p/p|Cracked nipple-del w p/p
C0157640|T047|PT|676.13|ICD9CM|Cracked nipple associated with childbirth, antepartum condition or complication|Cracked nipple associated with childbirth, antepartum condition or complication
C0157640|T047|AB|676.13|ICD9CM|Cracked nipple-antepart|Cracked nipple-antepart
C0157641|T047|PT|676.14|ICD9CM|Cracked nipple associated with childbirth, postpartum condition or complication|Cracked nipple associated with childbirth, postpartum condition or complication
C0157641|T047|AB|676.14|ICD9CM|Cracked nipple-postpart|Cracked nipple-postpart
C0157642|T046|HT|676.2|ICD9CM|Engorgement of breasts associated with childbirth|Engorgement of breasts associated with childbirth
C0157643|T047|AB|676.20|ICD9CM|Breast engorge-unspec|Breast engorge-unspec
C0157644|T047|AB|676.21|ICD9CM|Breast engorge-delivered|Breast engorge-delivered
C0157645|T047|AB|676.22|ICD9CM|Breast engorge-del w p/p|Breast engorge-del w p/p
C0157646|T047|AB|676.23|ICD9CM|Breast engorge-antepart|Breast engorge-antepart
C0157646|T047|PT|676.23|ICD9CM|Engorgement of breasts associated with childbirth, antepartum condition or complication|Engorgement of breasts associated with childbirth, antepartum condition or complication
C0157647|T047|AB|676.24|ICD9CM|Breast engorge-postpart|Breast engorge-postpart
C0157647|T047|PT|676.24|ICD9CM|Engorgement of breasts associated with childbirth, postpartum condition or complication|Engorgement of breasts associated with childbirth, postpartum condition or complication
C0157648|T047|HT|676.3|ICD9CM|Other and unspecified disorder of breast associated with childbirth|Other and unspecified disorder of breast associated with childbirth
C0157649|T047|AB|676.30|ICD9CM|Breast dis preg NEC-unsp|Breast dis preg NEC-unsp
C0157650|T047|AB|676.31|ICD9CM|Breast dis NEC-delivered|Breast dis NEC-delivered
C0157651|T047|AB|676.32|ICD9CM|Breast dis NEC-del w p/p|Breast dis NEC-del w p/p
C0157652|T047|AB|676.33|ICD9CM|Breast dis NEC-antepart|Breast dis NEC-antepart
C0157653|T047|AB|676.34|ICD9CM|Breast dis NEC-postpart|Breast dis NEC-postpart
C0152158|T046|HT|676.4|ICD9CM|Failure of lactation|Failure of lactation
C0152158|T046|PT|676.40|ICD9CM|Failure of lactation, unspecified as to episode of care or not applicable|Failure of lactation, unspecified as to episode of care or not applicable
C0152158|T046|AB|676.40|ICD9CM|Lactation fail-unspec|Lactation fail-unspec
C0157655|T033|PT|676.41|ICD9CM|Failure of lactation, delivered, with or without mention of antepartum condition|Failure of lactation, delivered, with or without mention of antepartum condition
C0157655|T033|AB|676.41|ICD9CM|Lactation fail-delivered|Lactation fail-delivered
C0157656|T046|PT|676.42|ICD9CM|Failure of lactation, delivered, with mention of postpartum complication|Failure of lactation, delivered, with mention of postpartum complication
C0157656|T046|AB|676.42|ICD9CM|Lactation fail-del w p/p|Lactation fail-del w p/p
C0157657|T046|PT|676.43|ICD9CM|Failure of lactation, antepartum condition or complication|Failure of lactation, antepartum condition or complication
C0157657|T046|AB|676.43|ICD9CM|Lactation fail-antepart|Lactation fail-antepart
C0157656|T046|PT|676.44|ICD9CM|Failure of lactation, postpartum condition or complication|Failure of lactation, postpartum condition or complication
C0157656|T046|AB|676.44|ICD9CM|Lactation fail-postpart|Lactation fail-postpart
C0269993|T047|HT|676.5|ICD9CM|Suppressed lactation|Suppressed lactation
C0269993|T047|AB|676.50|ICD9CM|Suppr lactation-unspec|Suppr lactation-unspec
C0269993|T047|PT|676.50|ICD9CM|Suppressed lactation, unspecified as to episode of care or not applicable|Suppressed lactation, unspecified as to episode of care or not applicable
C0157660|T047|AB|676.51|ICD9CM|Suppr lactation-deliver|Suppr lactation-deliver
C0157660|T047|PT|676.51|ICD9CM|Suppressed lactation, delivered, with or without mention of antepartum condition|Suppressed lactation, delivered, with or without mention of antepartum condition
C0157661|T047|AB|676.52|ICD9CM|Suppr lactat-del w p/p|Suppr lactat-del w p/p
C0157661|T047|PT|676.52|ICD9CM|Suppressed lactation, delivered, with mention of postpartum complication|Suppressed lactation, delivered, with mention of postpartum complication
C0157662|T047|AB|676.53|ICD9CM|Suppr lactation-antepar|Suppr lactation-antepar
C0157662|T047|PT|676.53|ICD9CM|Suppressed lactation, antepartum condition or complication|Suppressed lactation, antepartum condition or complication
C0157661|T047|AB|676.54|ICD9CM|Suppr lactation-postpart|Suppr lactation-postpart
C0157661|T047|PT|676.54|ICD9CM|Suppressed lactation, postpartum condition or complication|Suppressed lactation, postpartum condition or complication
C0269995|T047|HT|676.6|ICD9CM|Galactorrhea|Galactorrhea
C0269995|T047|PT|676.60|ICD9CM|Galactorrhea associated with childbirth, unspecified as to episode of care or not applicable|Galactorrhea associated with childbirth, unspecified as to episode of care or not applicable
C0269995|T047|AB|676.60|ICD9CM|Galactorrhea preg-unspec|Galactorrhea preg-unspec
C0157665|T047|PT|676.61|ICD9CM|Galactorrhea associated with childbirth, delivered, with or without mention of antepartum condition|Galactorrhea associated with childbirth, delivered, with or without mention of antepartum condition
C0157665|T047|AB|676.61|ICD9CM|Galactorrhea-delivered|Galactorrhea-delivered
C0157666|T047|PT|676.62|ICD9CM|Galactorrhea associated with childbirth, delivered, with mention of postpartum complication|Galactorrhea associated with childbirth, delivered, with mention of postpartum complication
C0157666|T047|AB|676.62|ICD9CM|Galactorrhea-del w p/p|Galactorrhea-del w p/p
C0157667|T047|PT|676.63|ICD9CM|Galactorrhea associated with childbirth, antepartum condition or complication|Galactorrhea associated with childbirth, antepartum condition or complication
C0157667|T047|AB|676.63|ICD9CM|Galactorrhea-antepartum|Galactorrhea-antepartum
C0157668|T047|PT|676.64|ICD9CM|Galactorrhea associated with childbirth, postpartum condition or complication|Galactorrhea associated with childbirth, postpartum condition or complication
C0157668|T047|AB|676.64|ICD9CM|Galactorrhea-postpartum|Galactorrhea-postpartum
C0157669|T047|HT|676.8|ICD9CM|Other disorders of lactation|Other disorders of lactation
C0157669|T047|AB|676.80|ICD9CM|Lactation dis NEC-unspec|Lactation dis NEC-unspec
C0157669|T047|PT|676.80|ICD9CM|Other disorders of lactation, unspecified as to episode of care or not applicable|Other disorders of lactation, unspecified as to episode of care or not applicable
C0157671|T047|AB|676.81|ICD9CM|Lactation dis NEC-deliv|Lactation dis NEC-deliv
C0157671|T047|PT|676.81|ICD9CM|Other disorders of lactation, delivered, with or without mention of antepartum condition|Other disorders of lactation, delivered, with or without mention of antepartum condition
C0157672|T047|AB|676.82|ICD9CM|Lactat dis NEC-del w p/p|Lactat dis NEC-del w p/p
C0157672|T047|PT|676.82|ICD9CM|Other disorders of lactation, delivered, with mention of postpartum complication|Other disorders of lactation, delivered, with mention of postpartum complication
C0157673|T047|AB|676.83|ICD9CM|Lactat dis NEC-antepart|Lactat dis NEC-antepart
C0157673|T047|PT|676.83|ICD9CM|Other disorders of lactation, antepartum condition or complication|Other disorders of lactation, antepartum condition or complication
C0157672|T047|AB|676.84|ICD9CM|Lactat dis NEC-postpart|Lactat dis NEC-postpart
C0157672|T047|PT|676.84|ICD9CM|Other disorders of lactation, postpartum condition or complication|Other disorders of lactation, postpartum condition or complication
C0022927|T047|HT|676.9|ICD9CM|Unspecified disorder of lactation|Unspecified disorder of lactation
C0022927|T047|AB|676.90|ICD9CM|Lactation dis NOS-unspec|Lactation dis NOS-unspec
C0022927|T047|PT|676.90|ICD9CM|Unspecified disorder of lactation, unspecified as to episode of care or not applicable|Unspecified disorder of lactation, unspecified as to episode of care or not applicable
C0157676|T047|AB|676.91|ICD9CM|Lactation dis NOS-deliv|Lactation dis NOS-deliv
C0157676|T047|PT|676.91|ICD9CM|Unspecified disorder of lactation, delivered, with or without mention of antepartum condition|Unspecified disorder of lactation, delivered, with or without mention of antepartum condition
C0157677|T047|AB|676.92|ICD9CM|Lactat dis NOS-del w p/p|Lactat dis NOS-del w p/p
C0157677|T047|PT|676.92|ICD9CM|Unspecified disorder of lactation, delivered, with mention of postpartum complication|Unspecified disorder of lactation, delivered, with mention of postpartum complication
C0157678|T047|AB|676.93|ICD9CM|Lactat dis NOS-antepart|Lactat dis NOS-antepart
C0157678|T047|PT|676.93|ICD9CM|Unspecified disorder of lactation, antepartum condition or complication|Unspecified disorder of lactation, antepartum condition or complication
C0157679|T047|AB|676.94|ICD9CM|Lactat dis NOS-postpart|Lactat dis NOS-postpart
C0157679|T047|PT|676.94|ICD9CM|Unspecified disorder of lactation, postpartum condition or complication|Unspecified disorder of lactation, postpartum condition or complication
C0375480|T047|AB|677|ICD9CM|Late effct cmplcatn preg|Late effct cmplcatn preg
C0375480|T047|PT|677|ICD9CM|Late effect of complication of pregnancy, childbirth, and the puerperium|Late effect of complication of pregnancy, childbirth, and the puerperium
C2349601|T033|HT|678|ICD9CM|Other fetal conditions|Other fetal conditions
C2349590|T033|HT|678-679.99|ICD9CM|OTHER MATERNAL AND FETAL COMPLICATIONS|OTHER MATERNAL AND FETAL COMPLICATIONS
C2349594|T046|HT|678.0|ICD9CM|Fetal hematologic conditions|Fetal hematologic conditions
C2349591|T046|PT|678.00|ICD9CM|Fetal hematologic conditions, unspecified as to episode of care or not applicable|Fetal hematologic conditions, unspecified as to episode of care or not applicable
C2349591|T046|AB|678.00|ICD9CM|Fetal hematologic-unspec|Fetal hematologic-unspec
C2349592|T046|PT|678.01|ICD9CM|Fetal hematologic conditions, delivered, with or without mention of antepartum condition|Fetal hematologic conditions, delivered, with or without mention of antepartum condition
C2349592|T046|AB|678.01|ICD9CM|Fetal hematologic-deliv|Fetal hematologic-deliv
C2349593|T046|PT|678.03|ICD9CM|Fetal hematologic conditions, antepartum condition or complication|Fetal hematologic conditions, antepartum condition or complication
C2349593|T046|AB|678.03|ICD9CM|Fetal hematologic-ante|Fetal hematologic-ante
C2349600|T046|HT|678.1|ICD9CM|Fetal conjoined twins|Fetal conjoined twins
C2349597|T046|AB|678.10|ICD9CM|Fetal conjoin twins-unsp|Fetal conjoin twins-unsp
C2349597|T046|PT|678.10|ICD9CM|Fetal conjoined twins, unspecified as to episode of care or not applicable|Fetal conjoined twins, unspecified as to episode of care or not applicable
C2349598|T046|AB|678.11|ICD9CM|Fetal conjoin twins-del|Fetal conjoin twins-del
C2349598|T046|PT|678.11|ICD9CM|Fetal conjoined twins, delivered, with or without mention of antepartum condition|Fetal conjoined twins, delivered, with or without mention of antepartum condition
C2349599|T046|AB|678.13|ICD9CM|Fetal conjoin twins-ante|Fetal conjoin twins-ante
C2349599|T046|PT|678.13|ICD9CM|Fetal conjoined twins, antepartum condition or complication|Fetal conjoined twins, antepartum condition or complication
C2349615|T046|HT|679|ICD9CM|Complications of in utero procedures|Complications of in utero procedures
C2349607|T046|HT|679.0|ICD9CM|Maternal complications from in utero procedure|Maternal complications from in utero procedure
C2349602|T046|AB|679.00|ICD9CM|Mat comp in utero-unsp|Mat comp in utero-unsp
C2349602|T046|PT|679.00|ICD9CM|Maternal complications from in utero procedure, unspecified as to episode of care or not applicable|Maternal complications from in utero procedure, unspecified as to episode of care or not applicable
C2349603|T046|AB|679.01|ICD9CM|Mat comp in utero-del|Mat comp in utero-del
C2349604|T046|AB|679.02|ICD9CM|Mat comp in utro-del-p/p|Mat comp in utro-del-p/p
C2349604|T046|PT|679.02|ICD9CM|Maternal complications from in utero procedure, delivered, with mention of postpartum complication|Maternal complications from in utero procedure, delivered, with mention of postpartum complication
C2349605|T046|AB|679.03|ICD9CM|Mat comp in utero-ante|Mat comp in utero-ante
C2349605|T046|PT|679.03|ICD9CM|Maternal complications from in utero procedure, antepartum condition or complication|Maternal complications from in utero procedure, antepartum condition or complication
C2349606|T046|AB|679.04|ICD9CM|Mat comp in utero-p/p|Mat comp in utero-p/p
C2349606|T046|PT|679.04|ICD9CM|Maternal complications from in utero procedure, postpartum condition or complication|Maternal complications from in utero procedure, postpartum condition or complication
C2349613|T046|HT|679.1|ICD9CM|Fetal complications from in utero procedure|Fetal complications from in utero procedure
C2349608|T046|AB|679.10|ICD9CM|Fetal comp in utero-unsp|Fetal comp in utero-unsp
C2349608|T046|PT|679.10|ICD9CM|Fetal complications from in utero procedure, unspecified as to episode of care or not applicable|Fetal complications from in utero procedure, unspecified as to episode of care or not applicable
C2349609|T046|AB|679.11|ICD9CM|Fetal comp in utero-del|Fetal comp in utero-del
C2349610|T046|PT|679.12|ICD9CM|Fetal complications from in utero procedure, delivered, with mention of postpartum complication|Fetal complications from in utero procedure, delivered, with mention of postpartum complication
C2349610|T046|AB|679.12|ICD9CM|Ftl cmp in utro-del-p/p|Ftl cmp in utro-del-p/p
C2349611|T046|AB|679.13|ICD9CM|Fetal comp in utero-ante|Fetal comp in utero-ante
C2349611|T046|PT|679.13|ICD9CM|Fetal complications from in utero procedure, antepartum condition or complication|Fetal complications from in utero procedure, antepartum condition or complication
C2349612|T046|AB|679.14|ICD9CM|Fetal comp in utero-p/p|Fetal comp in utero-p/p
C2349612|T046|PT|679.14|ICD9CM|Fetal complications from in utero procedure, postpartum condition or complication|Fetal complications from in utero procedure, postpartum condition or complication
C0157680|T047|HT|680|ICD9CM|Carbuncle and furuncle|Carbuncle and furuncle
C0037278|T047|HT|680-686.99|ICD9CM|INFECTIONS OF SKIN AND SUBCUTANEOUS TISSUE|INFECTIONS OF SKIN AND SUBCUTANEOUS TISSUE
C0178298|T047|HT|680-709.99|ICD9CM|DISEASES OF THE SKIN AND SUBCUTANEOUS TISSUE|DISEASES OF THE SKIN AND SUBCUTANEOUS TISSUE
C0157681|T047|PT|680.0|ICD9CM|Carbuncle and furuncle of face|Carbuncle and furuncle of face
C0157681|T047|AB|680.0|ICD9CM|Carbuncle of face|Carbuncle of face
C0157682|T047|PT|680.1|ICD9CM|Carbuncle and furuncle of neck|Carbuncle and furuncle of neck
C0157682|T047|AB|680.1|ICD9CM|Carbuncle of neck|Carbuncle of neck
C0157683|T047|PT|680.2|ICD9CM|Carbuncle and furuncle of trunk|Carbuncle and furuncle of trunk
C0157683|T047|AB|680.2|ICD9CM|Carbuncle of trunk|Carbuncle of trunk
C0157684|T047|PT|680.3|ICD9CM|Carbuncle and furuncle of upper arm and forearm|Carbuncle and furuncle of upper arm and forearm
C0157684|T047|AB|680.3|ICD9CM|Carbuncle of arm|Carbuncle of arm
C0157685|T047|PT|680.4|ICD9CM|Carbuncle and furuncle of hand|Carbuncle and furuncle of hand
C0157685|T047|AB|680.4|ICD9CM|Carbuncle of hand|Carbuncle of hand
C0157686|T047|PT|680.5|ICD9CM|Carbuncle and furuncle of buttock|Carbuncle and furuncle of buttock
C0157686|T047|AB|680.5|ICD9CM|Carbuncle of buttock|Carbuncle of buttock
C0157687|T047|PT|680.6|ICD9CM|Carbuncle and furuncle of leg, except foot|Carbuncle and furuncle of leg, except foot
C0157687|T047|AB|680.6|ICD9CM|Carbuncle of leg|Carbuncle of leg
C0157688|T047|PT|680.7|ICD9CM|Carbuncle and furuncle of foot|Carbuncle and furuncle of foot
C0157688|T047|AB|680.7|ICD9CM|Carbuncle of foot|Carbuncle of foot
C0157689|T047|PT|680.8|ICD9CM|Carbuncle and furuncle of other specified sites|Carbuncle and furuncle of other specified sites
C0157689|T047|AB|680.8|ICD9CM|Carbuncle, site NEC|Carbuncle, site NEC
C0007079|T047|PT|680.9|ICD9CM|Carbuncle and furuncle of unspecified site|Carbuncle and furuncle of unspecified site
C0007079|T047|AB|680.9|ICD9CM|Carbuncle NOS|Carbuncle NOS
C0157690|T047|HT|681|ICD9CM|Cellulitis and abscess of finger and toe|Cellulitis and abscess of finger and toe
C0157691|T047|HT|681.0|ICD9CM|Cellulitis and abscess of finger|Cellulitis and abscess of finger
C0157691|T047|PT|681.00|ICD9CM|Cellulitis and abscess of finger, unspecified|Cellulitis and abscess of finger, unspecified
C0157691|T047|AB|681.00|ICD9CM|Cellulitis, finger NOS|Cellulitis, finger NOS
C0152448|T046|AB|681.01|ICD9CM|Felon|Felon
C0152448|T046|PT|681.01|ICD9CM|Felon|Felon
C0157692|T047|PT|681.02|ICD9CM|Onychia and paronychia of finger|Onychia and paronychia of finger
C0157692|T047|AB|681.02|ICD9CM|Onychia of finger|Onychia of finger
C0157693|T047|HT|681.1|ICD9CM|Cellulitis and abscess of toe|Cellulitis and abscess of toe
C0157693|T047|PT|681.10|ICD9CM|Cellulitis and abscess of toe, unspecified|Cellulitis and abscess of toe, unspecified
C0157693|T047|AB|681.10|ICD9CM|Cellulitis, toe NOS|Cellulitis, toe NOS
C0157694|T047|PT|681.11|ICD9CM|Onychia and paronychia of toe|Onychia and paronychia of toe
C0157694|T047|AB|681.11|ICD9CM|Onychia of toe|Onychia of toe
C0007644|T047|PT|681.9|ICD9CM|Cellulitis and abscess of unspecified digit|Cellulitis and abscess of unspecified digit
C0007644|T047|AB|681.9|ICD9CM|Cellulitis of digit NOS|Cellulitis of digit NOS
C0157695|T047|HT|682|ICD9CM|Other cellulitis and abscess|Other cellulitis and abscess
C0157696|T047|PT|682.0|ICD9CM|Cellulitis and abscess of face|Cellulitis and abscess of face
C0157696|T047|AB|682.0|ICD9CM|Cellulitis of face|Cellulitis of face
C0157697|T047|PT|682.1|ICD9CM|Cellulitis and abscess of neck|Cellulitis and abscess of neck
C0157697|T047|AB|682.1|ICD9CM|Cellulitis of neck|Cellulitis of neck
C0157698|T047|PT|682.2|ICD9CM|Cellulitis and abscess of trunk|Cellulitis and abscess of trunk
C0157698|T047|AB|682.2|ICD9CM|Cellulitis of trunk|Cellulitis of trunk
C0157699|T047|PT|682.3|ICD9CM|Cellulitis and abscess of upper arm and forearm|Cellulitis and abscess of upper arm and forearm
C0157699|T047|AB|682.3|ICD9CM|Cellulitis of arm|Cellulitis of arm
C0406078|T047|PT|682.4|ICD9CM|Cellulitis and abscess of hand, except fingers and thumb|Cellulitis and abscess of hand, except fingers and thumb
C0406078|T047|AB|682.4|ICD9CM|Cellulitis of hand|Cellulitis of hand
C0157701|T047|PT|682.5|ICD9CM|Cellulitis and abscess of buttock|Cellulitis and abscess of buttock
C0157701|T047|AB|682.5|ICD9CM|Cellulitis of buttock|Cellulitis of buttock
C0157702|T047|PT|682.6|ICD9CM|Cellulitis and abscess of leg, except foot|Cellulitis and abscess of leg, except foot
C0157702|T047|AB|682.6|ICD9CM|Cellulitis of leg|Cellulitis of leg
C0406089|T047|PT|682.7|ICD9CM|Cellulitis and abscess of foot, except toes|Cellulitis and abscess of foot, except toes
C0406089|T047|AB|682.7|ICD9CM|Cellulitis of foot|Cellulitis of foot
C0157704|T047|PT|682.8|ICD9CM|Cellulitis and abscess of other specified sites|Cellulitis and abscess of other specified sites
C0157704|T047|AB|682.8|ICD9CM|Cellulitis, site NEC|Cellulitis, site NEC
C0007645|T047|PT|682.9|ICD9CM|Cellulitis and abscess of unspecified sites|Cellulitis and abscess of unspecified sites
C0007645|T047|AB|682.9|ICD9CM|Cellulitis NOS|Cellulitis NOS
C0157705|T047|AB|683|ICD9CM|Acute lymphadenitis|Acute lymphadenitis
C0157705|T047|PT|683|ICD9CM|Acute lymphadenitis|Acute lymphadenitis
C0021099|T047|AB|684|ICD9CM|Impetigo|Impetigo
C0021099|T047|PT|684|ICD9CM|Impetigo|Impetigo
C0031925|T047|HT|685|ICD9CM|Pilonidal cyst|Pilonidal cyst
C3537055|T046|AB|685.0|ICD9CM|Pilonidal cyst w abscess|Pilonidal cyst w abscess
C3537055|T046|PT|685.0|ICD9CM|Pilonidal cyst with abscess|Pilonidal cyst with abscess
C0520556|T190|AB|685.1|ICD9CM|Pilonidal cyst w/o absc|Pilonidal cyst w/o absc
C0520556|T190|PT|685.1|ICD9CM|Pilonidal cyst without mention of abscess|Pilonidal cyst without mention of abscess
C0157707|T047|HT|686|ICD9CM|Other local infections of skin and subcutaneous tissue|Other local infections of skin and subcutaneous tissue
C0034212|T047|HT|686.0|ICD9CM|Pyoderma|Pyoderma
C0034212|T047|AB|686.00|ICD9CM|Pyoderma NOS|Pyoderma NOS
C0034212|T047|PT|686.00|ICD9CM|Pyoderma, unspecified|Pyoderma, unspecified
C0085652|T047|AB|686.01|ICD9CM|Pyoderma gangrenosum|Pyoderma gangrenosum
C0085652|T047|PT|686.01|ICD9CM|Pyoderma gangrenosum|Pyoderma gangrenosum
C0490009|T047|PT|686.09|ICD9CM|Other pyoderma|Other pyoderma
C0490009|T047|AB|686.09|ICD9CM|Pyoderma NEC|Pyoderma NEC
C0034214|T046|AB|686.1|ICD9CM|Pyogenic granuloma|Pyogenic granuloma
C0034214|T046|PT|686.1|ICD9CM|Pyogenic granuloma of skin and subcutaneous tissue|Pyogenic granuloma of skin and subcutaneous tissue
C0029813|T046|AB|686.8|ICD9CM|Local skin infection NEC|Local skin infection NEC
C0029813|T046|PT|686.8|ICD9CM|Other specified local infections of skin and subcutaneous tissue|Other specified local infections of skin and subcutaneous tissue
C0406047|T047|AB|686.9|ICD9CM|Local skin infection NOS|Local skin infection NOS
C0406047|T047|PT|686.9|ICD9CM|Unspecified local infection of skin and subcutaneous tissue|Unspecified local infection of skin and subcutaneous tissue
C0014747|T047|HT|690|ICD9CM|Erythematosquamous dermatosis|Erythematosquamous dermatosis
C0178300|T047|HT|690-698.99|ICD9CM|OTHER INFLAMMATORY CONDITIONS OF SKIN AND SUBCUTANEOUS TISSUE|OTHER INFLAMMATORY CONDITIONS OF SKIN AND SUBCUTANEOUS TISSUE
C0036508|T047|HT|690.1|ICD9CM|Seborrheic dermatitis|Seborrheic dermatitis
C0036508|T047|PT|690.10|ICD9CM|Seborrheic dermatitis, unspecified|Seborrheic dermatitis, unspecified
C0036508|T047|AB|690.10|ICD9CM|Sebrrheic dermatitis NOS|Sebrrheic dermatitis NOS
C0221244|T047|AB|690.11|ICD9CM|Seborrhea capitis|Seborrhea capitis
C0221244|T047|PT|690.11|ICD9CM|Seborrhea capitis|Seborrhea capitis
C0343047|T047|AB|690.12|ICD9CM|Sbrheic infantl drmtitis|Sbrheic infantl drmtitis
C0343047|T047|PT|690.12|ICD9CM|Seborrheic infantile dermatitis|Seborrheic infantile dermatitis
C0348768|T047|PT|690.18|ICD9CM|Other seborrheic dermatitis|Other seborrheic dermatitis
C0348768|T047|AB|690.18|ICD9CM|Sebrrheic dermatitis NEC|Sebrrheic dermatitis NEC
C0375481|T047|AB|690.8|ICD9CM|Erythmtsquamous derm NEC|Erythmtsquamous derm NEC
C0375481|T047|PT|690.8|ICD9CM|Other erythematosquamous dermatosis|Other erythematosquamous dermatosis
C0004187|T047|HT|691|ICD9CM|Atopic dermatitis and related conditions|Atopic dermatitis and related conditions
C0011974|T047|AB|691.0|ICD9CM|Diaper or napkin rash|Diaper or napkin rash
C0011974|T047|PT|691.0|ICD9CM|Diaper or napkin rash|Diaper or napkin rash
C0494831|T047|AB|691.8|ICD9CM|Other atopic dermatitis|Other atopic dermatitis
C0494831|T047|PT|691.8|ICD9CM|Other atopic dermatitis and related conditions|Other atopic dermatitis and related conditions
C0009833|T047|HT|692|ICD9CM|Contact dermatitis and other eczema|Contact dermatitis and other eczema
C0157708|T047|PT|692.0|ICD9CM|Contact dermatitis and other eczema due to detergents|Contact dermatitis and other eczema due to detergents
C0157708|T047|AB|692.0|ICD9CM|Detergent dermatitis|Detergent dermatitis
C0157709|T047|PT|692.1|ICD9CM|Contact dermatitis and other eczema due to oils and greases|Contact dermatitis and other eczema due to oils and greases
C0157709|T047|AB|692.1|ICD9CM|Oil & grease dermatitis|Oil & grease dermatitis
C0157710|T047|PT|692.2|ICD9CM|Contact dermatitis and other eczema due to solvents|Contact dermatitis and other eczema due to solvents
C0157710|T047|AB|692.2|ICD9CM|Solvent dermatitis|Solvent dermatitis
C0157711|T047|PT|692.3|ICD9CM|Contact dermatitis and other eczema due to drugs and medicines in contact with skin|Contact dermatitis and other eczema due to drugs and medicines in contact with skin
C0157711|T047|AB|692.3|ICD9CM|Topical med dermatitis|Topical med dermatitis
C0157712|T047|AB|692.4|ICD9CM|Chemical dermatitis NEC|Chemical dermatitis NEC
C0157712|T047|PT|692.4|ICD9CM|Contact dermatitis and other eczema due to other chemical products|Contact dermatitis and other eczema due to other chemical products
C0157713|T047|PT|692.5|ICD9CM|Contact dermatitis and other eczema due to food in contact with skin|Contact dermatitis and other eczema due to food in contact with skin
C0157713|T047|AB|692.5|ICD9CM|Topical food dermatitis|Topical food dermatitis
C0157714|T047|PT|692.6|ICD9CM|Contact dermatitis and other eczema due to plants [except food]|Contact dermatitis and other eczema due to plants [except food]
C0157714|T047|AB|692.6|ICD9CM|Dermatitis due to plant|Dermatitis due to plant
C0157715|T037|HT|692.7|ICD9CM|Contact dermatitis and other eczema due to solar radiation|Contact dermatitis and other eczema due to solar radiation
C0263292|T047|AB|692.70|ICD9CM|Solar dermatitis NOS|Solar dermatitis NOS
C0263292|T047|PT|692.70|ICD9CM|Unspecified dermatitis due to sun|Unspecified dermatitis due to sun
C0038814|T037|AB|692.71|ICD9CM|Sunburn|Sunburn
C0038814|T037|PT|692.71|ICD9CM|Sunburn|Sunburn
C0375482|T047|AB|692.72|ICD9CM|Act drmtitis solar rdiat|Act drmtitis solar rdiat
C0375482|T047|PT|692.72|ICD9CM|Acute dermatitis due to solar radiation|Acute dermatitis due to solar radiation
C0375483|T047|PT|692.73|ICD9CM|Actinic reticuloid and actinic granuloma|Actinic reticuloid and actinic granuloma
C0375483|T047|AB|692.73|ICD9CM|Actnc retic actnc grnlma|Actnc retic actnc grnlma
C0375484|T047|AB|692.74|ICD9CM|Oth chr drmtit solar rad|Oth chr drmtit solar rad
C0375484|T047|PT|692.74|ICD9CM|Other chronic dermatitis due to solar radiation|Other chronic dermatitis due to solar radiation
C0265970|T047|AB|692.75|ICD9CM|Dis sup actnc porokrtsis|Dis sup actnc porokrtsis
C0265970|T047|PT|692.75|ICD9CM|Disseminated superficial actinic porokeratosis (DSAP)|Disseminated superficial actinic porokeratosis (DSAP)
C0451998|T037|AB|692.76|ICD9CM|2nd degree sunburn|2nd degree sunburn
C0451998|T037|PT|692.76|ICD9CM|Sunburn of second degree|Sunburn of second degree
C0452001|T037|AB|692.77|ICD9CM|3rd degree sunburn|3rd degree sunburn
C0452001|T037|PT|692.77|ICD9CM|Sunburn of third degree|Sunburn of third degree
C0375485|T047|AB|692.79|ICD9CM|Oth dermatitis solar rad|Oth dermatitis solar rad
C0375485|T047|PT|692.79|ICD9CM|Other dermatitis due to solar radiation|Other dermatitis due to solar radiation
C0009834|T047|HT|692.8|ICD9CM|Contact dermatitis and other eczema due to other specified agents|Contact dermatitis and other eczema due to other specified agents
C0263296|T047|AB|692.81|ICD9CM|Cosmetic dermatitis|Cosmetic dermatitis
C0263296|T047|PT|692.81|ICD9CM|Dermatitis due to cosmetics|Dermatitis due to cosmetics
C0375486|T047|PT|692.82|ICD9CM|Dermatitis due to other radiation|Dermatitis due to other radiation
C0375486|T047|AB|692.82|ICD9CM|Dermatitis oth radiation|Dermatitis oth radiation
C0263304|T047|PT|692.83|ICD9CM|Dermatitis due to metals|Dermatitis due to metals
C0263304|T047|AB|692.83|ICD9CM|Dermatitis metals|Dermatitis metals
C1456114|T047|PT|692.84|ICD9CM|Contact dermatitis and other eczema due to animal (cat) (dog) dander|Contact dermatitis and other eczema due to animal (cat) (dog) dander
C1456114|T047|AB|692.84|ICD9CM|Contact drmatitis-animal|Contact drmatitis-animal
C0009834|T047|PT|692.89|ICD9CM|Contact dermatitis and other eczema due to other specified agents|Contact dermatitis and other eczema due to other specified agents
C0009834|T047|AB|692.89|ICD9CM|Dermatitis NEC|Dermatitis NEC
C0375487|T047|PT|692.9|ICD9CM|Contact dermatitis and other eczema, unspecified cause|Contact dermatitis and other eczema, unspecified cause
C0375487|T047|AB|692.9|ICD9CM|Dermatitis NOS|Dermatitis NOS
C0157718|T047|HT|693|ICD9CM|Dermatitis due to substances taken internally|Dermatitis due to substances taken internally
C0011604|T046|PT|693.0|ICD9CM|Dermatitis due to drugs and medicines taken internally|Dermatitis due to drugs and medicines taken internally
C0011604|T046|AB|693.0|ICD9CM|Drug dermatitis NOS|Drug dermatitis NOS
C0494843|T047|AB|693.1|ICD9CM|Dermat d/t food ingest|Dermat d/t food ingest
C0494843|T047|PT|693.1|ICD9CM|Dermatitis due to food taken internally|Dermatitis due to food taken internally
C0157719|T046|AB|693.8|ICD9CM|Dermat d/t int agent NEC|Dermat d/t int agent NEC
C0157719|T046|PT|693.8|ICD9CM|Dermatitis due to other specified substances taken internally|Dermatitis due to other specified substances taken internally
C0157718|T047|AB|693.9|ICD9CM|Dermat d/t int agent NOS|Dermat d/t int agent NOS
C0157718|T047|PT|693.9|ICD9CM|Dermatitis due to unspecified substance taken internally|Dermatitis due to unspecified substance taken internally
C0085932|T047|HT|694|ICD9CM|Bullous dermatoses|Bullous dermatoses
C0011608|T047|AB|694.0|ICD9CM|Dermatitis herpetiformis|Dermatitis herpetiformis
C0011608|T047|PT|694.0|ICD9CM|Dermatitis herpetiformis|Dermatitis herpetiformis
C0600336|T047|AB|694.1|ICD9CM|Subcorneal pust dermatos|Subcorneal pust dermatos
C0600336|T047|PT|694.1|ICD9CM|Subcorneal pustular dermatosis|Subcorneal pustular dermatosis
C0152092|T047|AB|694.2|ICD9CM|Juven dermat herpetiform|Juven dermat herpetiform
C0152092|T047|PT|694.2|ICD9CM|Juvenile dermatitis herpetiformis|Juvenile dermatitis herpetiformis
C1314968|T047|AB|694.3|ICD9CM|Impetigo herpetiformis|Impetigo herpetiformis
C1314968|T047|PT|694.3|ICD9CM|Impetigo herpetiformis|Impetigo herpetiformis
C0030807|T047|AB|694.4|ICD9CM|Pemphigus|Pemphigus
C0030807|T047|PT|694.4|ICD9CM|Pemphigus|Pemphigus
C0030805|T047|AB|694.5|ICD9CM|Pemphigoid|Pemphigoid
C0030805|T047|PT|694.5|ICD9CM|Pemphigoid|Pemphigoid
C0030804|T047|HT|694.6|ICD9CM|Benign mucous membrane pemphigoid|Benign mucous membrane pemphigoid
C1367974|T047|PT|694.60|ICD9CM|Benign mucous membrane pemphigoid without mention of ocular involvement|Benign mucous membrane pemphigoid without mention of ocular involvement
C1367974|T047|AB|694.60|ICD9CM|Bn mucous memb pemph NOS|Bn mucous memb pemph NOS
C0157721|T047|PT|694.61|ICD9CM|Benign mucous membrane pemphigoid with ocular involvement|Benign mucous membrane pemphigoid with ocular involvement
C0157721|T047|AB|694.61|ICD9CM|Ocular pemphigus|Ocular pemphigus
C0079957|T047|AB|694.8|ICD9CM|Bullous dermatoses NEC|Bullous dermatoses NEC
C0079957|T047|PT|694.8|ICD9CM|Other specified bullous dermatoses|Other specified bullous dermatoses
C0085932|T047|AB|694.9|ICD9CM|Bullous dermatoses NOS|Bullous dermatoses NOS
C0085932|T047|PT|694.9|ICD9CM|Unspecified bullous dermatoses|Unspecified bullous dermatoses
C0041834|T047|HT|695|ICD9CM|Erythematous conditions|Erythematous conditions
C0152251|T047|AB|695.0|ICD9CM|Toxic erythema|Toxic erythema
C0152251|T047|PT|695.0|ICD9CM|Toxic erythema|Toxic erythema
C0014742|T047|HT|695.1|ICD9CM|Erythema multiforme|Erythema multiforme
C0014742|T047|AB|695.10|ICD9CM|Erythema multiforme NOS|Erythema multiforme NOS
C0014742|T047|PT|695.10|ICD9CM|Erythema multiforme, unspecified|Erythema multiforme, unspecified
C0857751|T047|PT|695.11|ICD9CM|Erythema multiforme minor|Erythema multiforme minor
C0857751|T047|AB|695.11|ICD9CM|Erythma multiforme minor|Erythma multiforme minor
C3241919|T047|AB|695.12|ICD9CM|Erythema multiforme maj|Erythema multiforme maj
C3241919|T047|PT|695.12|ICD9CM|Erythema multiforme major|Erythema multiforme major
C0038325|T047|PT|695.13|ICD9CM|Stevens-Johnson syndrome|Stevens-Johnson syndrome
C0038325|T047|AB|695.13|ICD9CM|Stevens-Johnson syndrome|Stevens-Johnson syndrome
C2349616|T047|PT|695.14|ICD9CM|Stevens-Johnson syndrome-toxic epidermal necrolysis overlap syndrome|Stevens-Johnson syndrome-toxic epidermal necrolysis overlap syndrome
C2349616|T047|AB|695.14|ICD9CM|Stevens-Johnson-TEN syn|Stevens-Johnson-TEN syn
C0014518|T047|PT|695.15|ICD9CM|Toxic epidermal necrolysis|Toxic epidermal necrolysis
C0014518|T047|AB|695.15|ICD9CM|Toxic epidrml necrolysis|Toxic epidrml necrolysis
C0477492|T047|AB|695.19|ICD9CM|Erythema multiforme NEC|Erythema multiforme NEC
C0477492|T047|PT|695.19|ICD9CM|Other erythema multiforme|Other erythema multiforme
C0014743|T047|AB|695.2|ICD9CM|Erythema nodosum|Erythema nodosum
C0014743|T047|PT|695.2|ICD9CM|Erythema nodosum|Erythema nodosum
C0035854|T047|AB|695.3|ICD9CM|Rosacea|Rosacea
C0035854|T047|PT|695.3|ICD9CM|Rosacea|Rosacea
C0409974|T047|AB|695.4|ICD9CM|Lupus erythematosus|Lupus erythematosus
C0409974|T047|PT|695.4|ICD9CM|Lupus erythematosus|Lupus erythematosus
C2349629|T047|HT|695.5|ICD9CM|Exfoliation due to erythematous conditions according to extent of body surface involved|Exfoliation due to erythematous conditions according to extent of body surface involved
C2349618|T047|AB|695.50|ICD9CM|Exfol d/t eryth <10% bdy|Exfol d/t eryth <10% bdy
C2349618|T047|PT|695.50|ICD9CM|Exfoliation due to erythematous condition involving less than 10 percent of body surface|Exfoliation due to erythematous condition involving less than 10 percent of body surface
C2349620|T047|AB|695.51|ICD9CM|Exfl d/t eryth 10-19 bdy|Exfl d/t eryth 10-19 bdy
C2349620|T047|PT|695.51|ICD9CM|Exfoliation due to erythematous condition involving 10-19 percent of body surface|Exfoliation due to erythematous condition involving 10-19 percent of body surface
C2349621|T047|AB|695.52|ICD9CM|Exfl d/t eryth 20-29 bdy|Exfl d/t eryth 20-29 bdy
C2349621|T047|PT|695.52|ICD9CM|Exfoliation due to erythematous condition involving 20-29 percent of body surface|Exfoliation due to erythematous condition involving 20-29 percent of body surface
C2349622|T047|AB|695.53|ICD9CM|Exfl d/t eryth 30-39 bdy|Exfl d/t eryth 30-39 bdy
C2349622|T047|PT|695.53|ICD9CM|Exfoliation due to erythematous condition involving 30-39 percent of body surface|Exfoliation due to erythematous condition involving 30-39 percent of body surface
C2349623|T047|AB|695.54|ICD9CM|Exfl d/t eryth 40-49 bdy|Exfl d/t eryth 40-49 bdy
C2349623|T047|PT|695.54|ICD9CM|Exfoliation due to erythematous condition involving 40-49 percent of body surface|Exfoliation due to erythematous condition involving 40-49 percent of body surface
C2349624|T047|AB|695.55|ICD9CM|Exfl d/t eryth 50-59 bdy|Exfl d/t eryth 50-59 bdy
C2349624|T047|PT|695.55|ICD9CM|Exfoliation due to erythematous condition involving 50-59 percent of body surface|Exfoliation due to erythematous condition involving 50-59 percent of body surface
C2349625|T047|AB|695.56|ICD9CM|Exfl d/t eryth 60-69 bdy|Exfl d/t eryth 60-69 bdy
C2349625|T047|PT|695.56|ICD9CM|Exfoliation due to erythematous condition involving 60-69 percent of body surface|Exfoliation due to erythematous condition involving 60-69 percent of body surface
C2349626|T047|AB|695.57|ICD9CM|Exfl d/t eryth 70-79 bdy|Exfl d/t eryth 70-79 bdy
C2349626|T047|PT|695.57|ICD9CM|Exfoliation due to erythematous condition involving 70-79 percent of body surface|Exfoliation due to erythematous condition involving 70-79 percent of body surface
C2349627|T047|AB|695.58|ICD9CM|Exfl d/t eryth 80-89 bdy|Exfl d/t eryth 80-89 bdy
C2349627|T047|PT|695.58|ICD9CM|Exfoliation due to erythematous condition involving 80-89 percent of body surface|Exfoliation due to erythematous condition involving 80-89 percent of body surface
C2349628|T047|AB|695.59|ICD9CM|Exfl d/t eryth >=90% bdy|Exfl d/t eryth >=90% bdy
C2349628|T047|PT|695.59|ICD9CM|Exfoliation due to erythematous condition involving 90 percent or more of body surface|Exfoliation due to erythematous condition involving 90 percent or more of body surface
C0029794|T047|HT|695.8|ICD9CM|Other specified erythematous conditions|Other specified erythematous conditions
C0038165|T047|AB|695.81|ICD9CM|Ritter's disease|Ritter's disease
C0038165|T047|PT|695.81|ICD9CM|Ritter's disease|Ritter's disease
C0029794|T047|AB|695.89|ICD9CM|Erythematous cond NEC|Erythematous cond NEC
C0029794|T047|PT|695.89|ICD9CM|Other specified erythematous conditions|Other specified erythematous conditions
C0041834|T047|AB|695.9|ICD9CM|Erythematous cond NOS|Erythematous cond NOS
C0041834|T047|PT|695.9|ICD9CM|Unspecified erythematous condition|Unspecified erythematous condition
C0157723|T047|HT|696|ICD9CM|Psoriasis and similar disorders|Psoriasis and similar disorders
C0003872|T047|AB|696.0|ICD9CM|Psoriatic arthropathy|Psoriatic arthropathy
C0003872|T047|PT|696.0|ICD9CM|Psoriatic arthropathy|Psoriatic arthropathy
C0490052|T047|AB|696.1|ICD9CM|Other psoriasis|Other psoriasis
C0490052|T047|PT|696.1|ICD9CM|Other psoriasis|Other psoriasis
C0030491|T047|AB|696.2|ICD9CM|Parapsoriasis|Parapsoriasis
C0030491|T047|PT|696.2|ICD9CM|Parapsoriasis|Parapsoriasis
C0032026|T047|AB|696.3|ICD9CM|Pityriasis rosea|Pityriasis rosea
C0032026|T047|PT|696.3|ICD9CM|Pityriasis rosea|Pityriasis rosea
C0032027|T047|AB|696.4|ICD9CM|Pityriasis rubra pilaris|Pityriasis rubra pilaris
C0032027|T047|PT|696.4|ICD9CM|Pityriasis rubra pilaris|Pityriasis rubra pilaris
C0029514|T047|PT|696.5|ICD9CM|Other and unspecified pityriasis|Other and unspecified pityriasis
C0029514|T047|AB|696.5|ICD9CM|Pityriasis NEC & NOS|Pityriasis NEC & NOS
C0029717|T047|PT|696.8|ICD9CM|Other psoriasis and similar disorders|Other psoriasis and similar disorders
C0029717|T047|AB|696.8|ICD9CM|Psorias related dis NEC|Psorias related dis NEC
C0023643|T047|HT|697|ICD9CM|Lichen|Lichen
C0023646|T047|AB|697.0|ICD9CM|Lichen planus|Lichen planus
C0023646|T047|PT|697.0|ICD9CM|Lichen planus|Lichen planus
C0162849|T047|AB|697.1|ICD9CM|Lichen nitidus|Lichen nitidus
C0162849|T047|PT|697.1|ICD9CM|Lichen nitidus|Lichen nitidus
C0868870|T047|AB|697.8|ICD9CM|Lichen NEC|Lichen NEC
C0868870|T047|PT|697.8|ICD9CM|Other lichen, not elsewhere classified|Other lichen, not elsewhere classified
C0023643|T047|AB|697.9|ICD9CM|Lichen NOS|Lichen NOS
C0023643|T047|PT|697.9|ICD9CM|Lichen, unspecified|Lichen, unspecified
C0157724|T184|HT|698|ICD9CM|Pruritus and related conditions|Pruritus and related conditions
C0033775|T184|AB|698.0|ICD9CM|Pruritus ani|Pruritus ani
C0033775|T184|PT|698.0|ICD9CM|Pruritus ani|Pruritus ani
C0033777|T184|PT|698.1|ICD9CM|Pruritus of genital organs|Pruritus of genital organs
C0033777|T184|AB|698.1|ICD9CM|Pruritus of genitalia|Pruritus of genitalia
C0033771|T047|AB|698.2|ICD9CM|Prurigo|Prurigo
C0033771|T047|PT|698.2|ICD9CM|Prurigo|Prurigo
C0023654|T047|AB|698.3|ICD9CM|Lichenification|Lichenification
C0023654|T047|PT|698.3|ICD9CM|Lichenification and lichen simplex chronicus|Lichenification and lichen simplex chronicus
C1274184|T047|AB|698.4|ICD9CM|Dermatitis factitia|Dermatitis factitia
C1274184|T047|PT|698.4|ICD9CM|Dermatitis factitia [artefacta]|Dermatitis factitia [artefacta]
C0157725|T184|PT|698.8|ICD9CM|Other specified pruritic conditions|Other specified pruritic conditions
C0157725|T184|AB|698.8|ICD9CM|Pruritic conditions NEC|Pruritic conditions NEC
C0033774|T033|AB|698.9|ICD9CM|Pruritic disorder NOS|Pruritic disorder NOS
C0033774|T033|PT|698.9|ICD9CM|Unspecified pruritic disorder|Unspecified pruritic disorder
C0157726|T020|AB|700|ICD9CM|Corns and callosities|Corns and callosities
C0157726|T020|PT|700|ICD9CM|Corns and callosities|Corns and callosities
C0178301|T047|HT|700-709.99|ICD9CM|OTHER DISEASES OF SKIN AND SUBCUTANEOUS TISSUE|OTHER DISEASES OF SKIN AND SUBCUTANEOUS TISSUE
C0157727|T046|HT|701|ICD9CM|Other hypertrophic and atrophic conditions of skin|Other hypertrophic and atrophic conditions of skin
C0036420|T047|AB|701.0|ICD9CM|Circumscribe scleroderma|Circumscribe scleroderma
C0036420|T047|PT|701.0|ICD9CM|Circumscribed scleroderma|Circumscribed scleroderma
C0022581|T020|AB|701.1|ICD9CM|Keratoderma, acquired|Keratoderma, acquired
C0022581|T020|PT|701.1|ICD9CM|Keratoderma, acquired|Keratoderma, acquired
C0392440|T020|AB|701.2|ICD9CM|Acq acanthosis nigricans|Acq acanthosis nigricans
C0392440|T020|PT|701.2|ICD9CM|Acquired acanthosis nigricans|Acquired acanthosis nigricans
C0152459|T020|AB|701.3|ICD9CM|Striae atrophicae|Striae atrophicae
C0152459|T020|PT|701.3|ICD9CM|Striae atrophicae|Striae atrophicae
C0022548|T020|AB|701.4|ICD9CM|Keloid scar|Keloid scar
C0022548|T020|PT|701.4|ICD9CM|Keloid scar|Keloid scar
C0157729|T047|AB|701.5|ICD9CM|Abnormal granulation NEC|Abnormal granulation NEC
C0157729|T047|PT|701.5|ICD9CM|Other abnormal granulation tissue|Other abnormal granulation tissue
C0029805|T047|PT|701.8|ICD9CM|Other specified hypertrophic and atrophic conditions of skin|Other specified hypertrophic and atrophic conditions of skin
C0029805|T047|AB|701.8|ICD9CM|Skin hypertro/atroph NEC|Skin hypertro/atroph NEC
C0041847|T047|AB|701.9|ICD9CM|Skin hypertro/atroph NOS|Skin hypertro/atroph NOS
C0041847|T047|PT|701.9|ICD9CM|Unspecified hypertrophic and atrophic conditions of skin|Unspecified hypertrophic and atrophic conditions of skin
C0029574|T047|HT|702|ICD9CM|Other dermatoses|Other dermatoses
C0022602|T191|AB|702.0|ICD9CM|Actinic keratosis|Actinic keratosis
C0022602|T191|PT|702.0|ICD9CM|Actinic keratosis|Actinic keratosis
C0022603|T191|HT|702.1|ICD9CM|Seborrheic keratosis|Seborrheic keratosis
C0376117|T191|AB|702.11|ICD9CM|Inflamed sbrheic keratos|Inflamed sbrheic keratos
C0376117|T191|PT|702.11|ICD9CM|Inflamed seborrheic keratosis|Inflamed seborrheic keratosis
C0375488|T047|AB|702.19|ICD9CM|Other sborheic keratosis|Other sborheic keratosis
C0375488|T047|PT|702.19|ICD9CM|Other seborrheic keratosis|Other seborrheic keratosis
C0157730|T047|AB|702.8|ICD9CM|Other specf dermatoses|Other specf dermatoses
C0157730|T047|PT|702.8|ICD9CM|Other specified dermatoses|Other specified dermatoses
C0027339|T047|HT|703|ICD9CM|Diseases of nail|Diseases of nail
C0027343|T033|AB|703.0|ICD9CM|Ingrowing nail|Ingrowing nail
C0027343|T033|PT|703.0|ICD9CM|Ingrowing nail|Ingrowing nail
C0157731|T047|AB|703.8|ICD9CM|Diseases of nail NEC|Diseases of nail NEC
C0157731|T047|PT|703.8|ICD9CM|Other specified diseases of nail|Other specified diseases of nail
C0027339|T047|AB|703.9|ICD9CM|Disease of nail NOS|Disease of nail NOS
C0027339|T047|PT|703.9|ICD9CM|Unspecified disease of nail|Unspecified disease of nail
C0554472|T047|HT|704|ICD9CM|Diseases of hair and hair follicles|Diseases of hair and hair follicles
C0002170|T047|HT|704.0|ICD9CM|Alopecia|Alopecia
C0002170|T047|AB|704.00|ICD9CM|Alopecia NOS|Alopecia NOS
C0002170|T047|PT|704.00|ICD9CM|Alopecia, unspecified|Alopecia, unspecified
C0002171|T047|AB|704.01|ICD9CM|Alopecia areata|Alopecia areata
C0002171|T047|PT|704.01|ICD9CM|Alopecia areata|Alopecia areata
C0263518|T047|AB|704.02|ICD9CM|Telogen effluvium|Telogen effluvium
C0263518|T047|PT|704.02|ICD9CM|Telogen effluvium|Telogen effluvium
C0029489|T047|AB|704.09|ICD9CM|Alopecia NEC|Alopecia NEC
C0029489|T047|PT|704.09|ICD9CM|Other alopecia|Other alopecia
C0019572|T033|AB|704.1|ICD9CM|Hirsutism|Hirsutism
C0019572|T033|PT|704.1|ICD9CM|Hirsutism|Hirsutism
C0157733|T033|AB|704.2|ICD9CM|Abnormalities of hair|Abnormalities of hair
C0157733|T033|PT|704.2|ICD9CM|Abnormalities of the hair|Abnormalities of the hair
C0157734|T033|AB|704.3|ICD9CM|Variations in hair color|Variations in hair color
C0157734|T033|PT|704.3|ICD9CM|Variations in hair color|Variations in hair color
C3161259|T047|HT|704.4|ICD9CM|Pilar and trichilemmal cysts|Pilar and trichilemmal cysts
C0086809|T190|PT|704.41|ICD9CM|Pilar cyst|Pilar cyst
C0086809|T190|AB|704.41|ICD9CM|Pilar cyst|Pilar cyst
C2266788|T047|AB|704.42|ICD9CM|Trichilemmal cyst|Trichilemmal cyst
C2266788|T047|PT|704.42|ICD9CM|Trichilemmal cyst|Trichilemmal cyst
C0029769|T047|AB|704.8|ICD9CM|Hair diseases NEC|Hair diseases NEC
C0029769|T047|PT|704.8|ICD9CM|Other specified diseases of hair and hair follicles|Other specified diseases of hair and hair follicles
C0554472|T047|AB|704.9|ICD9CM|Hair disease NOS|Hair disease NOS
C0554472|T047|PT|704.9|ICD9CM|Unspecified disease of hair and hair follicles|Unspecified disease of hair and hair follicles
C0038986|T047|HT|705|ICD9CM|Disorders of sweat glands|Disorders of sweat glands
C0003028|T047|AB|705.0|ICD9CM|Anhidrosis|Anhidrosis
C0003028|T047|PT|705.0|ICD9CM|Anhidrosis|Anhidrosis
C0162423|T047|AB|705.1|ICD9CM|Prickly heat|Prickly heat
C0162423|T047|PT|705.1|ICD9CM|Prickly heat|Prickly heat
C0476475|T033|HT|705.2|ICD9CM|Focal hyperhidrosis|Focal hyperhidrosis
C1456132|T047|PT|705.21|ICD9CM|Primary focal hyperhidrosis|Primary focal hyperhidrosis
C1456132|T047|AB|705.21|ICD9CM|Primary focal hyprhidros|Primary focal hyprhidros
C1456136|T047|AB|705.22|ICD9CM|Sec focal hyperhidrosis|Sec focal hyperhidrosis
C1456136|T047|PT|705.22|ICD9CM|Secondary focal hyperhidrosis|Secondary focal hyperhidrosis
C0157735|T047|HT|705.8|ICD9CM|Other specified disorders of sweat glands|Other specified disorders of sweat glands
C0032633|T047|AB|705.81|ICD9CM|Dyshidrosis|Dyshidrosis
C0032633|T047|PT|705.81|ICD9CM|Dyshidrosis|Dyshidrosis
C0016632|T047|AB|705.82|ICD9CM|Fox-fordyce disease|Fox-fordyce disease
C0016632|T047|PT|705.82|ICD9CM|Fox-Fordyce disease|Fox-Fordyce disease
C0085160|T047|AB|705.83|ICD9CM|Hidradenitis|Hidradenitis
C0085160|T047|PT|705.83|ICD9CM|Hidradenitis|Hidradenitis
C0157735|T047|PT|705.89|ICD9CM|Other specified disorders of sweat glands|Other specified disorders of sweat glands
C0157735|T047|AB|705.89|ICD9CM|Sweat gland disorder NEC|Sweat gland disorder NEC
C0038986|T047|AB|705.9|ICD9CM|Sweat gland disorder NOS|Sweat gland disorder NOS
C0038986|T047|PT|705.9|ICD9CM|Unspecified disorder of sweat glands|Unspecified disorder of sweat glands
C0036502|T047|HT|706|ICD9CM|Diseases of sebaceous glands|Diseases of sebaceous glands
C0152249|T047|AB|706.0|ICD9CM|Acne varioliformis|Acne varioliformis
C0152249|T047|PT|706.0|ICD9CM|Acne varioliformis|Acne varioliformis
C0029485|T047|AB|706.1|ICD9CM|Acne NEC|Acne NEC
C0029485|T047|PT|706.1|ICD9CM|Other acne|Other acne
C0014511|T190|AB|706.2|ICD9CM|Sebaceous cyst|Sebaceous cyst
C0014511|T190|PT|706.2|ICD9CM|Sebaceous cyst|Sebaceous cyst
C0036508|T047|AB|706.3|ICD9CM|Seborrhea|Seborrhea
C0036508|T047|PT|706.3|ICD9CM|Seborrhea|Seborrhea
C0157736|T047|PT|706.8|ICD9CM|Other specified diseases of sebaceous glands|Other specified diseases of sebaceous glands
C0157736|T047|AB|706.8|ICD9CM|Sebaceous gland dis NEC|Sebaceous gland dis NEC
C0036502|T047|AB|706.9|ICD9CM|Sebaceous gland dis NOS|Sebaceous gland dis NOS
C0036502|T047|PT|706.9|ICD9CM|Unspecified disease of sebaceous glands|Unspecified disease of sebaceous glands
C0157738|T047|HT|707|ICD9CM|Chronic ulcer of skin|Chronic ulcer of skin
C0011127|T047|HT|707.0|ICD9CM|Pressure ulcer|Pressure ulcer
C0011127|T047|AB|707.00|ICD9CM|Pressure ulcer, site NOS|Pressure ulcer, site NOS
C0011127|T047|PT|707.00|ICD9CM|Pressure ulcer, unspecified site|Pressure ulcer, unspecified site
C0558156|T047|AB|707.01|ICD9CM|Pressure ulcer, elbow|Pressure ulcer, elbow
C0558156|T047|PT|707.01|ICD9CM|Pressure ulcer, elbow|Pressure ulcer, elbow
C1456139|T046|PT|707.02|ICD9CM|Pressure ulcer, upper back|Pressure ulcer, upper back
C1456139|T046|AB|707.02|ICD9CM|Pressure ulcer, upr back|Pressure ulcer, upr back
C1456141|T047|AB|707.03|ICD9CM|Pressure ulcer, low back|Pressure ulcer, low back
C1456141|T047|PT|707.03|ICD9CM|Pressure ulcer, lower back|Pressure ulcer, lower back
C0577712|T046|AB|707.04|ICD9CM|Pressure ulcer, hip|Pressure ulcer, hip
C0577712|T046|PT|707.04|ICD9CM|Pressure ulcer, hip|Pressure ulcer, hip
C0558160|T047|AB|707.05|ICD9CM|Pressure ulcer, buttock|Pressure ulcer, buttock
C0558160|T047|PT|707.05|ICD9CM|Pressure ulcer, buttock|Pressure ulcer, buttock
C0577713|T047|AB|707.06|ICD9CM|Pressure ulcer, ankle|Pressure ulcer, ankle
C0577713|T047|PT|707.06|ICD9CM|Pressure ulcer, ankle|Pressure ulcer, ankle
C0558158|T047|AB|707.07|ICD9CM|Pressure ulcer, heel|Pressure ulcer, heel
C0558158|T047|PT|707.07|ICD9CM|Pressure ulcer, heel|Pressure ulcer, heel
C1456142|T047|PT|707.09|ICD9CM|Pressure ulcer, other site|Pressure ulcer, other site
C1456142|T047|AB|707.09|ICD9CM|Pressure ulcer, site NEC|Pressure ulcer, site NEC
C2349630|T047|HT|707.1|ICD9CM|Ulcer of lower limbs, except pressure ulcer|Ulcer of lower limbs, except pressure ulcer
C0878700|T047|AB|707.10|ICD9CM|Ulcer of lower limb NOS|Ulcer of lower limb NOS
C0878700|T047|PT|707.10|ICD9CM|Ulcer of lower limb, unspecified|Ulcer of lower limb, unspecified
C0878701|T047|AB|707.11|ICD9CM|Ulcer of thigh|Ulcer of thigh
C0878701|T047|PT|707.11|ICD9CM|Ulcer of thigh|Ulcer of thigh
C0577719|T047|AB|707.12|ICD9CM|Ulcer of calf|Ulcer of calf
C0577719|T047|PT|707.12|ICD9CM|Ulcer of calf|Ulcer of calf
C0741085|T047|AB|707.13|ICD9CM|Ulcer of ankle|Ulcer of ankle
C0741085|T047|PT|707.13|ICD9CM|Ulcer of ankle|Ulcer of ankle
C0878702|T047|AB|707.14|ICD9CM|Ulcer of heel & midfoot|Ulcer of heel & midfoot
C0878702|T047|PT|707.14|ICD9CM|Ulcer of heel and midfoot|Ulcer of heel and midfoot
C0878703|T047|PT|707.15|ICD9CM|Ulcer of other part of foot|Ulcer of other part of foot
C0878703|T047|AB|707.15|ICD9CM|Ulcer other part of foot|Ulcer other part of foot
C0878704|T047|PT|707.19|ICD9CM|Ulcer of other part of lower limb|Ulcer of other part of lower limb
C0878704|T047|AB|707.19|ICD9CM|Ulcer oth part low limb|Ulcer oth part low limb
C1718233|T033|HT|707.2|ICD9CM|Pressure ulcer stages|Pressure ulcer stages
C2349631|T047|PT|707.20|ICD9CM|Pressure ulcer, unspecified stage|Pressure ulcer, unspecified stage
C2349631|T047|AB|707.20|ICD9CM|Pressure ulcer,stage NOS|Pressure ulcer,stage NOS
C1720599|T047|AB|707.21|ICD9CM|Pressure ulcer, stage I|Pressure ulcer, stage I
C1720599|T047|PT|707.21|ICD9CM|Pressure ulcer, stage I|Pressure ulcer, stage I
C1720518|T047|AB|707.22|ICD9CM|Pressure ulcer, stage II|Pressure ulcer, stage II
C1720518|T047|PT|707.22|ICD9CM|Pressure ulcer, stage II|Pressure ulcer, stage II
C1719811|T047|PT|707.23|ICD9CM|Pressure ulcer, stage III|Pressure ulcer, stage III
C1719811|T047|AB|707.23|ICD9CM|Pressure ulcer,stage III|Pressure ulcer,stage III
C1719910|T047|AB|707.24|ICD9CM|Pressure ulcer, stage IV|Pressure ulcer, stage IV
C1719910|T047|PT|707.24|ICD9CM|Pressure ulcer, stage IV|Pressure ulcer, stage IV
C2368027|T047|PT|707.25|ICD9CM|Pressure ulcer, unstageable|Pressure ulcer, unstageable
C2368027|T047|AB|707.25|ICD9CM|Pressure ulcer,unstagebl|Pressure ulcer,unstagebl
C0157740|T047|AB|707.8|ICD9CM|Chronic skin ulcer NEC|Chronic skin ulcer NEC
C0157740|T047|PT|707.8|ICD9CM|Chronic ulcer of other specified sites|Chronic ulcer of other specified sites
C0333297|T047|AB|707.9|ICD9CM|Chronic skin ulcer NOS|Chronic skin ulcer NOS
C0333297|T047|PT|707.9|ICD9CM|Chronic ulcer of unspecified site|Chronic ulcer of unspecified site
C0042109|T047|HT|708|ICD9CM|Urticaria|Urticaria
C0149526|T047|AB|708.0|ICD9CM|Allergic urticaria|Allergic urticaria
C0149526|T047|PT|708.0|ICD9CM|Allergic urticaria|Allergic urticaria
C0157741|T047|AB|708.1|ICD9CM|Idiopathic urticaria|Idiopathic urticaria
C0157741|T047|PT|708.1|ICD9CM|Idiopathic urticaria|Idiopathic urticaria
C0157742|T037|PT|708.2|ICD9CM|Urticaria due to cold and heat|Urticaria due to cold and heat
C0157742|T037|AB|708.2|ICD9CM|Urticaria from cold/heat|Urticaria from cold/heat
C0343065|T047|AB|708.3|ICD9CM|Dermatographic urticaria|Dermatographic urticaria
C0343065|T047|PT|708.3|ICD9CM|Dermatographic urticaria|Dermatographic urticaria
C0157743|T047|AB|708.4|ICD9CM|Vibratory urticaria|Vibratory urticaria
C0157743|T047|PT|708.4|ICD9CM|Vibratory urticaria|Vibratory urticaria
C0152230|T047|AB|708.5|ICD9CM|Cholinergic urticaria|Cholinergic urticaria
C0152230|T047|PT|708.5|ICD9CM|Cholinergic urticaria|Cholinergic urticaria
C0029839|T047|PT|708.8|ICD9CM|Other specified urticaria|Other specified urticaria
C0029839|T047|AB|708.8|ICD9CM|Urticaria NEC|Urticaria NEC
C0042109|T047|AB|708.9|ICD9CM|Urticaria NOS|Urticaria NOS
C0042109|T047|PT|708.9|ICD9CM|Urticaria, unspecified|Urticaria, unspecified
C0178301|T047|HT|709|ICD9CM|Other disorders of skin and subcutaneous tissue|Other disorders of skin and subcutaneous tissue
C0151907|T033|HT|709.0|ICD9CM|Dyschromia|Dyschromia
C0151907|T033|AB|709.00|ICD9CM|Dyschromia, unspecified|Dyschromia, unspecified
C0151907|T033|PT|709.00|ICD9CM|Dyschromia, unspecified|Dyschromia, unspecified
C0042900|T047|AB|709.01|ICD9CM|Vitiligo|Vitiligo
C0042900|T047|PT|709.01|ICD9CM|Vitiligo|Vitiligo
C0375489|T047|AB|709.09|ICD9CM|Other dyschromia|Other dyschromia
C0375489|T047|PT|709.09|ICD9CM|Other dyschromia|Other dyschromia
C0162819|T047|AB|709.1|ICD9CM|Vascular disord of skin|Vascular disord of skin
C0162819|T047|PT|709.1|ICD9CM|Vascular disorders of skin|Vascular disorders of skin
C0036278|T020|AB|709.2|ICD9CM|Scar & fibrosis of skin|Scar & fibrosis of skin
C0036278|T020|PT|709.2|ICD9CM|Scar conditions and fibrosis of skin|Scar conditions and fibrosis of skin
C0342981|T047|AB|709.3|ICD9CM|Degenerative skin disord|Degenerative skin disord
C0342981|T047|PT|709.3|ICD9CM|Degenerative skin disorders|Degenerative skin disorders
C0157746|T047|AB|709.4|ICD9CM|Foreign body granul-skin|Foreign body granul-skin
C0157746|T047|PT|709.4|ICD9CM|Foreign body granuloma of skin and subcutaneous tissue|Foreign body granuloma of skin and subcutaneous tissue
C0029788|T047|PT|709.8|ICD9CM|Other specified disorders of skin|Other specified disorders of skin
C0029788|T047|AB|709.8|ICD9CM|Skin disorders NEC|Skin disorders NEC
C0178298|T047|AB|709.9|ICD9CM|Skin disorder NOS|Skin disorder NOS
C0178298|T047|PT|709.9|ICD9CM|Unspecified disorder of skin and subcutaneous tissue|Unspecified disorder of skin and subcutaneous tissue
C0041785|T047|HT|710|ICD9CM|Diffuse diseases of connective tissue|Diffuse diseases of connective tissue
C0178303|T047|HT|710-719.99|ICD9CM|ARTHROPATHIES AND RELATED DISORDERS|ARTHROPATHIES AND RELATED DISORDERS
C0263660|T047|HT|710-739.99|ICD9CM|DISEASES OF THE MUSCULOSKELETAL SYSTEM AND CONNECTIVE TISSUE|DISEASES OF THE MUSCULOSKELETAL SYSTEM AND CONNECTIVE TISSUE
C0024141|T047|AB|710.0|ICD9CM|Syst lupus erythematosus|Syst lupus erythematosus
C0024141|T047|PT|710.0|ICD9CM|Systemic lupus erythematosus|Systemic lupus erythematosus
C0036421|T047|AB|710.1|ICD9CM|Systemic sclerosis|Systemic sclerosis
C0036421|T047|PT|710.1|ICD9CM|Systemic sclerosis|Systemic sclerosis
C0086981|T047|AB|710.2|ICD9CM|Sicca syndrome|Sicca syndrome
C0086981|T047|PT|710.2|ICD9CM|Sicca syndrome|Sicca syndrome
C0011633|T047|AB|710.3|ICD9CM|Dermatomyositis|Dermatomyositis
C0011633|T047|PT|710.3|ICD9CM|Dermatomyositis|Dermatomyositis
C0085655|T047|AB|710.4|ICD9CM|Polymyositis|Polymyositis
C0085655|T047|PT|710.4|ICD9CM|Polymyositis|Polymyositis
C0085179|T047|AB|710.5|ICD9CM|Eosinophilia myalgia snd|Eosinophilia myalgia snd
C0085179|T047|PT|710.5|ICD9CM|Eosinophilia myalgia syndrome|Eosinophilia myalgia syndrome
C0157748|T047|AB|710.8|ICD9CM|Diff connect tis dis NEC|Diff connect tis dis NEC
C0157748|T047|PT|710.8|ICD9CM|Other specified diffuse diseases of connective tissue|Other specified diffuse diseases of connective tissue
C0041785|T047|AB|710.9|ICD9CM|Diff connect tis dis NOS|Diff connect tis dis NOS
C0041785|T047|PT|710.9|ICD9CM|Unspecified diffuse connective tissue disease|Unspecified diffuse connective tissue disease
C0157749|T047|HT|711|ICD9CM|Arthropathy associated with infections|Arthropathy associated with infections
C0003869|T047|HT|711.0|ICD9CM|Pyogenic arthritis|Pyogenic arthritis
C0343175|T047|AB|711.00|ICD9CM|Pyogen arthritis-unspec|Pyogen arthritis-unspec
C0343175|T047|PT|711.00|ICD9CM|Pyogenic arthritis, site unspecified|Pyogenic arthritis, site unspecified
C0263681|T047|AB|711.01|ICD9CM|Pyogen arthritis-shlder|Pyogen arthritis-shlder
C0263681|T047|PT|711.01|ICD9CM|Pyogenic arthritis, shoulder region|Pyogenic arthritis, shoulder region
C0263682|T047|AB|711.02|ICD9CM|Pyogen arthritis-up/arm|Pyogen arthritis-up/arm
C0263682|T047|PT|711.02|ICD9CM|Pyogenic arthritis, upper arm|Pyogenic arthritis, upper arm
C0263683|T047|AB|711.03|ICD9CM|Pyogen arthritis-forearm|Pyogen arthritis-forearm
C0263683|T047|PT|711.03|ICD9CM|Pyogenic arthritis, forearm|Pyogenic arthritis, forearm
C0263684|T047|AB|711.04|ICD9CM|Pyogen arthritis-hand|Pyogen arthritis-hand
C0263684|T047|PT|711.04|ICD9CM|Pyogenic arthritis, hand|Pyogenic arthritis, hand
C0409544|T047|AB|711.05|ICD9CM|Pyogen arthritis-pelvis|Pyogen arthritis-pelvis
C0409544|T047|PT|711.05|ICD9CM|Pyogenic arthritis, pelvic region and thigh|Pyogenic arthritis, pelvic region and thigh
C0263687|T047|AB|711.06|ICD9CM|Pyogen arthritis-l/leg|Pyogen arthritis-l/leg
C0263687|T047|PT|711.06|ICD9CM|Pyogenic arthritis, lower leg|Pyogenic arthritis, lower leg
C0157756|T047|AB|711.07|ICD9CM|Pyogen arthritis-ankle|Pyogen arthritis-ankle
C0157756|T047|PT|711.07|ICD9CM|Pyogenic arthritis, ankle and foot|Pyogenic arthritis, ankle and foot
C0409540|T047|AB|711.08|ICD9CM|Pyogen arthritis NEC|Pyogen arthritis NEC
C0409540|T047|PT|711.08|ICD9CM|Pyogenic arthritis, other specified sites|Pyogenic arthritis, other specified sites
C0263690|T047|AB|711.09|ICD9CM|Pyogen arthritis-mult|Pyogen arthritis-mult
C0263690|T047|PT|711.09|ICD9CM|Pyogenic arthritis, multiple sites|Pyogenic arthritis, multiple sites
C0157760|T047|HT|711.1|ICD9CM|Arthropathy associated with Reiter's disease and nonspecific urethritis|Arthropathy associated with Reiter's disease and nonspecific urethritis
C0157760|T047|PT|711.10|ICD9CM|Arthropathy associated with Reiter's disease and nonspecific urethritis, site unspecified|Arthropathy associated with Reiter's disease and nonspecific urethritis, site unspecified
C0157760|T047|AB|711.10|ICD9CM|Reiter arthritis-unspec|Reiter arthritis-unspec
C0157761|T047|PT|711.11|ICD9CM|Arthropathy associated with Reiter's disease and nonspecific urethritis, shoulder region|Arthropathy associated with Reiter's disease and nonspecific urethritis, shoulder region
C0157761|T047|AB|711.11|ICD9CM|Reiter arthritis-shlder|Reiter arthritis-shlder
C0157762|T047|PT|711.12|ICD9CM|Arthropathy associated with Reiter's disease and nonspecific urethritis, upper arm|Arthropathy associated with Reiter's disease and nonspecific urethritis, upper arm
C0157762|T047|AB|711.12|ICD9CM|Reiter arthritis-up/arm|Reiter arthritis-up/arm
C0157763|T047|PT|711.13|ICD9CM|Arthropathy associated with Reiter's disease and nonspecific urethritis, forearm|Arthropathy associated with Reiter's disease and nonspecific urethritis, forearm
C0157763|T047|AB|711.13|ICD9CM|Reiter arthritis-forearm|Reiter arthritis-forearm
C0157764|T047|PT|711.14|ICD9CM|Arthropathy associated with Reiter's disease and nonspecific urethritis, hand|Arthropathy associated with Reiter's disease and nonspecific urethritis, hand
C0157764|T047|AB|711.14|ICD9CM|Reiter arthritis-hand|Reiter arthritis-hand
C0157765|T047|PT|711.15|ICD9CM|Arthropathy associated with Reiter's disease and nonspecific urethritis, pelvic region and thigh|Arthropathy associated with Reiter's disease and nonspecific urethritis, pelvic region and thigh
C0157765|T047|AB|711.15|ICD9CM|Reiter arthritis-pelvis|Reiter arthritis-pelvis
C0157766|T047|PT|711.16|ICD9CM|Arthropathy associated with Reiter's disease and nonspecific urethritis, lower leg|Arthropathy associated with Reiter's disease and nonspecific urethritis, lower leg
C0157766|T047|AB|711.16|ICD9CM|Reiter arthritis-l/leg|Reiter arthritis-l/leg
C0157767|T047|PT|711.17|ICD9CM|Arthropathy associated with Reiter's disease and nonspecific urethritis, ankle and foot|Arthropathy associated with Reiter's disease and nonspecific urethritis, ankle and foot
C0157767|T047|AB|711.17|ICD9CM|Reiter arthritis-ankle|Reiter arthritis-ankle
C0157768|T047|PT|711.18|ICD9CM|Arthropathy associated with Reiter's disease and nonspecific urethritis, other specified sites|Arthropathy associated with Reiter's disease and nonspecific urethritis, other specified sites
C0157768|T047|AB|711.18|ICD9CM|Reiter arthritis NEC|Reiter arthritis NEC
C0157769|T047|PT|711.19|ICD9CM|Arthropathy associated with Reiter's disease and nonspecific urethritis, multiple sites|Arthropathy associated with Reiter's disease and nonspecific urethritis, multiple sites
C0157769|T047|AB|711.19|ICD9CM|Reiter arthritis-mult|Reiter arthritis-mult
C0157770|T047|HT|711.2|ICD9CM|Arthropathy in Behcet's syndrome|Arthropathy in Behcet's syndrome
C0157770|T047|PT|711.20|ICD9CM|Arthropathy in Behcet's syndrome, site unspecified|Arthropathy in Behcet's syndrome, site unspecified
C0157770|T047|AB|711.20|ICD9CM|Behcet arthritis-unspec|Behcet arthritis-unspec
C0409692|T047|PT|711.21|ICD9CM|Arthropathy in Behcet's syndrome, shoulder region|Arthropathy in Behcet's syndrome, shoulder region
C0409692|T047|AB|711.21|ICD9CM|Behcet arthritis-shlder|Behcet arthritis-shlder
C0409691|T047|PT|711.22|ICD9CM|Arthropathy in Behcet's syndrome, upper arm|Arthropathy in Behcet's syndrome, upper arm
C0409691|T047|AB|711.22|ICD9CM|Behcet arthritis-up/arm|Behcet arthritis-up/arm
C0409690|T047|PT|711.23|ICD9CM|Arthropathy in Behcet's syndrome, forearm|Arthropathy in Behcet's syndrome, forearm
C0409690|T047|AB|711.23|ICD9CM|Behcet arthritis-forearm|Behcet arthritis-forearm
C0409689|T047|PT|711.24|ICD9CM|Arthropathy in Behcet's syndrome, hand|Arthropathy in Behcet's syndrome, hand
C0409689|T047|AB|711.24|ICD9CM|Behcet arthritis-hand|Behcet arthritis-hand
C0409688|T047|PT|711.25|ICD9CM|Arthropathy in Behcet's syndrome, pelvic region and thigh|Arthropathy in Behcet's syndrome, pelvic region and thigh
C0409688|T047|AB|711.25|ICD9CM|Behcet arthritis-pelvis|Behcet arthritis-pelvis
C0409687|T047|PT|711.26|ICD9CM|Arthropathy in Behcet's syndrome, lower leg|Arthropathy in Behcet's syndrome, lower leg
C0409687|T047|AB|711.26|ICD9CM|Behcet arthritis-l/leg|Behcet arthritis-l/leg
C0409686|T047|PT|711.27|ICD9CM|Arthropathy in Behcet's syndrome, ankle and foot|Arthropathy in Behcet's syndrome, ankle and foot
C0409686|T047|AB|711.27|ICD9CM|Behcet arthritis-ankle|Behcet arthritis-ankle
C0409684|T047|PT|711.28|ICD9CM|Arthropathy in Behcet's syndrome, other specified sites|Arthropathy in Behcet's syndrome, other specified sites
C0409684|T047|AB|711.28|ICD9CM|Behcet arthritis NEC|Behcet arthritis NEC
C0409685|T047|PT|711.29|ICD9CM|Arthropathy in Behcet's syndrome, multiple sites|Arthropathy in Behcet's syndrome, multiple sites
C0409685|T047|AB|711.29|ICD9CM|Behcet arthritis-mult|Behcet arthritis-mult
C0152085|T046|HT|711.3|ICD9CM|Postdysenteric arthropathy|Postdysenteric arthropathy
C0152085|T046|AB|711.30|ICD9CM|Dysenter arthrit-unspec|Dysenter arthrit-unspec
C0152085|T046|PT|711.30|ICD9CM|Postdysenteric arthropathy, site unspecified|Postdysenteric arthropathy, site unspecified
C0837419|T047|AB|711.31|ICD9CM|Dysenter arthrit-shlder|Dysenter arthrit-shlder
C0837419|T047|PT|711.31|ICD9CM|Postdysenteric arthropathy, shoulder region|Postdysenteric arthropathy, shoulder region
C0837420|T047|AB|711.32|ICD9CM|Dysenter arthrit-up/arm|Dysenter arthrit-up/arm
C0837420|T047|PT|711.32|ICD9CM|Postdysenteric arthropathy, upper arm|Postdysenteric arthropathy, upper arm
C0837421|T047|AB|711.33|ICD9CM|Dysenter arthrit-forearm|Dysenter arthrit-forearm
C0837421|T047|PT|711.33|ICD9CM|Postdysenteric arthropathy, forearm|Postdysenteric arthropathy, forearm
C0837422|T046|AB|711.34|ICD9CM|Dysenter arthrit-hand|Dysenter arthrit-hand
C0837422|T046|PT|711.34|ICD9CM|Postdysenteric arthropathy, hand|Postdysenteric arthropathy, hand
C0837423|T047|AB|711.35|ICD9CM|Dysenter arthrit-pelvis|Dysenter arthrit-pelvis
C0837423|T047|PT|711.35|ICD9CM|Postdysenteric arthropathy, pelvic region and thigh|Postdysenteric arthropathy, pelvic region and thigh
C0837424|T047|AB|711.36|ICD9CM|Dysenter arthrit-l/leg|Dysenter arthrit-l/leg
C0837424|T047|PT|711.36|ICD9CM|Postdysenteric arthropathy, lower leg|Postdysenteric arthropathy, lower leg
C0837425|T046|AB|711.37|ICD9CM|Dysenter arthrit-ankle|Dysenter arthrit-ankle
C0837425|T046|PT|711.37|ICD9CM|Postdysenteric arthropathy, ankle and foot|Postdysenteric arthropathy, ankle and foot
C0157787|T047|AB|711.38|ICD9CM|Dysenter arthrit NEC|Dysenter arthrit NEC
C0157787|T047|PT|711.38|ICD9CM|Postdysenteric arthropathy, other specified sites|Postdysenteric arthropathy, other specified sites
C0837418|T046|AB|711.39|ICD9CM|Dysenter arthrit-mult|Dysenter arthrit-mult
C0837418|T046|PT|711.39|ICD9CM|Postdysenteric arthropathy, multiple sites|Postdysenteric arthropathy, multiple sites
C0157790|T047|HT|711.4|ICD9CM|Arthropathy associated with other bacterial diseases|Arthropathy associated with other bacterial diseases
C0157790|T047|PT|711.40|ICD9CM|Arthropathy associated with other bacterial diseases, site unspecified|Arthropathy associated with other bacterial diseases, site unspecified
C0157790|T047|AB|711.40|ICD9CM|Bact arthritis-unspec|Bact arthritis-unspec
C0409539|T047|PT|711.41|ICD9CM|Arthropathy associated with other bacterial diseases, shoulder region|Arthropathy associated with other bacterial diseases, shoulder region
C0409539|T047|AB|711.41|ICD9CM|Bact arthritis-shlder|Bact arthritis-shlder
C0409538|T047|PT|711.42|ICD9CM|Arthropathy associated with other bacterial diseases, upper arm|Arthropathy associated with other bacterial diseases, upper arm
C0409538|T047|AB|711.42|ICD9CM|Bact arthritis-up/arm|Bact arthritis-up/arm
C0409537|T047|PT|711.43|ICD9CM|Arthropathy associated with other bacterial diseases, forearm|Arthropathy associated with other bacterial diseases, forearm
C0409537|T047|AB|711.43|ICD9CM|Bact arthritis-forearm|Bact arthritis-forearm
C0409536|T047|PT|711.44|ICD9CM|Arthropathy associated with other bacterial diseases, hand|Arthropathy associated with other bacterial diseases, hand
C0409536|T047|AB|711.44|ICD9CM|Bact arthritis-hand|Bact arthritis-hand
C0409535|T047|PT|711.45|ICD9CM|Arthropathy associated with other bacterial diseases, pelvic region and thigh|Arthropathy associated with other bacterial diseases, pelvic region and thigh
C0409535|T047|AB|711.45|ICD9CM|Bact arthritis-pelvis|Bact arthritis-pelvis
C0409534|T047|PT|711.46|ICD9CM|Arthropathy associated with other bacterial diseases, lower leg|Arthropathy associated with other bacterial diseases, lower leg
C0409534|T047|AB|711.46|ICD9CM|Bact arthritis-l/leg|Bact arthritis-l/leg
C0409533|T047|PT|711.47|ICD9CM|Arthropathy associated with other bacterial diseases, ankle and foot|Arthropathy associated with other bacterial diseases, ankle and foot
C0409533|T047|AB|711.47|ICD9CM|Bact arthritis-ankle|Bact arthritis-ankle
C0409531|T047|PT|711.48|ICD9CM|Arthropathy associated with other bacterial diseases, other specified sites|Arthropathy associated with other bacterial diseases, other specified sites
C0409531|T047|AB|711.48|ICD9CM|Bact arthritis NEC|Bact arthritis NEC
C0409532|T047|PT|711.49|ICD9CM|Arthropathy associated with other bacterial diseases, multiple sites|Arthropathy associated with other bacterial diseases, multiple sites
C0409532|T047|AB|711.49|ICD9CM|Bact arthritis-mult|Bact arthritis-mult
C0157801|T047|HT|711.5|ICD9CM|Arthropathy associated with other viral diseases|Arthropathy associated with other viral diseases
C0157801|T047|PT|711.50|ICD9CM|Arthropathy associated with other viral diseases, site unspecified|Arthropathy associated with other viral diseases, site unspecified
C0157801|T047|AB|711.50|ICD9CM|Viral arthritis-unspec|Viral arthritis-unspec
C0409556|T047|PT|711.51|ICD9CM|Arthropathy associated with other viral diseases, shoulder region|Arthropathy associated with other viral diseases, shoulder region
C0409556|T047|AB|711.51|ICD9CM|Viral arthritis-shlder|Viral arthritis-shlder
C0409555|T047|PT|711.52|ICD9CM|Arthropathy associated with other viral diseases, upper arm|Arthropathy associated with other viral diseases, upper arm
C0409555|T047|AB|711.52|ICD9CM|Viral arthritis-up/arm|Viral arthritis-up/arm
C0409554|T047|PT|711.53|ICD9CM|Arthropathy associated with other viral diseases, forearm|Arthropathy associated with other viral diseases, forearm
C0409554|T047|AB|711.53|ICD9CM|Viral arthritis-forearm|Viral arthritis-forearm
C0157805|T047|PT|711.54|ICD9CM|Arthropathy associated with other viral diseases, hand|Arthropathy associated with other viral diseases, hand
C0157805|T047|AB|711.54|ICD9CM|Viral arthritis-hand|Viral arthritis-hand
C0409552|T047|PT|711.55|ICD9CM|Arthropathy associated with other viral diseases, pelvic region and thigh|Arthropathy associated with other viral diseases, pelvic region and thigh
C0409552|T047|AB|711.55|ICD9CM|Viral arthritis-pelvis|Viral arthritis-pelvis
C0409551|T047|PT|711.56|ICD9CM|Arthropathy associated with other viral diseases, lower leg|Arthropathy associated with other viral diseases, lower leg
C0409551|T047|AB|711.56|ICD9CM|Viral arthritis-l/leg|Viral arthritis-l/leg
C0409550|T047|PT|711.57|ICD9CM|Arthropathy associated with other viral diseases, ankle and foot|Arthropathy associated with other viral diseases, ankle and foot
C0409550|T047|AB|711.57|ICD9CM|Viral arthritis-ankle|Viral arthritis-ankle
C0409548|T047|PT|711.58|ICD9CM|Arthropathy associated with other viral diseases, other specified sites|Arthropathy associated with other viral diseases, other specified sites
C0409548|T047|AB|711.58|ICD9CM|Viral arthritis NEC|Viral arthritis NEC
C0409549|T047|PT|711.59|ICD9CM|Arthropathy associated with other viral diseases, multiple sites|Arthropathy associated with other viral diseases, multiple sites
C0409549|T047|AB|711.59|ICD9CM|Viral arthritis-mult|Viral arthritis-mult
C0869528|T047|HT|711.6|ICD9CM|Arthropathy associated with mycoses|Arthropathy associated with mycoses
C0869528|T047|PT|711.60|ICD9CM|Arthropathy associated with mycoses, site unspecified|Arthropathy associated with mycoses, site unspecified
C0869528|T047|AB|711.60|ICD9CM|Mycotic arthritis-unspec|Mycotic arthritis-unspec
C0409567|T047|PT|711.61|ICD9CM|Arthropathy associated with mycoses, shoulder region|Arthropathy associated with mycoses, shoulder region
C0409567|T047|AB|711.61|ICD9CM|Mycotic arthritis-shlder|Mycotic arthritis-shlder
C0409566|T047|PT|711.62|ICD9CM|Arthropathy associated with mycoses, upper arm|Arthropathy associated with mycoses, upper arm
C0409566|T047|AB|711.62|ICD9CM|Mycotic arthritis-up/arm|Mycotic arthritis-up/arm
C0409565|T047|PT|711.63|ICD9CM|Arthropathy associated with mycoses, forearm|Arthropathy associated with mycoses, forearm
C0409565|T047|AB|711.63|ICD9CM|Mycotic arthrit-forearm|Mycotic arthrit-forearm
C0409564|T047|PT|711.64|ICD9CM|Arthropathy associated with mycoses, hand|Arthropathy associated with mycoses, hand
C0409564|T047|AB|711.64|ICD9CM|Mycotic arthritis-hand|Mycotic arthritis-hand
C0409563|T047|PT|711.65|ICD9CM|Arthropathy associated with mycoses, pelvic region and thigh|Arthropathy associated with mycoses, pelvic region and thigh
C0409563|T047|AB|711.65|ICD9CM|Mycotic arthritis-pelvis|Mycotic arthritis-pelvis
C0409562|T047|PT|711.66|ICD9CM|Arthropathy associated with mycoses, lower leg|Arthropathy associated with mycoses, lower leg
C0409562|T047|AB|711.66|ICD9CM|Mycotic arthritis-l/leg|Mycotic arthritis-l/leg
C0409561|T047|PT|711.67|ICD9CM|Arthropathy associated with mycoses, ankle and foot|Arthropathy associated with mycoses, ankle and foot
C0409561|T047|AB|711.67|ICD9CM|Mycotic arthritis-ankle|Mycotic arthritis-ankle
C0409559|T047|PT|711.68|ICD9CM|Arthropathy associated with mycoses, other specified sites|Arthropathy associated with mycoses, other specified sites
C0409559|T047|AB|711.68|ICD9CM|Mycotic arthritis NEC|Mycotic arthritis NEC
C0157821|T047|PT|711.69|ICD9CM|Arthropathy associated with mycoses, involving multiple sites|Arthropathy associated with mycoses, involving multiple sites
C0157821|T047|AB|711.69|ICD9CM|Mycotic arthritis-mult|Mycotic arthritis-mult
C0157822|T047|HT|711.7|ICD9CM|Arthropathy associated with helminthiasis|Arthropathy associated with helminthiasis
C0409569|T047|PT|711.70|ICD9CM|Arthropathy associated with helminthiasis, site unspecified|Arthropathy associated with helminthiasis, site unspecified
C0409569|T047|AB|711.70|ICD9CM|Helminth arthrit-unspec|Helminth arthrit-unspec
C0157824|T047|PT|711.71|ICD9CM|Arthropathy associated with helminthiasis, shoulder region|Arthropathy associated with helminthiasis, shoulder region
C0157824|T047|AB|711.71|ICD9CM|Helminth arthrit-shlder|Helminth arthrit-shlder
C0409577|T047|PT|711.72|ICD9CM|Arthropathy associated with helminthiasis, upper arm|Arthropathy associated with helminthiasis, upper arm
C0409577|T047|AB|711.72|ICD9CM|Helminth arthrit-up/arm|Helminth arthrit-up/arm
C0409576|T047|PT|711.73|ICD9CM|Arthropathy associated with helminthiasis, forearm|Arthropathy associated with helminthiasis, forearm
C0409576|T047|AB|711.73|ICD9CM|Helminth arthrit-forearm|Helminth arthrit-forearm
C0409575|T047|PT|711.74|ICD9CM|Arthropathy associated with helminthiasis, hand|Arthropathy associated with helminthiasis, hand
C0409575|T047|AB|711.74|ICD9CM|Helminth arthrit-hand|Helminth arthrit-hand
C0409574|T047|PT|711.75|ICD9CM|Arthropathy associated with helminthiasis, pelvic region and thigh|Arthropathy associated with helminthiasis, pelvic region and thigh
C0409574|T047|AB|711.75|ICD9CM|Helminth arthrit-pelvis|Helminth arthrit-pelvis
C0409573|T047|PT|711.76|ICD9CM|Arthropathy associated with helminthiasis, lower leg|Arthropathy associated with helminthiasis, lower leg
C0409573|T047|AB|711.76|ICD9CM|Helminth arthrit-l/leg|Helminth arthrit-l/leg
C0409572|T047|PT|711.77|ICD9CM|Arthropathy associated with helminthiasis, ankle and foot|Arthropathy associated with helminthiasis, ankle and foot
C0409572|T047|AB|711.77|ICD9CM|Helminth arthrit-ankle|Helminth arthrit-ankle
C0409570|T047|PT|711.78|ICD9CM|Arthropathy associated with helminthiasis, other specified sites|Arthropathy associated with helminthiasis, other specified sites
C0409570|T047|AB|711.78|ICD9CM|Helminth arthrit NEC|Helminth arthrit NEC
C0409571|T047|PT|711.79|ICD9CM|Arthropathy associated with helminthiasis, multiple sites|Arthropathy associated with helminthiasis, multiple sites
C0409571|T047|AB|711.79|ICD9CM|Helminth arthrit-mult|Helminth arthrit-mult
C0157833|T047|HT|711.8|ICD9CM|Arthropathy associated with other infectious and parasitic diseases|Arthropathy associated with other infectious and parasitic diseases
C0157833|T047|PT|711.80|ICD9CM|Arthropathy associated with other infectious and parasitic diseases, site unspecified|Arthropathy associated with other infectious and parasitic diseases, site unspecified
C0157833|T047|AB|711.80|ICD9CM|Inf arthritis NEC-unspec|Inf arthritis NEC-unspec
C0157834|T047|PT|711.81|ICD9CM|Arthropathy associated with other infectious and parasitic diseases, shoulder region|Arthropathy associated with other infectious and parasitic diseases, shoulder region
C0157834|T047|AB|711.81|ICD9CM|Inf arthritis NEC-shlder|Inf arthritis NEC-shlder
C0157835|T047|PT|711.82|ICD9CM|Arthropathy associated with other infectious and parasitic diseases, upper arm|Arthropathy associated with other infectious and parasitic diseases, upper arm
C0157835|T047|AB|711.82|ICD9CM|Inf arthritis NEC-up/arm|Inf arthritis NEC-up/arm
C0157836|T047|PT|711.83|ICD9CM|Arthropathy associated with other infectious and parasitic diseases, forearm|Arthropathy associated with other infectious and parasitic diseases, forearm
C0157836|T047|AB|711.83|ICD9CM|Inf arthrit NEC-forearm|Inf arthrit NEC-forearm
C0157837|T047|PT|711.84|ICD9CM|Arthropathy associated with other infectious and parasitic diseases, hand|Arthropathy associated with other infectious and parasitic diseases, hand
C0157837|T047|AB|711.84|ICD9CM|Inf arthritis NEC-hand|Inf arthritis NEC-hand
C0157838|T047|PT|711.85|ICD9CM|Arthropathy associated with other infectious and parasitic diseases, pelvic region and thigh|Arthropathy associated with other infectious and parasitic diseases, pelvic region and thigh
C0157838|T047|AB|711.85|ICD9CM|Inf arthritis NEC-pelvis|Inf arthritis NEC-pelvis
C0157839|T047|PT|711.86|ICD9CM|Arthropathy associated with other infectious and parasitic diseases, lower leg|Arthropathy associated with other infectious and parasitic diseases, lower leg
C0157839|T047|AB|711.86|ICD9CM|Inf arthritis NEC-l/leg|Inf arthritis NEC-l/leg
C0157840|T047|PT|711.87|ICD9CM|Arthropathy associated with other infectious and parasitic diseases, ankle and foot|Arthropathy associated with other infectious and parasitic diseases, ankle and foot
C0157840|T047|AB|711.87|ICD9CM|Inf arthritis NEC-ankle|Inf arthritis NEC-ankle
C0157841|T047|PT|711.88|ICD9CM|Arthropathy associated with other infectious and parasitic diseases, other specified sites|Arthropathy associated with other infectious and parasitic diseases, other specified sites
C0157841|T047|AB|711.88|ICD9CM|Inf arthrit NEC-oth site|Inf arthrit NEC-oth site
C0157842|T047|PT|711.89|ICD9CM|Arthropathy associated with other infectious and parasitic diseases, multiple sites|Arthropathy associated with other infectious and parasitic diseases, multiple sites
C0157842|T047|AB|711.89|ICD9CM|Inf arthritis NEC-mult|Inf arthritis NEC-mult
C0003869|T047|HT|711.9|ICD9CM|Unspecified infective arthritis|Unspecified infective arthritis
C0003869|T047|AB|711.90|ICD9CM|Inf arthritis NOS-unspec|Inf arthritis NOS-unspec
C0003869|T047|PT|711.90|ICD9CM|Unspecified infective arthritis, site unspecified|Unspecified infective arthritis, site unspecified
C0157843|T047|AB|711.91|ICD9CM|Inf arthritis NOS-shlder|Inf arthritis NOS-shlder
C0157843|T047|PT|711.91|ICD9CM|Unspecified infective arthritis, shoulder region|Unspecified infective arthritis, shoulder region
C0157844|T047|AB|711.92|ICD9CM|Inf arthritis NOS-up/arm|Inf arthritis NOS-up/arm
C0157844|T047|PT|711.92|ICD9CM|Unspecified infective arthritis, upper arm|Unspecified infective arthritis, upper arm
C0157845|T047|AB|711.93|ICD9CM|Inf arthrit NOS-forearm|Inf arthrit NOS-forearm
C0157845|T047|PT|711.93|ICD9CM|Unspecified infective arthritis, forearm|Unspecified infective arthritis, forearm
C0157846|T047|AB|711.94|ICD9CM|Inf arthrit NOS-hand|Inf arthrit NOS-hand
C0157846|T047|PT|711.94|ICD9CM|Unspecified infective arthritis, hand|Unspecified infective arthritis, hand
C0157847|T047|AB|711.95|ICD9CM|Inf arthrit NOS-pelvis|Inf arthrit NOS-pelvis
C0157847|T047|PT|711.95|ICD9CM|Unspecified infective arthritis, pelvic region and thigh|Unspecified infective arthritis, pelvic region and thigh
C0157848|T047|AB|711.96|ICD9CM|Inf arthrit NOS-l/leg|Inf arthrit NOS-l/leg
C0157848|T047|PT|711.96|ICD9CM|Unspecified infective arthritis, lower leg|Unspecified infective arthritis, lower leg
C0157849|T047|AB|711.97|ICD9CM|Inf arthrit NOS-ankle|Inf arthrit NOS-ankle
C0157849|T047|PT|711.97|ICD9CM|Unspecified infective arthritis, ankle and foot|Unspecified infective arthritis, ankle and foot
C0157850|T047|AB|711.98|ICD9CM|Inf arthrit NOS-oth site|Inf arthrit NOS-oth site
C0157850|T047|PT|711.98|ICD9CM|Unspecified infective arthritis, other specified sites|Unspecified infective arthritis, other specified sites
C0157851|T047|AB|711.99|ICD9CM|Inf arthritis NOS-mult|Inf arthritis NOS-mult
C0157851|T047|PT|711.99|ICD9CM|Unspecified infective arthritis, multiple sites|Unspecified infective arthritis, multiple sites
C0152087|T047|HT|712|ICD9CM|Crystal arthropathies|Crystal arthropathies
C0157852|T047|HT|712.1|ICD9CM|Chondrocalcinosis due to dicalcium phosphate crystals|Chondrocalcinosis due to dicalcium phosphate crystals
C0409882|T047|PT|712.10|ICD9CM|Chondrocalcinosis, due to dicalcium phosphate crystals, site unspecified|Chondrocalcinosis, due to dicalcium phosphate crystals, site unspecified
C0409882|T047|AB|712.10|ICD9CM|Dicalc phos cryst-unspec|Dicalc phos cryst-unspec
C0409881|T047|PT|712.11|ICD9CM|Chondrocalcinosis, due to dicalcium phosphate crystals, shoulder region|Chondrocalcinosis, due to dicalcium phosphate crystals, shoulder region
C0409881|T047|AB|712.11|ICD9CM|Dicalc phos cryst-shlder|Dicalc phos cryst-shlder
C0409880|T047|PT|712.12|ICD9CM|Chondrocalcinosis, due to dicalcium phosphate crystals, upper arm|Chondrocalcinosis, due to dicalcium phosphate crystals, upper arm
C0409880|T047|AB|712.12|ICD9CM|Dicalc phos cryst-up/arm|Dicalc phos cryst-up/arm
C0409879|T047|PT|712.13|ICD9CM|Chondrocalcinosis, due to dicalcium phosphate crystals, forearm|Chondrocalcinosis, due to dicalcium phosphate crystals, forearm
C0409879|T047|AB|712.13|ICD9CM|Dicalc phos crys-forearm|Dicalc phos crys-forearm
C0409878|T047|PT|712.14|ICD9CM|Chondrocalcinosis, due to dicalcium phosphate crystals, hand|Chondrocalcinosis, due to dicalcium phosphate crystals, hand
C0409878|T047|AB|712.14|ICD9CM|Dicalc phos cryst-hand|Dicalc phos cryst-hand
C0409877|T047|PT|712.15|ICD9CM|Chondrocalcinosis, due to dicalcium phosphate crystals, pelvic region and thigh|Chondrocalcinosis, due to dicalcium phosphate crystals, pelvic region and thigh
C0409877|T047|AB|712.15|ICD9CM|Dicalc phos cryst-pelvis|Dicalc phos cryst-pelvis
C0409876|T047|PT|712.16|ICD9CM|Chondrocalcinosis, due to dicalcium phosphate crystals, lower leg|Chondrocalcinosis, due to dicalcium phosphate crystals, lower leg
C0409876|T047|AB|712.16|ICD9CM|Dicalc phos cryst-l/leg|Dicalc phos cryst-l/leg
C0409875|T047|PT|712.17|ICD9CM|Chondrocalcinosis, due to dicalcium phosphate crystals, ankle and foot|Chondrocalcinosis, due to dicalcium phosphate crystals, ankle and foot
C0409875|T047|AB|712.17|ICD9CM|Dicalc phos cryst-ankle|Dicalc phos cryst-ankle
C0409873|T047|PT|712.18|ICD9CM|Chondrocalcinosis, due to dicalcium phosphate crystals, other specified sites|Chondrocalcinosis, due to dicalcium phosphate crystals, other specified sites
C0409873|T047|AB|712.18|ICD9CM|Dicalc phos cry-site NEC|Dicalc phos cry-site NEC
C0409874|T047|PT|712.19|ICD9CM|Chondrocalcinosis, due to dicalcium phosphate crystals, multiple sites|Chondrocalcinosis, due to dicalcium phosphate crystals, multiple sites
C0409874|T047|AB|712.19|ICD9CM|Dicalc phos cryst-mult|Dicalc phos cryst-mult
C0553730|T047|HT|712.2|ICD9CM|Chondrocalcinosis due to pyrophosphate crystals|Chondrocalcinosis due to pyrophosphate crystals
C0553730|T047|PT|712.20|ICD9CM|Chondrocalcinosis, due to pyrophosphate crystals, site unspecified|Chondrocalcinosis, due to pyrophosphate crystals, site unspecified
C0553730|T047|AB|712.20|ICD9CM|Pyrophosph cryst-unspec|Pyrophosph cryst-unspec
C0409871|T047|PT|712.21|ICD9CM|Chondrocalcinosis, due to pyrophosphate crystals, shoulder region|Chondrocalcinosis, due to pyrophosphate crystals, shoulder region
C0409871|T047|AB|712.21|ICD9CM|Pyrophosph cryst-shlder|Pyrophosph cryst-shlder
C0409870|T047|PT|712.22|ICD9CM|Chondrocalcinosis, due to pyrophosphate crystals, upper arm|Chondrocalcinosis, due to pyrophosphate crystals, upper arm
C0409870|T047|AB|712.22|ICD9CM|Pyrophosph cryst-up/arm|Pyrophosph cryst-up/arm
C0409869|T047|PT|712.23|ICD9CM|Chondrocalcinosis, due to pyrophosphate crystals, forearm|Chondrocalcinosis, due to pyrophosphate crystals, forearm
C0409869|T047|AB|712.23|ICD9CM|Pyrophosph cryst-forearm|Pyrophosph cryst-forearm
C0409868|T047|PT|712.24|ICD9CM|Chondrocalcinosis, due to pyrophosphate crystals, hand|Chondrocalcinosis, due to pyrophosphate crystals, hand
C0409868|T047|AB|712.24|ICD9CM|Pyrophosph cryst-hand|Pyrophosph cryst-hand
C0409867|T047|PT|712.25|ICD9CM|Chondrocalcinosis, due to pyrophosphate crystals, pelvic region and thigh|Chondrocalcinosis, due to pyrophosphate crystals, pelvic region and thigh
C0409867|T047|AB|712.25|ICD9CM|Pyrophosph cryst-pelvis|Pyrophosph cryst-pelvis
C0409865|T047|PT|712.26|ICD9CM|Chondrocalcinosis, due to pyrophosphate crystals, lower leg|Chondrocalcinosis, due to pyrophosphate crystals, lower leg
C0409865|T047|AB|712.26|ICD9CM|Pyrophosph cryst-l/leg|Pyrophosph cryst-l/leg
C0409864|T047|PT|712.27|ICD9CM|Chondrocalcinosis, due to pyrophosphate crystals, ankle and foot|Chondrocalcinosis, due to pyrophosphate crystals, ankle and foot
C0409864|T047|AB|712.27|ICD9CM|Pyrophosph cryst-ankle|Pyrophosph cryst-ankle
C0409862|T047|PT|712.28|ICD9CM|Chondrocalcinosis, due to pyrophosphate crystals, other specified sites|Chondrocalcinosis, due to pyrophosphate crystals, other specified sites
C0409862|T047|AB|712.28|ICD9CM|Pyrophos cryst-site NEC|Pyrophos cryst-site NEC
C0409863|T047|PT|712.29|ICD9CM|Chondrocalcinosis, due to pyrophosphate crystals, multiple sites|Chondrocalcinosis, due to pyrophosphate crystals, multiple sites
C0409863|T047|AB|712.29|ICD9CM|Pyrophos cryst-mult|Pyrophos cryst-mult
C0553730|T047|HT|712.3|ICD9CM|Chondrocalcinosis, cause unspecified|Chondrocalcinosis, cause unspecified
C0157874|T047|AB|712.30|ICD9CM|Chondrocalcin NOS-unspec|Chondrocalcin NOS-unspec
C0157874|T047|PT|712.30|ICD9CM|Chondrocalcinosis, unspecified, site unspecified|Chondrocalcinosis, unspecified, site unspecified
C0409894|T047|AB|712.31|ICD9CM|Chondrocalcin NOS-shlder|Chondrocalcin NOS-shlder
C0409894|T047|PT|712.31|ICD9CM|Chondrocalcinosis, unspecified, shoulder region|Chondrocalcinosis, unspecified, shoulder region
C0409893|T047|AB|712.32|ICD9CM|Chondrocalcin NOS-up/arm|Chondrocalcin NOS-up/arm
C0409893|T047|PT|712.32|ICD9CM|Chondrocalcinosis, unspecified, upper arm|Chondrocalcinosis, unspecified, upper arm
C0409892|T047|AB|712.33|ICD9CM|Chondrocalc NOS-forearm|Chondrocalc NOS-forearm
C0409892|T047|PT|712.33|ICD9CM|Chondrocalcinosis, unspecified, forearm|Chondrocalcinosis, unspecified, forearm
C0409891|T047|AB|712.34|ICD9CM|Chondrocalcin NOS-hand|Chondrocalcin NOS-hand
C0409891|T047|PT|712.34|ICD9CM|Chondrocalcinosis, unspecified, hand|Chondrocalcinosis, unspecified, hand
C0409890|T047|AB|712.35|ICD9CM|Chondrocalcin NOS-pelvis|Chondrocalcin NOS-pelvis
C0409890|T047|PT|712.35|ICD9CM|Chondrocalcinosis, unspecified, pelvic region and thigh|Chondrocalcinosis, unspecified, pelvic region and thigh
C0409889|T047|AB|712.36|ICD9CM|Chondrocalcin NOS-l/leg|Chondrocalcin NOS-l/leg
C0409889|T047|PT|712.36|ICD9CM|Chondrocalcinosis, unspecified, lower leg|Chondrocalcinosis, unspecified, lower leg
C0409888|T047|AB|712.37|ICD9CM|Chondrocalcin NOS-ankle|Chondrocalcin NOS-ankle
C0409888|T047|PT|712.37|ICD9CM|Chondrocalcinosis, unspecified, ankle and foot|Chondrocalcinosis, unspecified, ankle and foot
C0409886|T047|AB|712.38|ICD9CM|Chondrocalc NOS-oth site|Chondrocalc NOS-oth site
C0409886|T047|PT|712.38|ICD9CM|Chondrocalcinosis, unspecified, other specified sites|Chondrocalcinosis, unspecified, other specified sites
C0409887|T047|AB|712.39|ICD9CM|Chondrocalcin NOS-mult|Chondrocalcin NOS-mult
C0409887|T047|PT|712.39|ICD9CM|Chondrocalcinosis, unspecified, multiple sites|Chondrocalcinosis, unspecified, multiple sites
C0157884|T047|HT|712.8|ICD9CM|Other specified crystal arthropathies|Other specified crystal arthropathies
C0157884|T047|AB|712.80|ICD9CM|Cryst arthrop NEC-unspec|Cryst arthrop NEC-unspec
C0157884|T047|PT|712.80|ICD9CM|Other specified crystal arthropathies, site unspecified|Other specified crystal arthropathies, site unspecified
C0837882|T047|AB|712.81|ICD9CM|Cryst arthrop NEC-shlder|Cryst arthrop NEC-shlder
C0837882|T047|PT|712.81|ICD9CM|Other specified crystal arthropathies, shoulder region|Other specified crystal arthropathies, shoulder region
C0837883|T047|AB|712.82|ICD9CM|Cryst arthrop NEC-up/arm|Cryst arthrop NEC-up/arm
C0837883|T047|PT|712.82|ICD9CM|Other specified crystal arthropathies, upper arm|Other specified crystal arthropathies, upper arm
C0837884|T047|AB|712.83|ICD9CM|Crys arthrop NEC-forearm|Crys arthrop NEC-forearm
C0837884|T047|PT|712.83|ICD9CM|Other specified crystal arthropathies, forearm|Other specified crystal arthropathies, forearm
C0837885|T047|AB|712.84|ICD9CM|Cryst arthrop NEC-hand|Cryst arthrop NEC-hand
C0837885|T047|PT|712.84|ICD9CM|Other specified crystal arthropathies, hand|Other specified crystal arthropathies, hand
C0837886|T047|AB|712.85|ICD9CM|Cryst arthrop NEC-pelvis|Cryst arthrop NEC-pelvis
C0837886|T047|PT|712.85|ICD9CM|Other specified crystal arthropathies, pelvic region and thigh|Other specified crystal arthropathies, pelvic region and thigh
C0837887|T047|AB|712.86|ICD9CM|Cryst arthrop NEC-l/leg|Cryst arthrop NEC-l/leg
C0837887|T047|PT|712.86|ICD9CM|Other specified crystal arthropathies, lower leg|Other specified crystal arthropathies, lower leg
C0837888|T047|AB|712.87|ICD9CM|Cryst arthrop NEC-ankle|Cryst arthrop NEC-ankle
C0837888|T047|PT|712.87|ICD9CM|Other specified crystal arthropathies, ankle and foot|Other specified crystal arthropathies, ankle and foot
C0157892|T047|AB|712.88|ICD9CM|Cry arthrop NEC-oth site|Cry arthrop NEC-oth site
C0157892|T047|PT|712.88|ICD9CM|Other specified crystal arthropathies, other specified sites|Other specified crystal arthropathies, other specified sites
C0837881|T047|AB|712.89|ICD9CM|Cryst arthrop NEC-mult|Cryst arthrop NEC-mult
C0837881|T047|PT|712.89|ICD9CM|Other specified crystal arthropathies, multiple sites|Other specified crystal arthropathies, multiple sites
C0152087|T047|HT|712.9|ICD9CM|Unspecified crystal arthropathy|Unspecified crystal arthropathy
C0152087|T047|AB|712.90|ICD9CM|Cryst arthrop NOS-unspec|Cryst arthrop NOS-unspec
C0152087|T047|PT|712.90|ICD9CM|Unspecified crystal arthropathy, site unspecified|Unspecified crystal arthropathy, site unspecified
C0263708|T047|AB|712.91|ICD9CM|Cryst arthrop NOS-shldr|Cryst arthrop NOS-shldr
C0263708|T047|PT|712.91|ICD9CM|Unspecified crystal arthropathy, shoulder region|Unspecified crystal arthropathy, shoulder region
C0263709|T047|AB|712.92|ICD9CM|Cryst arthrop NOS-up/arm|Cryst arthrop NOS-up/arm
C0263709|T047|PT|712.92|ICD9CM|Unspecified crystal arthropathy, upper arm|Unspecified crystal arthropathy, upper arm
C0263710|T047|AB|712.93|ICD9CM|Crys arthrop NOS-forearm|Crys arthrop NOS-forearm
C0263710|T047|PT|712.93|ICD9CM|Unspecified crystal arthropathy, forearm|Unspecified crystal arthropathy, forearm
C0263711|T047|AB|712.94|ICD9CM|Cryst arthrop NOS-hand|Cryst arthrop NOS-hand
C0263711|T047|PT|712.94|ICD9CM|Unspecified crystal arthropathy, hand|Unspecified crystal arthropathy, hand
C0409843|T047|AB|712.95|ICD9CM|Cryst arthrop NOS-pelvis|Cryst arthrop NOS-pelvis
C0409843|T047|PT|712.95|ICD9CM|Unspecified crystal arthropathy, pelvic region and thigh|Unspecified crystal arthropathy, pelvic region and thigh
C0263714|T047|AB|712.96|ICD9CM|Cryst arthrop NOS-l/leg|Cryst arthrop NOS-l/leg
C0263714|T047|PT|712.96|ICD9CM|Unspecified crystal arthropathy, lower leg|Unspecified crystal arthropathy, lower leg
C0263715|T047|AB|712.97|ICD9CM|Cryst arthrop NOS-ankle|Cryst arthrop NOS-ankle
C0263715|T047|PT|712.97|ICD9CM|Unspecified crystal arthropathy, ankle and foot|Unspecified crystal arthropathy, ankle and foot
C0263716|T047|AB|712.98|ICD9CM|Cry arthrop NOS-oth site|Cry arthrop NOS-oth site
C0263716|T047|PT|712.98|ICD9CM|Unspecified crystal arthropathy, other specified sites|Unspecified crystal arthropathy, other specified sites
C0263717|T047|AB|712.99|ICD9CM|Cryst arthrop NOS-mult|Cryst arthrop NOS-mult
C0263717|T047|PT|712.99|ICD9CM|Unspecified crystal arthropathy, multiple sites|Unspecified crystal arthropathy, multiple sites
C0157904|T047|HT|713|ICD9CM|Arthropathy associated with other disorders classified elsewhere|Arthropathy associated with other disorders classified elsewhere
C0409729|T047|AB|713.0|ICD9CM|Arthrop w endocr/met dis|Arthrop w endocr/met dis
C0409729|T047|PT|713.0|ICD9CM|Arthropathy associated with other endocrine and metabolic disorders|Arthropathy associated with other endocrine and metabolic disorders
C0263723|T047|AB|713.1|ICD9CM|Arthrop w noninf GI dis|Arthrop w noninf GI dis
C0263723|T047|PT|713.1|ICD9CM|Arthropathy associated with gastrointestinal conditions other than infections|Arthropathy associated with gastrointestinal conditions other than infections
C0263724|T047|AB|713.2|ICD9CM|Arthropath w hematol dis|Arthropath w hematol dis
C0263724|T047|PT|713.2|ICD9CM|Arthropathy associated with hematological disorders|Arthropathy associated with hematological disorders
C0263726|T047|PT|713.3|ICD9CM|Arthropathy associated with dermatological disorders|Arthropathy associated with dermatological disorders
C0263726|T047|AB|713.3|ICD9CM|Arthropathy w skin dis|Arthropathy w skin dis
C0263727|T047|PT|713.4|ICD9CM|Arthropathy associated with respiratory disorders|Arthropathy associated with respiratory disorders
C0263727|T047|AB|713.4|ICD9CM|Arthropathy w resp dis|Arthropathy w resp dis
C0003892|T047|PT|713.5|ICD9CM|Arthropathy associated with neurological disorders|Arthropathy associated with neurological disorders
C0003892|T047|AB|713.5|ICD9CM|Arthropathy w nerve dis|Arthropathy w nerve dis
C0263730|T047|AB|713.6|ICD9CM|Arthrop w hypersen react|Arthrop w hypersen react
C0263730|T047|PT|713.6|ICD9CM|Arthropathy associated with hypersensitivity reaction|Arthropathy associated with hypersensitivity reaction
C0157911|T047|AB|713.7|ICD9CM|Arthrop w system dis NEC|Arthrop w system dis NEC
C0157911|T047|PT|713.7|ICD9CM|Other general diseases with articular involvement|Other general diseases with articular involvement
C0263732|T047|AB|713.8|ICD9CM|Arthrop w oth dis NEC|Arthrop w oth dis NEC
C0263732|T047|PT|713.8|ICD9CM|Arthropathy associated with other conditions classifiable elsewhere|Arthropathy associated with other conditions classifiable elsewhere
C0157913|T047|HT|714|ICD9CM|Rheumatoid arthritis and other inflammatory polyarthropathies|Rheumatoid arthritis and other inflammatory polyarthropathies
C0003873|T047|AB|714.0|ICD9CM|Rheumatoid arthritis|Rheumatoid arthritis
C0003873|T047|PT|714.0|ICD9CM|Rheumatoid arthritis|Rheumatoid arthritis
C0015773|T047|AB|714.1|ICD9CM|Felty's syndrome|Felty's syndrome
C0015773|T047|PT|714.1|ICD9CM|Felty's syndrome|Felty's syndrome
C0157914|T047|PT|714.2|ICD9CM|Other rheumatoid arthritis with visceral or systemic involvement|Other rheumatoid arthritis with visceral or systemic involvement
C0157914|T047|AB|714.2|ICD9CM|Syst rheum arthritis NEC|Syst rheum arthritis NEC
C0409667|T047|HT|714.3|ICD9CM|Juvenile chronic polyarthritis|Juvenile chronic polyarthritis
C0837691|T047|AB|714.30|ICD9CM|Juv rheum arthritis NOS|Juv rheum arthritis NOS
C0837691|T047|PT|714.30|ICD9CM|Polyarticular juvenile rheumatoid arthritis, chronic or unspecified|Polyarticular juvenile rheumatoid arthritis, chronic or unspecified
C0157916|T047|AB|714.31|ICD9CM|Polyart juv rheum arthr|Polyart juv rheum arthr
C0157916|T047|PT|714.31|ICD9CM|Polyarticular juvenile rheumatoid arthritis, acute|Polyarticular juvenile rheumatoid arthritis, acute
C0157917|T047|AB|714.32|ICD9CM|Pauciart juv rheum arthr|Pauciart juv rheum arthr
C0157917|T047|PT|714.32|ICD9CM|Pauciarticular juvenile rheumatoid arthritis|Pauciarticular juvenile rheumatoid arthritis
C0157918|T047|AB|714.33|ICD9CM|Monoart juv rheum arthr|Monoart juv rheum arthr
C0157918|T047|PT|714.33|ICD9CM|Monoarticular juvenile rheumatoid arthritis|Monoarticular juvenile rheumatoid arthritis
C0152084|T047|AB|714.4|ICD9CM|Chr postrheum arthritis|Chr postrheum arthritis
C0152084|T047|PT|714.4|ICD9CM|Chronic postrheumatic arthropathy|Chronic postrheumatic arthropathy
C0157919|T047|HT|714.8|ICD9CM|Other specified inflammatory polyarthropathies|Other specified inflammatory polyarthropathies
C0994344|T047|AB|714.81|ICD9CM|Rheumatoid lung|Rheumatoid lung
C0994344|T047|PT|714.81|ICD9CM|Rheumatoid lung|Rheumatoid lung
C0157919|T047|AB|714.89|ICD9CM|Inflamm polyarthrop NEC|Inflamm polyarthrop NEC
C0157919|T047|PT|714.89|ICD9CM|Other specified inflammatory polyarthropathies|Other specified inflammatory polyarthropathies
C0162323|T047|AB|714.9|ICD9CM|Inflamm polyarthrop NOS|Inflamm polyarthrop NOS
C0162323|T047|PT|714.9|ICD9CM|Unspecified inflammatory polyarthropathy|Unspecified inflammatory polyarthropathy
C0263742|T047|HT|715|ICD9CM|Osteoarthrosis and allied disorders|Osteoarthrosis and allied disorders
C1384584|T047|HT|715.0|ICD9CM|Osteoarthrosis, generalized|Osteoarthrosis, generalized
C0157923|T047|AB|715.00|ICD9CM|General osteoarthrosis|General osteoarthrosis
C0157923|T047|PT|715.00|ICD9CM|Osteoarthrosis, generalized, site unspecified|Osteoarthrosis, generalized, site unspecified
C0157924|T047|AB|715.04|ICD9CM|Gen osteoarthros-hand|Gen osteoarthros-hand
C0157924|T047|PT|715.04|ICD9CM|Osteoarthrosis, generalized, hand|Osteoarthrosis, generalized, hand
C1384584|T047|AB|715.09|ICD9CM|General osteoarthrosis|General osteoarthrosis
C1384584|T047|PT|715.09|ICD9CM|Osteoarthrosis, generalized, multiple sites|Osteoarthrosis, generalized, multiple sites
C0157926|T047|HT|715.1|ICD9CM|Osteoarthrosis, localized, primary|Osteoarthrosis, localized, primary
C0157926|T047|AB|715.10|ICD9CM|Loc prim osteoart-unspec|Loc prim osteoart-unspec
C0157926|T047|PT|715.10|ICD9CM|Osteoarthrosis, localized, primary, site unspecified|Osteoarthrosis, localized, primary, site unspecified
C0263752|T047|AB|715.11|ICD9CM|Loc prim osteoart-shlder|Loc prim osteoart-shlder
C0263752|T047|PT|715.11|ICD9CM|Osteoarthrosis, localized, primary, shoulder region|Osteoarthrosis, localized, primary, shoulder region
C0263753|T047|AB|715.12|ICD9CM|Loc prim osteoart-up/arm|Loc prim osteoart-up/arm
C0263753|T047|PT|715.12|ICD9CM|Osteoarthrosis, localized, primary, upper arm|Osteoarthrosis, localized, primary, upper arm
C0263754|T047|AB|715.13|ICD9CM|Loc prim osteoart-forarm|Loc prim osteoart-forarm
C0263754|T047|PT|715.13|ICD9CM|Osteoarthrosis, localized, primary, forearm|Osteoarthrosis, localized, primary, forearm
C0263755|T047|AB|715.14|ICD9CM|Loc prim osteoarth-hand|Loc prim osteoarth-hand
C0263755|T047|PT|715.14|ICD9CM|Osteoarthrosis, localized, primary, hand|Osteoarthrosis, localized, primary, hand
C0473748|T047|AB|715.15|ICD9CM|Loc prim osteoart-pelvis|Loc prim osteoart-pelvis
C0473748|T047|PT|715.15|ICD9CM|Osteoarthrosis, localized, primary, pelvic region and thigh|Osteoarthrosis, localized, primary, pelvic region and thigh
C0263758|T047|AB|715.16|ICD9CM|Loc prim osteoart-l/leg|Loc prim osteoart-l/leg
C0263758|T047|PT|715.16|ICD9CM|Osteoarthrosis, localized, primary, lower leg|Osteoarthrosis, localized, primary, lower leg
C0263759|T047|AB|715.17|ICD9CM|Loc prim osteoarth-ankle|Loc prim osteoarth-ankle
C0263759|T047|PT|715.17|ICD9CM|Osteoarthrosis, localized, primary, ankle and foot|Osteoarthrosis, localized, primary, ankle and foot
C0701814|T047|AB|715.18|ICD9CM|Loc prim osteoarthr NEC|Loc prim osteoarthr NEC
C0701814|T047|PT|715.18|ICD9CM|Osteoarthrosis, localized, primary, other specified sites|Osteoarthrosis, localized, primary, other specified sites
C0473754|T047|HT|715.2|ICD9CM|Osteoarthrosis, localized, secondary|Osteoarthrosis, localized, secondary
C0157937|T047|AB|715.20|ICD9CM|Loc 2nd osteoarth-unspec|Loc 2nd osteoarth-unspec
C0157937|T047|PT|715.20|ICD9CM|Osteoarthrosis, localized, secondary, site unspecified|Osteoarthrosis, localized, secondary, site unspecified
C0157938|T047|AB|715.21|ICD9CM|Loc 2nd osteoarth-shlder|Loc 2nd osteoarth-shlder
C0157938|T047|PT|715.21|ICD9CM|Osteoarthrosis, localized, secondary, shoulder region|Osteoarthrosis, localized, secondary, shoulder region
C0157939|T047|AB|715.22|ICD9CM|Loc 2nd osteoarth-up/arm|Loc 2nd osteoarth-up/arm
C0157939|T047|PT|715.22|ICD9CM|Osteoarthrosis, localized, secondary, upper arm|Osteoarthrosis, localized, secondary, upper arm
C0157940|T047|AB|715.23|ICD9CM|Loc 2nd osteoart-forearm|Loc 2nd osteoart-forearm
C0157940|T047|PT|715.23|ICD9CM|Osteoarthrosis, localized, secondary, forearm|Osteoarthrosis, localized, secondary, forearm
C0157941|T047|AB|715.24|ICD9CM|Loc 2nd osteoarthro-hand|Loc 2nd osteoarthro-hand
C0157941|T047|PT|715.24|ICD9CM|Osteoarthrosis, localized, secondary, hand|Osteoarthrosis, localized, secondary, hand
C0157942|T047|AB|715.25|ICD9CM|Loc 2nd osteoarth-pelvis|Loc 2nd osteoarth-pelvis
C0157942|T047|PT|715.25|ICD9CM|Osteoarthrosis, localized, secondary, pelvic region and thigh|Osteoarthrosis, localized, secondary, pelvic region and thigh
C0157943|T047|AB|715.26|ICD9CM|Loc 2nd osteoarthr-l/leg|Loc 2nd osteoarthr-l/leg
C0157943|T047|PT|715.26|ICD9CM|Osteoarthrosis, localized, secondary, lower leg|Osteoarthrosis, localized, secondary, lower leg
C0157944|T047|AB|715.27|ICD9CM|Loc 2nd osteoarthr-ankle|Loc 2nd osteoarthr-ankle
C0157944|T047|PT|715.27|ICD9CM|Osteoarthrosis, localized, secondary, ankle and foot|Osteoarthrosis, localized, secondary, ankle and foot
C0157945|T047|AB|715.28|ICD9CM|Loc 2nd osteoarthros NEC|Loc 2nd osteoarthros NEC
C0157945|T047|PT|715.28|ICD9CM|Osteoarthrosis, localized, secondary, other specified sites|Osteoarthrosis, localized, secondary, other specified sites
C0157946|T047|HT|715.3|ICD9CM|Osteoarthrosis, localized, not specified whether primary or secondary|Osteoarthrosis, localized, not specified whether primary or secondary
C0157947|T047|AB|715.30|ICD9CM|Loc osteoarth NOS-unspec|Loc osteoarth NOS-unspec
C0157947|T047|PT|715.30|ICD9CM|Osteoarthrosis, localized, not specified whether primary or secondary, site unspecified|Osteoarthrosis, localized, not specified whether primary or secondary, site unspecified
C0157948|T047|AB|715.31|ICD9CM|Loc osteoarth NOS-shlder|Loc osteoarth NOS-shlder
C0157948|T047|PT|715.31|ICD9CM|Osteoarthrosis, localized, not specified whether primary or secondary, shoulder region|Osteoarthrosis, localized, not specified whether primary or secondary, shoulder region
C0157949|T047|AB|715.32|ICD9CM|Loc osteoarth NOS-up/arm|Loc osteoarth NOS-up/arm
C0157949|T047|PT|715.32|ICD9CM|Osteoarthrosis, localized, not specified whether primary or secondary, upper arm|Osteoarthrosis, localized, not specified whether primary or secondary, upper arm
C0157950|T047|AB|715.33|ICD9CM|Loc osteoart NOS-forearm|Loc osteoart NOS-forearm
C0157950|T047|PT|715.33|ICD9CM|Osteoarthrosis, localized, not specified whether primary or secondary, forearm|Osteoarthrosis, localized, not specified whether primary or secondary, forearm
C0157951|T047|AB|715.34|ICD9CM|Loc osteoarth NOS-hand|Loc osteoarth NOS-hand
C0157951|T047|PT|715.34|ICD9CM|Osteoarthrosis, localized, not specified whether primary or secondary, hand|Osteoarthrosis, localized, not specified whether primary or secondary, hand
C0157952|T047|AB|715.35|ICD9CM|Loc osteoarth NOS-pelvis|Loc osteoarth NOS-pelvis
C0157952|T047|PT|715.35|ICD9CM|Osteoarthrosis, localized, not specified whether primary or secondary, pelvic region and thigh|Osteoarthrosis, localized, not specified whether primary or secondary, pelvic region and thigh
C0157953|T047|AB|715.36|ICD9CM|Loc osteoarth NOS-l/leg|Loc osteoarth NOS-l/leg
C0157953|T047|PT|715.36|ICD9CM|Osteoarthrosis, localized, not specified whether primary or secondary, lower leg|Osteoarthrosis, localized, not specified whether primary or secondary, lower leg
C0157954|T047|AB|715.37|ICD9CM|Loc osteoarth NOS-ankle|Loc osteoarth NOS-ankle
C0157954|T047|PT|715.37|ICD9CM|Osteoarthrosis, localized, not specified whether primary or secondary, ankle and foot|Osteoarthrosis, localized, not specified whether primary or secondary, ankle and foot
C0157955|T047|AB|715.38|ICD9CM|Loc osteoar NOS-site NEC|Loc osteoar NOS-site NEC
C0157955|T047|PT|715.38|ICD9CM|Osteoarthrosis, localized, not specified whether primary or secondary, other specified sites|Osteoarthrosis, localized, not specified whether primary or secondary, other specified sites
C0263774|T047|HT|715.8|ICD9CM|Osteoarthrosis involving or with mention of more than one site, but not specified as generalized|Osteoarthrosis involving or with mention of more than one site, but not specified as generalized
C0157957|T047|AB|715.80|ICD9CM|Osteoarthrosis-mult site|Osteoarthrosis-mult site
C0157958|T047|AB|715.89|ICD9CM|Osteoarthrosis-mult site|Osteoarthrosis-mult site
C0029408|T047|HT|715.9|ICD9CM|Osteoarthrosis, unspecified whether generalized or localized|Osteoarthrosis, unspecified whether generalized or localized
C0157959|T047|AB|715.90|ICD9CM|Osteoarthros NOS-unspec|Osteoarthros NOS-unspec
C0157959|T047|PT|715.90|ICD9CM|Osteoarthrosis, unspecified whether generalized or localized, site unspecified|Osteoarthrosis, unspecified whether generalized or localized, site unspecified
C0157960|T047|AB|715.91|ICD9CM|Osteoarthros NOS-shlder|Osteoarthros NOS-shlder
C0157960|T047|PT|715.91|ICD9CM|Osteoarthrosis, unspecified whether generalized or localized, shoulder region|Osteoarthrosis, unspecified whether generalized or localized, shoulder region
C0157961|T047|AB|715.92|ICD9CM|Osteoarthros NOS-up/arm|Osteoarthros NOS-up/arm
C0157961|T047|PT|715.92|ICD9CM|Osteoarthrosis, unspecified whether generalized or localized, upper arm|Osteoarthrosis, unspecified whether generalized or localized, upper arm
C0157962|T047|AB|715.93|ICD9CM|Osteoarthros NOS-forearm|Osteoarthros NOS-forearm
C0157962|T047|PT|715.93|ICD9CM|Osteoarthrosis, unspecified whether generalized or localized, forearm|Osteoarthrosis, unspecified whether generalized or localized, forearm
C0157963|T047|AB|715.94|ICD9CM|Osteoarthros NOS-hand|Osteoarthros NOS-hand
C0157963|T047|PT|715.94|ICD9CM|Osteoarthrosis, unspecified whether generalized or localized, hand|Osteoarthrosis, unspecified whether generalized or localized, hand
C0157964|T047|AB|715.95|ICD9CM|Osteoarthros NOS-pelvis|Osteoarthros NOS-pelvis
C0157964|T047|PT|715.95|ICD9CM|Osteoarthrosis, unspecified whether generalized or localized, pelvic region and thigh|Osteoarthrosis, unspecified whether generalized or localized, pelvic region and thigh
C0157965|T047|AB|715.96|ICD9CM|Osteoarthros NOS-l/leg|Osteoarthros NOS-l/leg
C0157965|T047|PT|715.96|ICD9CM|Osteoarthrosis, unspecified whether generalized or localized, lower leg|Osteoarthrosis, unspecified whether generalized or localized, lower leg
C0157966|T047|AB|715.97|ICD9CM|Osteoarthros NOS-ankle|Osteoarthros NOS-ankle
C0157966|T047|PT|715.97|ICD9CM|Osteoarthrosis, unspecified whether generalized or localized, ankle and foot|Osteoarthrosis, unspecified whether generalized or localized, ankle and foot
C0157967|T047|AB|715.98|ICD9CM|Osteoarthro NOS-oth site|Osteoarthro NOS-oth site
C0157967|T047|PT|715.98|ICD9CM|Osteoarthrosis, unspecified whether generalized or localized, other specified sites|Osteoarthrosis, unspecified whether generalized or localized, other specified sites
C1442831|T047|HT|716|ICD9CM|Other and unspecified arthropathies|Other and unspecified arthropathies
C2745963|T047|HT|716.0|ICD9CM|Kaschin-Beck disease|Kaschin-Beck disease
C2745963|T047|AB|716.00|ICD9CM|Kaschin-beck dis-unspec|Kaschin-beck dis-unspec
C2745963|T047|PT|716.00|ICD9CM|Kaschin-Beck disease, site unspecified|Kaschin-Beck disease, site unspecified
C0157969|T047|AB|716.01|ICD9CM|Kaschin-beck dis-shlder|Kaschin-beck dis-shlder
C0157969|T047|PT|716.01|ICD9CM|Kaschin-Beck disease, shoulder region|Kaschin-Beck disease, shoulder region
C0157970|T047|AB|716.02|ICD9CM|Kaschin-beck dis-up/arm|Kaschin-beck dis-up/arm
C0157970|T047|PT|716.02|ICD9CM|Kaschin-Beck disease, upper arm|Kaschin-Beck disease, upper arm
C0157971|T047|AB|716.03|ICD9CM|Kaschin-beck dis-forearm|Kaschin-beck dis-forearm
C0157971|T047|PT|716.03|ICD9CM|Kaschin-Beck disease, forearm|Kaschin-Beck disease, forearm
C0157972|T047|AB|716.04|ICD9CM|Kaschin-beck dis-hand|Kaschin-beck dis-hand
C0157972|T047|PT|716.04|ICD9CM|Kaschin-Beck disease, hand|Kaschin-Beck disease, hand
C0409970|T047|AB|716.05|ICD9CM|Kaschin-beck dis-pelvis|Kaschin-beck dis-pelvis
C0409970|T047|PT|716.05|ICD9CM|Kaschin-Beck disease, pelvic region and thigh|Kaschin-Beck disease, pelvic region and thigh
C0157974|T047|AB|716.06|ICD9CM|Kaschin-beck dis-l/leg|Kaschin-beck dis-l/leg
C0157974|T047|PT|716.06|ICD9CM|Kaschin-Beck disease, lower leg|Kaschin-Beck disease, lower leg
C0409969|T047|AB|716.07|ICD9CM|Kaschin-beck dis-ankle|Kaschin-beck dis-ankle
C0409969|T047|PT|716.07|ICD9CM|Kaschin-Beck disease, ankle and foot|Kaschin-Beck disease, ankle and foot
C0409968|T047|AB|716.08|ICD9CM|Kaschin-beck dis NEC|Kaschin-beck dis NEC
C0409968|T047|PT|716.08|ICD9CM|Kaschin-Beck disease, other specified sites|Kaschin-Beck disease, other specified sites
C0157977|T047|AB|716.09|ICD9CM|Kaschin-beck dis-mult|Kaschin-beck dis-mult
C0157977|T047|PT|716.09|ICD9CM|Kaschin-Beck disease, multiple sites|Kaschin-Beck disease, multiple sites
C0152086|T037|HT|716.1|ICD9CM|Traumatic arthropathy|Traumatic arthropathy
C0152086|T037|AB|716.10|ICD9CM|Traum arthropathy-unspec|Traum arthropathy-unspec
C0152086|T037|PT|716.10|ICD9CM|Traumatic arthropathy, site unspecified|Traumatic arthropathy, site unspecified
C0409760|T037|AB|716.11|ICD9CM|Traum arthropathy-shlder|Traum arthropathy-shlder
C0409760|T037|PT|716.11|ICD9CM|Traumatic arthropathy, shoulder region|Traumatic arthropathy, shoulder region
C0409759|T037|AB|716.12|ICD9CM|Traum arthropathy-up/arm|Traum arthropathy-up/arm
C0409759|T037|PT|716.12|ICD9CM|Traumatic arthropathy, upper arm|Traumatic arthropathy, upper arm
C0409758|T037|AB|716.13|ICD9CM|Traum arthropath-forearm|Traum arthropath-forearm
C0409758|T037|PT|716.13|ICD9CM|Traumatic arthropathy, forearm|Traumatic arthropathy, forearm
C0409757|T037|AB|716.14|ICD9CM|Traum arthropathy-hand|Traum arthropathy-hand
C0409757|T037|PT|716.14|ICD9CM|Traumatic arthropathy, hand|Traumatic arthropathy, hand
C0409756|T047|AB|716.15|ICD9CM|Traum arthropathy-pelvis|Traum arthropathy-pelvis
C0409756|T047|PT|716.15|ICD9CM|Traumatic arthropathy, pelvic region and thigh|Traumatic arthropathy, pelvic region and thigh
C0409755|T037|AB|716.16|ICD9CM|Traum arthropathy-l/leg|Traum arthropathy-l/leg
C0409755|T037|PT|716.16|ICD9CM|Traumatic arthropathy, lower leg|Traumatic arthropathy, lower leg
C0409754|T037|AB|716.17|ICD9CM|Traum arthropathy-ankle|Traum arthropathy-ankle
C0409754|T037|PT|716.17|ICD9CM|Traumatic arthropathy, ankle and foot|Traumatic arthropathy, ankle and foot
C0409753|T037|AB|716.18|ICD9CM|Traum arthropathy NEC|Traum arthropathy NEC
C0409753|T037|PT|716.18|ICD9CM|Traumatic arthropathy, other specified sites|Traumatic arthropathy, other specified sites
C0409752|T037|AB|716.19|ICD9CM|Traum arthropathy-mult|Traum arthropathy-mult
C0409752|T037|PT|716.19|ICD9CM|Traumatic arthropathy, multiple sites|Traumatic arthropathy, multiple sites
C0157987|T047|HT|716.2|ICD9CM|Allergic arthritis|Allergic arthritis
C0157987|T047|AB|716.20|ICD9CM|Allerg arthritis-unspec|Allerg arthritis-unspec
C0157987|T047|PT|716.20|ICD9CM|Allergic arthritis, site unspecified|Allergic arthritis, site unspecified
C0409260|T047|AB|716.21|ICD9CM|Allerg arthritis-shlder|Allerg arthritis-shlder
C0409260|T047|PT|716.21|ICD9CM|Allergic arthritis, shoulder region|Allergic arthritis, shoulder region
C0409259|T047|AB|716.22|ICD9CM|Allerg arthritis-up/arm|Allerg arthritis-up/arm
C0409259|T047|PT|716.22|ICD9CM|Allergic arthritis, upper arm|Allergic arthritis, upper arm
C0409258|T047|AB|716.23|ICD9CM|Allerg arthritis-forearm|Allerg arthritis-forearm
C0409258|T047|PT|716.23|ICD9CM|Allergic arthritis, forearm|Allergic arthritis, forearm
C0409257|T047|AB|716.24|ICD9CM|Allerg arthritis-hand|Allerg arthritis-hand
C0409257|T047|PT|716.24|ICD9CM|Allergic arthritis, hand|Allergic arthritis, hand
C0409256|T047|AB|716.25|ICD9CM|Allerg arthritis-pelvis|Allerg arthritis-pelvis
C0409256|T047|PT|716.25|ICD9CM|Allergic arthritis, pelvic region and thigh|Allergic arthritis, pelvic region and thigh
C0409255|T047|AB|716.26|ICD9CM|Allerg arthritis-l/leg|Allerg arthritis-l/leg
C0409255|T047|PT|716.26|ICD9CM|Allergic arthritis, lower leg|Allergic arthritis, lower leg
C0409254|T047|AB|716.27|ICD9CM|Allerg arthritis-ankle|Allerg arthritis-ankle
C0409254|T047|PT|716.27|ICD9CM|Allergic arthritis, ankle and foot|Allergic arthritis, ankle and foot
C0409253|T047|AB|716.28|ICD9CM|Allerg arthritis NEC|Allerg arthritis NEC
C0409253|T047|PT|716.28|ICD9CM|Allergic arthritis, other specified sites|Allergic arthritis, other specified sites
C0409252|T047|AB|716.29|ICD9CM|Allerg arthritis-mult|Allerg arthritis-mult
C0409252|T047|PT|716.29|ICD9CM|Allergic arthritis, multiple sites|Allergic arthritis, multiple sites
C0157997|T047|HT|716.3|ICD9CM|Climacteric arthritis|Climacteric arthritis
C0157997|T047|AB|716.30|ICD9CM|Climact arthritis-unspec|Climact arthritis-unspec
C0157997|T047|PT|716.30|ICD9CM|Climacteric arthritis, site unspecified|Climacteric arthritis, site unspecified
C0409251|T047|AB|716.31|ICD9CM|Climact arthritis-shlder|Climact arthritis-shlder
C0409251|T047|PT|716.31|ICD9CM|Climacteric arthritis, shoulder region|Climacteric arthritis, shoulder region
C0409250|T047|AB|716.32|ICD9CM|Climact arthritis-up/arm|Climact arthritis-up/arm
C0409250|T047|PT|716.32|ICD9CM|Climacteric arthritis, upper arm|Climacteric arthritis, upper arm
C0409249|T047|AB|716.33|ICD9CM|Climact arthrit-forearm|Climact arthrit-forearm
C0409249|T047|PT|716.33|ICD9CM|Climacteric arthritis, forearm|Climacteric arthritis, forearm
C0409248|T047|AB|716.34|ICD9CM|Climact arthritis-hand|Climact arthritis-hand
C0409248|T047|PT|716.34|ICD9CM|Climacteric arthritis, hand|Climacteric arthritis, hand
C0409247|T047|AB|716.35|ICD9CM|Climact arthritis-pelvis|Climact arthritis-pelvis
C0409247|T047|PT|716.35|ICD9CM|Climacteric arthritis, pelvic region and thigh|Climacteric arthritis, pelvic region and thigh
C0409246|T047|AB|716.36|ICD9CM|Climact arthritis-l/leg|Climact arthritis-l/leg
C0409246|T047|PT|716.36|ICD9CM|Climacteric arthritis, lower leg|Climacteric arthritis, lower leg
C0158004|T047|AB|716.37|ICD9CM|Climact arthritis-ankle|Climact arthritis-ankle
C0158004|T047|PT|716.37|ICD9CM|Climacteric arthritis, ankle and foot|Climacteric arthritis, ankle and foot
C0409244|T047|AB|716.38|ICD9CM|Climact arthritis NEC|Climact arthritis NEC
C0409244|T047|PT|716.38|ICD9CM|Climacteric arthritis, other specified sites|Climacteric arthritis, other specified sites
C0409243|T047|AB|716.39|ICD9CM|Climact arthritis-mult|Climact arthritis-mult
C0409243|T047|PT|716.39|ICD9CM|Climacteric arthritis, multiple sites|Climacteric arthritis, multiple sites
C0152083|T047|HT|716.4|ICD9CM|Transient arthropathy|Transient arthropathy
C0152083|T047|AB|716.40|ICD9CM|Trans arthropathy-unspec|Trans arthropathy-unspec
C0152083|T047|PT|716.40|ICD9CM|Transient arthropathy, site unspecified|Transient arthropathy, site unspecified
C0158007|T047|AB|716.41|ICD9CM|Trans arthropathy-shlder|Trans arthropathy-shlder
C0158007|T047|PT|716.41|ICD9CM|Transient arthropathy, shoulder region|Transient arthropathy, shoulder region
C0409816|T047|AB|716.42|ICD9CM|Trans arthropathy-up/arm|Trans arthropathy-up/arm
C0409816|T047|PT|716.42|ICD9CM|Transient arthropathy, upper arm|Transient arthropathy, upper arm
C0409815|T047|AB|716.43|ICD9CM|Trans arthropath-forearm|Trans arthropath-forearm
C0409815|T047|PT|716.43|ICD9CM|Transient arthropathy, forearm|Transient arthropathy, forearm
C0409814|T047|AB|716.44|ICD9CM|Trans arthropathy-hand|Trans arthropathy-hand
C0409814|T047|PT|716.44|ICD9CM|Transient arthropathy, hand|Transient arthropathy, hand
C0409813|T047|AB|716.45|ICD9CM|Trans arthropathy-pelvis|Trans arthropathy-pelvis
C0409813|T047|PT|716.45|ICD9CM|Transient arthropathy, pelvic region and thigh|Transient arthropathy, pelvic region and thigh
C0409812|T047|AB|716.46|ICD9CM|Trans arthropathy-l/leg|Trans arthropathy-l/leg
C0409812|T047|PT|716.46|ICD9CM|Transient arthropathy, lower leg|Transient arthropathy, lower leg
C0409811|T047|AB|716.47|ICD9CM|Trans arthropathy-ankle|Trans arthropathy-ankle
C0409811|T047|PT|716.47|ICD9CM|Transient arthropathy, ankle and foot|Transient arthropathy, ankle and foot
C0409810|T047|AB|716.48|ICD9CM|Trans arthropathy NEC|Trans arthropathy NEC
C0409810|T047|PT|716.48|ICD9CM|Transient arthropathy, other specified sites|Transient arthropathy, other specified sites
C0409809|T047|AB|716.49|ICD9CM|Trans arthropathy-mult|Trans arthropathy-mult
C0409809|T047|PT|716.49|ICD9CM|Transient arthropathy, multiple sites|Transient arthropathy, multiple sites
C1692323|T047|HT|716.5|ICD9CM|Unspecified polyarthropathy or polyarthritis|Unspecified polyarthropathy or polyarthritis
C1692323|T047|AB|716.50|ICD9CM|Polyarthritis NOS-unspec|Polyarthritis NOS-unspec
C1692323|T047|PT|716.50|ICD9CM|Unspecified polyarthropathy or polyarthritis, site unspecified|Unspecified polyarthropathy or polyarthritis, site unspecified
C0158017|T047|AB|716.51|ICD9CM|Polyarthritis NOS-shlder|Polyarthritis NOS-shlder
C0158017|T047|PT|716.51|ICD9CM|Unspecified polyarthropathy or polyarthritis, shoulder region|Unspecified polyarthropathy or polyarthritis, shoulder region
C0158018|T047|AB|716.52|ICD9CM|Polyarthritis NOS-up/arm|Polyarthritis NOS-up/arm
C0158018|T047|PT|716.52|ICD9CM|Unspecified polyarthropathy or polyarthritis, upper arm|Unspecified polyarthropathy or polyarthritis, upper arm
C0158019|T047|AB|716.53|ICD9CM|Polyarthrit NOS-forearm|Polyarthrit NOS-forearm
C0158019|T047|PT|716.53|ICD9CM|Unspecified polyarthropathy or polyarthritis, forearm|Unspecified polyarthropathy or polyarthritis, forearm
C0158020|T047|AB|716.54|ICD9CM|Polyarthritis NOS-hand|Polyarthritis NOS-hand
C0158020|T047|PT|716.54|ICD9CM|Unspecified polyarthropathy or polyarthritis, hand|Unspecified polyarthropathy or polyarthritis, hand
C0158021|T047|AB|716.55|ICD9CM|Polyarthritis NOS-pelvis|Polyarthritis NOS-pelvis
C0158021|T047|PT|716.55|ICD9CM|Unspecified polyarthropathy or polyarthritis, pelvic region and thigh|Unspecified polyarthropathy or polyarthritis, pelvic region and thigh
C0158022|T047|AB|716.56|ICD9CM|Polyarthritis NOS-l/leg|Polyarthritis NOS-l/leg
C0158022|T047|PT|716.56|ICD9CM|Unspecified polyarthropathy or polyarthritis, lower leg|Unspecified polyarthropathy or polyarthritis, lower leg
C0158023|T047|AB|716.57|ICD9CM|Polyarthritis NOS-ankle|Polyarthritis NOS-ankle
C0158023|T047|PT|716.57|ICD9CM|Unspecified polyarthropathy or polyarthritis, ankle and foot|Unspecified polyarthropathy or polyarthritis, ankle and foot
C0158024|T047|AB|716.58|ICD9CM|Polyarthrit NOS-oth site|Polyarthrit NOS-oth site
C0158024|T047|PT|716.58|ICD9CM|Unspecified polyarthropathy or polyarthritis, other specified sites|Unspecified polyarthropathy or polyarthritis, other specified sites
C0546840|T047|AB|716.59|ICD9CM|Polyarthritis NOS-mult|Polyarthritis NOS-mult
C0546840|T047|PT|716.59|ICD9CM|Unspecified polyarthropathy or polyarthritis, multiple sites|Unspecified polyarthropathy or polyarthritis, multiple sites
C0158026|T047|HT|716.6|ICD9CM|Unspecified monoarthritis|Unspecified monoarthritis
C0158026|T047|AB|716.60|ICD9CM|Monoarthritis NOS-unspec|Monoarthritis NOS-unspec
C0158026|T047|PT|716.60|ICD9CM|Unspecified monoarthritis, site unspecified|Unspecified monoarthritis, site unspecified
C0409232|T047|AB|716.61|ICD9CM|Monoarthritis NOS-shlder|Monoarthritis NOS-shlder
C0409232|T047|PT|716.61|ICD9CM|Unspecified monoarthritis, shoulder region|Unspecified monoarthritis, shoulder region
C0409231|T047|AB|716.62|ICD9CM|Monoarthritis NOS-up/arm|Monoarthritis NOS-up/arm
C0409231|T047|PT|716.62|ICD9CM|Unspecified monoarthritis, upper arm|Unspecified monoarthritis, upper arm
C0409230|T047|AB|716.63|ICD9CM|Monoarthrit NOS-forearm|Monoarthrit NOS-forearm
C0409230|T047|PT|716.63|ICD9CM|Unspecified monoarthritis, forearm|Unspecified monoarthritis, forearm
C0409229|T047|AB|716.64|ICD9CM|Monoarthritis NOS-hand|Monoarthritis NOS-hand
C0409229|T047|PT|716.64|ICD9CM|Unspecified monoarthritis, hand|Unspecified monoarthritis, hand
C0409228|T047|AB|716.65|ICD9CM|Monoarthritis NOS-pelvis|Monoarthritis NOS-pelvis
C0409228|T047|PT|716.65|ICD9CM|Unspecified monoarthritis, pelvic region and thigh|Unspecified monoarthritis, pelvic region and thigh
C0409227|T047|AB|716.66|ICD9CM|Monoarthritis NOS-l/leg|Monoarthritis NOS-l/leg
C0409227|T047|PT|716.66|ICD9CM|Unspecified monoarthritis, lower leg|Unspecified monoarthritis, lower leg
C0409226|T047|AB|716.67|ICD9CM|Monoarthritis NOS-ankle|Monoarthritis NOS-ankle
C0409226|T047|PT|716.67|ICD9CM|Unspecified monoarthritis, ankle and foot|Unspecified monoarthritis, ankle and foot
C0409225|T047|AB|716.68|ICD9CM|Monoarthrit NOS-oth site|Monoarthrit NOS-oth site
C0409225|T047|PT|716.68|ICD9CM|Unspecified monoarthritis, other specified sites|Unspecified monoarthritis, other specified sites
C0029746|T047|HT|716.8|ICD9CM|Other specified arthropathy|Other specified arthropathy
C0869062|T047|AB|716.80|ICD9CM|Arthropathy NEC-unspec|Arthropathy NEC-unspec
C0869062|T047|PT|716.80|ICD9CM|Other specified arthropathy, site unspecified|Other specified arthropathy, site unspecified
C0409223|T047|AB|716.81|ICD9CM|Arthropathy NEC-shlder|Arthropathy NEC-shlder
C0409223|T047|PT|716.81|ICD9CM|Other specified arthropathy, shoulder region|Other specified arthropathy, shoulder region
C0409222|T047|AB|716.82|ICD9CM|Arthropathy NEC-up/arm|Arthropathy NEC-up/arm
C0409222|T047|PT|716.82|ICD9CM|Other specified arthropathy, upper arm|Other specified arthropathy, upper arm
C0409221|T047|AB|716.83|ICD9CM|Arthropathy NEC-forearm|Arthropathy NEC-forearm
C0409221|T047|PT|716.83|ICD9CM|Other specified arthropathy, forearm|Other specified arthropathy, forearm
C0409220|T047|AB|716.84|ICD9CM|Arthropathy NEC-hand|Arthropathy NEC-hand
C0409220|T047|PT|716.84|ICD9CM|Other specified arthropathy, hand|Other specified arthropathy, hand
C0409219|T047|AB|716.85|ICD9CM|Arthropathy NEC-pelvis|Arthropathy NEC-pelvis
C0409219|T047|PT|716.85|ICD9CM|Other specified arthropathy, pelvic region and thigh|Other specified arthropathy, pelvic region and thigh
C0409218|T047|AB|716.86|ICD9CM|Arthropathy NEC-l/leg|Arthropathy NEC-l/leg
C0409218|T047|PT|716.86|ICD9CM|Other specified arthropathy, lower leg|Other specified arthropathy, lower leg
C0409217|T047|AB|716.87|ICD9CM|Arthropathy NEC-ankle|Arthropathy NEC-ankle
C0409217|T047|PT|716.87|ICD9CM|Other specified arthropathy, ankle and foot|Other specified arthropathy, ankle and foot
C0409216|T047|AB|716.88|ICD9CM|Arthropathy NEC-oth site|Arthropathy NEC-oth site
C0409216|T047|PT|716.88|ICD9CM|Other specified arthropathy, other specified sites|Other specified arthropathy, other specified sites
C0409215|T047|AB|716.89|ICD9CM|Arthropathy NEC-mult|Arthropathy NEC-mult
C0409215|T047|PT|716.89|ICD9CM|Other specified arthropathy, multiple sites|Other specified arthropathy, multiple sites
C0022408|T047|HT|716.9|ICD9CM|Arthropathy, unspecified|Arthropathy, unspecified
C0022408|T047|AB|716.90|ICD9CM|Arthropathy NOS-unspec|Arthropathy NOS-unspec
C0022408|T047|PT|716.90|ICD9CM|Arthropathy, unspecified, site unspecified|Arthropathy, unspecified, site unspecified
C0158044|T047|AB|716.91|ICD9CM|Arthropathy NOS-shlder|Arthropathy NOS-shlder
C0158044|T047|PT|716.91|ICD9CM|Arthropathy, unspecified, shoulder region|Arthropathy, unspecified, shoulder region
C0158045|T047|AB|716.92|ICD9CM|Arthropathy NOS-up/arm|Arthropathy NOS-up/arm
C0158045|T047|PT|716.92|ICD9CM|Arthropathy, unspecified, upper arm|Arthropathy, unspecified, upper arm
C0409209|T047|AB|716.93|ICD9CM|Arthropathy NOS-forearm|Arthropathy NOS-forearm
C0409209|T047|PT|716.93|ICD9CM|Arthropathy, unspecified, forearm|Arthropathy, unspecified, forearm
C0158234|T047|AB|716.94|ICD9CM|Arthropathy NOS-hand|Arthropathy NOS-hand
C0158234|T047|PT|716.94|ICD9CM|Arthropathy, unspecified, hand|Arthropathy, unspecified, hand
C0158048|T047|AB|716.95|ICD9CM|Arthropathy NOS-pelvis|Arthropathy NOS-pelvis
C0158048|T047|PT|716.95|ICD9CM|Arthropathy, unspecified, pelvic region and thigh|Arthropathy, unspecified, pelvic region and thigh
C0158049|T047|AB|716.96|ICD9CM|Arthropathy NOS-l/leg|Arthropathy NOS-l/leg
C0158049|T047|PT|716.96|ICD9CM|Arthropathy, unspecified, lower leg|Arthropathy, unspecified, lower leg
C0158050|T047|AB|716.97|ICD9CM|Arthropathy NOS-ankle|Arthropathy NOS-ankle
C0158050|T047|PT|716.97|ICD9CM|Arthropathy, unspecified, ankle and foot|Arthropathy, unspecified, ankle and foot
C0158051|T047|AB|716.98|ICD9CM|Arthropathy NOS-oth site|Arthropathy NOS-oth site
C0158051|T047|PT|716.98|ICD9CM|Arthropathy, unspecified, other specified sites|Arthropathy, unspecified, other specified sites
C0158052|T047|AB|716.99|ICD9CM|Arthropathy NOS-mult|Arthropathy NOS-mult
C0158052|T047|PT|716.99|ICD9CM|Arthropathy, unspecified, multiple sites|Arthropathy, unspecified, multiple sites
C0158053|T047|HT|717|ICD9CM|Internal derangement of knee|Internal derangement of knee
C0158054|T033|PT|717.0|ICD9CM|Old bucket handle tear of medial meniscus|Old bucket handle tear of medial meniscus
C0158054|T033|AB|717.0|ICD9CM|Old bucket tear med men|Old bucket tear med men
C0158055|T037|AB|717.1|ICD9CM|Derang ant med meniscus|Derang ant med meniscus
C0158055|T037|PT|717.1|ICD9CM|Derangement of anterior horn of medial meniscus|Derangement of anterior horn of medial meniscus
C0158056|T037|AB|717.2|ICD9CM|Derang post med meniscus|Derang post med meniscus
C0158056|T037|PT|717.2|ICD9CM|Derangement of posterior horn of medial meniscus|Derangement of posterior horn of medial meniscus
C0158057|T190|AB|717.3|ICD9CM|Derang med meniscus NEC|Derang med meniscus NEC
C0158057|T190|PT|717.3|ICD9CM|Other and unspecified derangement of medial meniscus|Other and unspecified derangement of medial meniscus
C0158058|T037|HT|717.4|ICD9CM|Derangement of lateral meniscus|Derangement of lateral meniscus
C0158058|T037|AB|717.40|ICD9CM|Derang lat meniscus NOS|Derang lat meniscus NOS
C0158058|T037|PT|717.40|ICD9CM|Derangement of lateral meniscus, unspecified|Derangement of lateral meniscus, unspecified
C0434992|T037|PT|717.41|ICD9CM|Bucket handle tear of lateral meniscus|Bucket handle tear of lateral meniscus
C0434992|T037|AB|717.41|ICD9CM|Old bucket tear lat men|Old bucket tear lat men
C0158060|T037|AB|717.42|ICD9CM|Derange ant lat meniscus|Derange ant lat meniscus
C0158060|T037|PT|717.42|ICD9CM|Derangement of anterior horn of lateral meniscus|Derangement of anterior horn of lateral meniscus
C0158061|T037|AB|717.43|ICD9CM|Derang post lat meniscus|Derang post lat meniscus
C0158061|T037|PT|717.43|ICD9CM|Derangement of posterior horn of lateral meniscus|Derangement of posterior horn of lateral meniscus
C0158062|T037|AB|717.49|ICD9CM|Derang lat meniscus NEC|Derang lat meniscus NEC
C0158062|T037|PT|717.49|ICD9CM|Other derangement of lateral meniscus|Other derangement of lateral meniscus
C0868743|T190|AB|717.5|ICD9CM|Derangement meniscus NEC|Derangement meniscus NEC
C0868743|T190|PT|717.5|ICD9CM|Derangement of meniscus, not elsewhere classified|Derangement of meniscus, not elsewhere classified
C0343161|T020|AB|717.6|ICD9CM|Loose body in knee|Loose body in knee
C0343161|T020|PT|717.6|ICD9CM|Loose body in knee|Loose body in knee
C0008475|T047|PT|717.7|ICD9CM|Chondromalacia of patella|Chondromalacia of patella
C0008475|T047|AB|717.7|ICD9CM|Chondromalacia patellae|Chondromalacia patellae
C0158065|T047|HT|717.8|ICD9CM|Other internal derangement of knee|Other internal derangement of knee
C0158066|T037|AB|717.81|ICD9CM|Old disrupt lat collat|Old disrupt lat collat
C0158066|T037|PT|717.81|ICD9CM|Old disruption of lateral collateral ligament|Old disruption of lateral collateral ligament
C0158067|T037|AB|717.82|ICD9CM|Old disrupt med collat|Old disrupt med collat
C0158067|T037|PT|717.82|ICD9CM|Old disruption of medial collateral ligament|Old disruption of medial collateral ligament
C0158068|T037|AB|717.83|ICD9CM|Old disrupt ant cruciate|Old disrupt ant cruciate
C0158068|T037|PT|717.83|ICD9CM|Old disruption of anterior cruciate ligament|Old disruption of anterior cruciate ligament
C0158069|T037|AB|717.84|ICD9CM|Old disrupt post cruciat|Old disrupt post cruciat
C0158069|T037|PT|717.84|ICD9CM|Old disruption of posterior cruciate ligament|Old disruption of posterior cruciate ligament
C0158070|T037|AB|717.85|ICD9CM|Old disrupt knee lig NEC|Old disrupt knee lig NEC
C0158070|T037|PT|717.85|ICD9CM|Old disruption of other ligaments of knee|Old disruption of other ligaments of knee
C0158065|T047|AB|717.89|ICD9CM|Int derangement knee NEC|Int derangement knee NEC
C0158065|T047|PT|717.89|ICD9CM|Other internal derangement of knee|Other internal derangement of knee
C0158053|T047|AB|717.9|ICD9CM|Int derangement knee NOS|Int derangement knee NOS
C0158053|T047|PT|717.9|ICD9CM|Unspecified internal derangement of knee|Unspecified internal derangement of knee
C0158072|T037|HT|718|ICD9CM|Other derangement of joint|Other derangement of joint
C0158073|T047|HT|718.0|ICD9CM|Articular cartilage disorder|Articular cartilage disorder
C0158073|T047|AB|718.00|ICD9CM|Artic cartil dis-unspec|Artic cartil dis-unspec
C0158073|T047|PT|718.00|ICD9CM|Articular cartilage disorder, site unspecified|Articular cartilage disorder, site unspecified
C0263793|T047|AB|718.01|ICD9CM|Artic cartil dis-shlder|Artic cartil dis-shlder
C0263793|T047|PT|718.01|ICD9CM|Articular cartilage disorder, shoulder region|Articular cartilage disorder, shoulder region
C0263794|T047|AB|718.02|ICD9CM|Artic cartil dis-up/arm|Artic cartil dis-up/arm
C0263794|T047|PT|718.02|ICD9CM|Articular cartilage disorder, upper arm|Articular cartilage disorder, upper arm
C0263795|T047|AB|718.03|ICD9CM|Artic cartil dis-forearm|Artic cartil dis-forearm
C0263795|T047|PT|718.03|ICD9CM|Articular cartilage disorder, forearm|Articular cartilage disorder, forearm
C0158077|T047|AB|718.04|ICD9CM|Artic cartil dis-hand|Artic cartil dis-hand
C0158077|T047|PT|718.04|ICD9CM|Articular cartilage disorder, hand|Articular cartilage disorder, hand
C0410332|T047|AB|718.05|ICD9CM|Artic cartil dis-pelvis|Artic cartil dis-pelvis
C0410332|T047|PT|718.05|ICD9CM|Articular cartilage disorder, pelvic region and thigh|Articular cartilage disorder, pelvic region and thigh
C0263799|T047|AB|718.07|ICD9CM|Artic cartil dis-ankle|Artic cartil dis-ankle
C0263799|T047|PT|718.07|ICD9CM|Articular cartilage disorder, ankle and foot|Articular cartilage disorder, ankle and foot
C0410331|T047|AB|718.08|ICD9CM|Artic cartil dis-jt NEC|Artic cartil dis-jt NEC
C0410331|T047|PT|718.08|ICD9CM|Articular cartilage disorder, other specified sites|Articular cartilage disorder, other specified sites
C0263801|T047|AB|718.09|ICD9CM|Artic cartil dis-mult jt|Artic cartil dis-mult jt
C0263801|T047|PT|718.09|ICD9CM|Articular cartilage disorder, multiple sites|Articular cartilage disorder, multiple sites
C0022411|T020|HT|718.1|ICD9CM|Loose body in joint|Loose body in joint
C0022411|T020|PT|718.10|ICD9CM|Loose body in joint, site unspecified|Loose body in joint, site unspecified
C0022411|T020|AB|718.10|ICD9CM|Loose body-unspec|Loose body-unspec
C0158082|T020|PT|718.11|ICD9CM|Loose body in joint, shoulder region|Loose body in joint, shoulder region
C0158082|T020|AB|718.11|ICD9CM|Loose body-shlder|Loose body-shlder
C0158083|T020|PT|718.12|ICD9CM|Loose body in joint, upper arm|Loose body in joint, upper arm
C0158083|T020|AB|718.12|ICD9CM|Loose body-up/arm|Loose body-up/arm
C0158084|T020|PT|718.13|ICD9CM|Loose body in joint, forearm|Loose body in joint, forearm
C0158084|T020|AB|718.13|ICD9CM|Loose body-forearm|Loose body-forearm
C0158085|T020|PT|718.14|ICD9CM|Loose body in joint, hand|Loose body in joint, hand
C0158085|T020|AB|718.14|ICD9CM|Loose body-hand|Loose body-hand
C0158086|T020|PT|718.15|ICD9CM|Loose body in joint, pelvic region and thigh|Loose body in joint, pelvic region and thigh
C0158086|T020|AB|718.15|ICD9CM|Loose body-pelvis|Loose body-pelvis
C0158087|T020|PT|718.17|ICD9CM|Loose body in joint, ankle and foot|Loose body in joint, ankle and foot
C0158087|T020|AB|718.17|ICD9CM|Loose body-ankle|Loose body-ankle
C0023988|T020|PT|718.18|ICD9CM|Loose body in joint, other specified sites|Loose body in joint, other specified sites
C0023988|T020|AB|718.18|ICD9CM|Loose body-joint NEC|Loose body-joint NEC
C0158088|T020|PT|718.19|ICD9CM|Loose body in joint, multiple sites|Loose body in joint, multiple sites
C0158088|T020|AB|718.19|ICD9CM|Loose body-mult joints|Loose body-mult joints
C0158090|T046|HT|718.2|ICD9CM|Pathological dislocation|Pathological dislocation
C0158090|T046|AB|718.20|ICD9CM|Pathol dislocat-unspec|Pathol dislocat-unspec
C0158090|T046|PT|718.20|ICD9CM|Pathological dislocation of joint, site unspecified|Pathological dislocation of joint, site unspecified
C0158091|T020|AB|718.21|ICD9CM|Pathol dislocat-shlder|Pathol dislocat-shlder
C0158091|T020|PT|718.21|ICD9CM|Pathological dislocation of joint, shoulder region|Pathological dislocation of joint, shoulder region
C0263805|T047|AB|718.22|ICD9CM|Pathol dislocat-up/arm|Pathol dislocat-up/arm
C0263805|T047|PT|718.22|ICD9CM|Pathological dislocation of joint, upper arm|Pathological dislocation of joint, upper arm
C0263806|T047|AB|718.23|ICD9CM|Pathol dislocat-forearm|Pathol dislocat-forearm
C0263806|T047|PT|718.23|ICD9CM|Pathological dislocation of joint, forearm|Pathological dislocation of joint, forearm
C0158094|T046|AB|718.24|ICD9CM|Pathol dislocat-hand|Pathol dislocat-hand
C0158094|T046|PT|718.24|ICD9CM|Pathological dislocation of joint, hand|Pathological dislocation of joint, hand
C0158095|T047|AB|718.25|ICD9CM|Pathol dislocat-pelvis|Pathol dislocat-pelvis
C0158095|T047|PT|718.25|ICD9CM|Pathological dislocation of joint, pelvic region and thigh|Pathological dislocation of joint, pelvic region and thigh
C0263809|T047|AB|718.26|ICD9CM|Pathol dislocat-l/leg|Pathol dislocat-l/leg
C0263809|T047|PT|718.26|ICD9CM|Pathological dislocation of joint, lower leg|Pathological dislocation of joint, lower leg
C0263810|T046|AB|718.27|ICD9CM|Pathol dislocat-ankle|Pathol dislocat-ankle
C0263810|T046|PT|718.27|ICD9CM|Pathological dislocation of joint, ankle and foot|Pathological dislocation of joint, ankle and foot
C0158098|T047|AB|718.28|ICD9CM|Pathol dislocat-jt NEC|Pathol dislocat-jt NEC
C0158098|T047|PT|718.28|ICD9CM|Pathological dislocation of joint, other specified sites|Pathological dislocation of joint, other specified sites
C0263812|T046|AB|718.29|ICD9CM|Pathol dislocat-mult jts|Pathol dislocat-mult jts
C0263812|T046|PT|718.29|ICD9CM|Pathological dislocation of joint, multiple sites|Pathological dislocation of joint, multiple sites
C0158100|T037|HT|718.3|ICD9CM|Recurrent dislocation of joint|Recurrent dislocation of joint
C0158100|T037|AB|718.30|ICD9CM|Recur dislocat-unspec|Recur dislocat-unspec
C0158100|T037|PT|718.30|ICD9CM|Recurrent dislocation of joint, site unspecified|Recurrent dislocation of joint, site unspecified
C0409415|T037|AB|718.31|ICD9CM|Recur dislocat-shlder|Recur dislocat-shlder
C0409415|T037|PT|718.31|ICD9CM|Recurrent dislocation of joint, shoulder region|Recurrent dislocation of joint, shoulder region
C0263814|T037|AB|718.32|ICD9CM|Recur dislocat-up/arm|Recur dislocat-up/arm
C0263814|T037|PT|718.32|ICD9CM|Recurrent dislocation of joint, upper arm|Recurrent dislocation of joint, upper arm
C0263815|T037|AB|718.33|ICD9CM|Recur dislocat-forearm|Recur dislocat-forearm
C0263815|T037|PT|718.33|ICD9CM|Recurrent dislocation of joint, forearm|Recurrent dislocation of joint, forearm
C0263816|T037|AB|718.34|ICD9CM|Recur dislocat-hand|Recur dislocat-hand
C0263816|T037|PT|718.34|ICD9CM|Recurrent dislocation of joint, hand|Recurrent dislocation of joint, hand
C0158105|T046|AB|718.35|ICD9CM|Recur dislocat-pelvis|Recur dislocat-pelvis
C0158105|T046|PT|718.35|ICD9CM|Recurrent dislocation of joint, pelvic region and thigh|Recurrent dislocation of joint, pelvic region and thigh
C0263819|T037|AB|718.36|ICD9CM|Recur dislocat-l/leg|Recur dislocat-l/leg
C0263819|T037|PT|718.36|ICD9CM|Recurrent dislocation of joint, lower leg|Recurrent dislocation of joint, lower leg
C0263820|T046|AB|718.37|ICD9CM|Recur dislocat-ankle|Recur dislocat-ankle
C0263820|T046|PT|718.37|ICD9CM|Recurrent dislocation of joint, ankle and foot|Recurrent dislocation of joint, ankle and foot
C0158108|T037|AB|718.38|ICD9CM|Recur dislocat-jt NEC|Recur dislocat-jt NEC
C0158108|T037|PT|718.38|ICD9CM|Recurrent dislocation of joint, other specified sites|Recurrent dislocation of joint, other specified sites
C0263822|T037|AB|718.39|ICD9CM|Recur dislocat-mult jts|Recur dislocat-mult jts
C0263822|T037|PT|718.39|ICD9CM|Recurrent dislocation of joint, multiple sites|Recurrent dislocation of joint, multiple sites
C0009918|T190|HT|718.4|ICD9CM|Contracture of joint|Contracture of joint
C0009918|T190|PT|718.40|ICD9CM|Contracture of joint, site unspecified|Contracture of joint, site unspecified
C0009918|T190|AB|718.40|ICD9CM|Jt contracture-unspec|Jt contracture-unspec
C0158110|T020|PT|718.41|ICD9CM|Contracture of joint, shoulder region|Contracture of joint, shoulder region
C0158110|T020|AB|718.41|ICD9CM|Jt contracture-shlder|Jt contracture-shlder
C0158111|T020|PT|718.42|ICD9CM|Contracture of joint, upper arm|Contracture of joint, upper arm
C0158111|T020|AB|718.42|ICD9CM|Jt contracture-up/arm|Jt contracture-up/arm
C0158112|T190|PT|718.43|ICD9CM|Contracture of joint, forearm|Contracture of joint, forearm
C0158112|T190|AB|718.43|ICD9CM|Jt contracture-forearm|Jt contracture-forearm
C0158113|T190|PT|718.44|ICD9CM|Contracture of joint, hand|Contracture of joint, hand
C0158113|T190|AB|718.44|ICD9CM|Jt contracture-hand|Jt contracture-hand
C1306306|T047|PT|718.45|ICD9CM|Contracture of joint, pelvic region and thigh|Contracture of joint, pelvic region and thigh
C1306306|T047|AB|718.45|ICD9CM|Jt contracture-pelvis|Jt contracture-pelvis
C0158115|T020|PT|718.46|ICD9CM|Contracture of joint, lower leg|Contracture of joint, lower leg
C0158115|T020|AB|718.46|ICD9CM|Jt contracture-l/leg|Jt contracture-l/leg
C1963664|T020|PT|718.47|ICD9CM|Contracture of joint, ankle and foot|Contracture of joint, ankle and foot
C1963664|T020|AB|718.47|ICD9CM|Jt contracture-ankle|Jt contracture-ankle
C0158117|T020|PT|718.48|ICD9CM|Contracture of joint, other specified sites|Contracture of joint, other specified sites
C0158117|T020|AB|718.48|ICD9CM|Jt contracture-jt NEC|Jt contracture-jt NEC
C0158118|T020|PT|718.49|ICD9CM|Contracture of joint, multiple sites|Contracture of joint, multiple sites
C0158118|T020|AB|718.49|ICD9CM|Jt contracture-mult jts|Jt contracture-mult jts
C0003090|T046|HT|718.5|ICD9CM|Ankylosis of joint|Ankylosis of joint
C0003090|T046|PT|718.50|ICD9CM|Ankylosis of joint, site unspecified|Ankylosis of joint, site unspecified
C0003090|T046|AB|718.50|ICD9CM|Ankylosis-unspec|Ankylosis-unspec
C0158119|T020|PT|718.51|ICD9CM|Ankylosis of joint, shoulder region|Ankylosis of joint, shoulder region
C0158119|T020|AB|718.51|ICD9CM|Ankylosis-shoulder|Ankylosis-shoulder
C0158120|T020|PT|718.52|ICD9CM|Ankylosis of joint, upper arm|Ankylosis of joint, upper arm
C0158120|T020|AB|718.52|ICD9CM|Ankylosis-upper/arm|Ankylosis-upper/arm
C0158121|T020|PT|718.53|ICD9CM|Ankylosis of joint, forearm|Ankylosis of joint, forearm
C0158121|T020|AB|718.53|ICD9CM|Ankylosis-forearm|Ankylosis-forearm
C0158122|T020|PT|718.54|ICD9CM|Ankylosis of joint, hand|Ankylosis of joint, hand
C0158122|T020|AB|718.54|ICD9CM|Ankylosis-hand|Ankylosis-hand
C0158123|T047|PT|718.55|ICD9CM|Ankylosis of joint, pelvic region and thigh|Ankylosis of joint, pelvic region and thigh
C0158123|T047|AB|718.55|ICD9CM|Ankylosis-pelvis|Ankylosis-pelvis
C0158124|T020|PT|718.56|ICD9CM|Ankylosis of joint, lower leg|Ankylosis of joint, lower leg
C0158124|T020|AB|718.56|ICD9CM|Ankylosis-lower/leg|Ankylosis-lower/leg
C1963544|T020|PT|718.57|ICD9CM|Ankylosis of joint, ankle and foot|Ankylosis of joint, ankle and foot
C1963544|T020|AB|718.57|ICD9CM|Ankylosis-ankle|Ankylosis-ankle
C0158126|T047|PT|718.58|ICD9CM|Ankylosis of joint, other specified sites|Ankylosis of joint, other specified sites
C0158126|T047|AB|718.58|ICD9CM|Ankylosis-joint NEC|Ankylosis-joint NEC
C0158127|T047|PT|718.59|ICD9CM|Ankylosis of joint, multiple sites|Ankylosis of joint, multiple sites
C0158127|T047|AB|718.59|ICD9CM|Ankylosis-mult joints|Ankylosis-mult joints
C0158128|T047|HT|718.6|ICD9CM|Unspecified intrapelvic protrusion of acetabulum|Unspecified intrapelvic protrusion of acetabulum
C0158129|T047|AB|718.65|ICD9CM|Protrusio acetabuli NOS|Protrusio acetabuli NOS
C0158129|T047|PT|718.65|ICD9CM|Unspecified intrapelvic protrusion of acetabulum, pelvic region and thigh|Unspecified intrapelvic protrusion of acetabulum, pelvic region and thigh
C1145757|T047|HT|718.7|ICD9CM|Developmental dislocation of joint|Developmental dislocation of joint
C1176349|T047|AB|718.70|ICD9CM|Dev dislocat jt site NOS|Dev dislocat jt site NOS
C1176349|T047|PT|718.70|ICD9CM|Developmental dislocation of joint, site unspecified|Developmental dislocation of joint, site unspecified
C1176350|T047|AB|718.71|ICD9CM|Dev dislocat joint-shldr|Dev dislocat joint-shldr
C1176350|T047|PT|718.71|ICD9CM|Developmental dislocation of joint, shoulder region|Developmental dislocation of joint, shoulder region
C1176351|T047|AB|718.72|ICD9CM|Dev dislocat jt-up/arm|Dev dislocat jt-up/arm
C1176351|T047|PT|718.72|ICD9CM|Developmental dislocation of joint, upper arm|Developmental dislocation of joint, upper arm
C1176352|T047|AB|718.73|ICD9CM|Dev dislocat jt-forearm|Dev dislocat jt-forearm
C1176352|T047|PT|718.73|ICD9CM|Developmental dislocation of joint, forearm|Developmental dislocation of joint, forearm
C1176353|T047|AB|718.74|ICD9CM|Dev dislocat joint-hand|Dev dislocat joint-hand
C1176353|T047|PT|718.74|ICD9CM|Developmental dislocation of joint, hand|Developmental dislocation of joint, hand
C1176354|T047|AB|718.75|ICD9CM|Dev dis jt-pelvic/thigh|Dev dis jt-pelvic/thigh
C1176354|T047|PT|718.75|ICD9CM|Developmental dislocation of joint, pelvic region and thigh|Developmental dislocation of joint, pelvic region and thigh
C1176355|T047|AB|718.76|ICD9CM|Dev disloc jt-lower leg|Dev disloc jt-lower leg
C1176355|T047|PT|718.76|ICD9CM|Developmental dislocation of joint, lower leg|Developmental dislocation of joint, lower leg
C1176356|T047|AB|718.77|ICD9CM|Dev disloc jt-ankle/foot|Dev disloc jt-ankle/foot
C1176356|T047|PT|718.77|ICD9CM|Developmental dislocation of joint, ankle and foot|Developmental dislocation of joint, ankle and foot
C1176357|T047|AB|718.78|ICD9CM|Dev disloc jt-site NEC|Dev disloc jt-site NEC
C1176357|T047|PT|718.78|ICD9CM|Developmental dislocation of joint, other specified sites|Developmental dislocation of joint, other specified sites
C1176358|T047|AB|718.79|ICD9CM|Dev disloc jt-mult sites|Dev disloc jt-mult sites
C1176358|T047|PT|718.79|ICD9CM|Developmental dislocation of joint, multiple sites|Developmental dislocation of joint, multiple sites
C0869063|T047|HT|718.8|ICD9CM|Other joint derangement, not elsewhere classified|Other joint derangement, not elsewhere classified
C0869063|T047|AB|718.80|ICD9CM|Jt derangmnt NEC-unsp jt|Jt derangmnt NEC-unsp jt
C0869063|T047|PT|718.80|ICD9CM|Other joint derangement, not elsewhere classified, site unspecified|Other joint derangement, not elsewhere classified, site unspecified
C0869296|T190|AB|718.81|ICD9CM|Jt derangment NEC-shlder|Jt derangment NEC-shlder
C0869296|T190|PT|718.81|ICD9CM|Other joint derangement, not elsewhere classified, shoulder region|Other joint derangement, not elsewhere classified, shoulder region
C0869298|T190|AB|718.82|ICD9CM|Jt derangment NEC-up/arm|Jt derangment NEC-up/arm
C0869298|T190|PT|718.82|ICD9CM|Other joint derangement, not elsewhere classified, upper arm|Other joint derangement, not elsewhere classified, upper arm
C0869300|T190|AB|718.83|ICD9CM|Jt derangmnt NEC-forearm|Jt derangmnt NEC-forearm
C0869300|T190|PT|718.83|ICD9CM|Other joint derangement, not elsewhere classified, forearm|Other joint derangement, not elsewhere classified, forearm
C0869426|T190|AB|718.84|ICD9CM|Jt derangement NEC-hand|Jt derangement NEC-hand
C0869426|T190|PT|718.84|ICD9CM|Other joint derangement, not elsewhere classified, hand|Other joint derangement, not elsewhere classified, hand
C0869428|T190|AB|718.85|ICD9CM|Jt derangment NEC-pelvis|Jt derangment NEC-pelvis
C0869428|T190|PT|718.85|ICD9CM|Other joint derangement, not elsewhere classified, pelvic region and thigh|Other joint derangement, not elsewhere classified, pelvic region and thigh
C0869430|T190|AB|718.86|ICD9CM|Jt derangement NEC-l/leg|Jt derangement NEC-l/leg
C0869430|T190|PT|718.86|ICD9CM|Other joint derangement, not elsewhere classified, lower leg|Other joint derangement, not elsewhere classified, lower leg
C0869432|T190|AB|718.87|ICD9CM|Jt derangement NEC-ankle|Jt derangement NEC-ankle
C0869432|T190|PT|718.87|ICD9CM|Other joint derangement, not elsewhere classified, ankle and foot|Other joint derangement, not elsewhere classified, ankle and foot
C0869434|T190|AB|718.88|ICD9CM|Jt derangment NEC-oth jt|Jt derangment NEC-oth jt
C0869434|T190|PT|718.88|ICD9CM|Other joint derangement, not elsewhere classified, other specified sites|Other joint derangement, not elsewhere classified, other specified sites
C0869436|T190|AB|718.89|ICD9CM|Jt derangement NEC-mult|Jt derangement NEC-mult
C0869436|T190|PT|718.89|ICD9CM|Other joint derangement, not elsewhere classified, multiple sites|Other joint derangement, not elsewhere classified, multiple sites
C0158140|T047|HT|718.9|ICD9CM|Unspecified derangement of joint|Unspecified derangement of joint
C0158140|T047|AB|718.90|ICD9CM|Jt derangmnt NOS-unsp jt|Jt derangmnt NOS-unsp jt
C0158140|T047|PT|718.90|ICD9CM|Unspecified derangement of joint, site unspecified|Unspecified derangement of joint, site unspecified
C0409278|T190|AB|718.91|ICD9CM|Jt derangment NOS-shlder|Jt derangment NOS-shlder
C0409278|T190|PT|718.91|ICD9CM|Unspecified derangement of joint, shoulder region|Unspecified derangement of joint, shoulder region
C0409277|T190|AB|718.92|ICD9CM|Jt derangment NOS-up/arm|Jt derangment NOS-up/arm
C0409277|T190|PT|718.92|ICD9CM|Unspecified derangement of joint, upper arm|Unspecified derangement of joint, upper arm
C0409276|T190|AB|718.93|ICD9CM|Jt derangmnt NOS-forearm|Jt derangmnt NOS-forearm
C0409276|T190|PT|718.93|ICD9CM|Unspecified derangement of joint, forearm|Unspecified derangement of joint, forearm
C0409275|T047|AB|718.94|ICD9CM|Jt derangement NOS-hand|Jt derangement NOS-hand
C0409275|T047|PT|718.94|ICD9CM|Unspecified derangement of joint, hand|Unspecified derangement of joint, hand
C0409274|T190|AB|718.95|ICD9CM|Jt derangment NOS-pelvis|Jt derangment NOS-pelvis
C0409274|T190|PT|718.95|ICD9CM|Unspecified derangement of joint, pelvic region and thigh|Unspecified derangement of joint, pelvic region and thigh
C0409273|T047|AB|718.97|ICD9CM|Jt derangement NOS-ankle|Jt derangement NOS-ankle
C0409273|T047|PT|718.97|ICD9CM|Unspecified derangement of joint, ankle and foot|Unspecified derangement of joint, ankle and foot
C0409272|T190|AB|718.98|ICD9CM|Jt derangment NOS-oth jt|Jt derangment NOS-oth jt
C0409272|T190|PT|718.98|ICD9CM|Unspecified derangement of joint, other specified sites|Unspecified derangement of joint, other specified sites
C0409271|T047|AB|718.99|ICD9CM|Jt derangement NOS-mult|Jt derangement NOS-mult
C0409271|T047|PT|718.99|ICD9CM|Unspecified derangement of joint, multiple sites|Unspecified derangement of joint, multiple sites
C1442831|T047|HT|719|ICD9CM|Other and unspecified disorders of joint|Other and unspecified disorders of joint
C1253936|T046|HT|719.0|ICD9CM|Effusion of joint|Effusion of joint
C1253936|T046|PT|719.00|ICD9CM|Effusion of joint, site unspecified|Effusion of joint, site unspecified
C1253936|T046|AB|719.00|ICD9CM|Joint effusion-unspec|Joint effusion-unspec
C0158150|T046|PT|719.01|ICD9CM|Effusion of joint, shoulder region|Effusion of joint, shoulder region
C0158150|T046|AB|719.01|ICD9CM|Joint effusion-shlder|Joint effusion-shlder
C0158151|T046|PT|719.02|ICD9CM|Effusion of joint, upper arm|Effusion of joint, upper arm
C0158151|T046|AB|719.02|ICD9CM|Joint effusion-up/arm|Joint effusion-up/arm
C0158152|T046|PT|719.03|ICD9CM|Effusion of joint, forearm|Effusion of joint, forearm
C0158152|T046|AB|719.03|ICD9CM|Joint effusion-forearm|Joint effusion-forearm
C0158153|T046|PT|719.04|ICD9CM|Effusion of joint, hand|Effusion of joint, hand
C0158153|T046|AB|719.04|ICD9CM|Joint effusion-hand|Joint effusion-hand
C0554588|T046|PT|719.05|ICD9CM|Effusion of joint, pelvic region and thigh|Effusion of joint, pelvic region and thigh
C0554588|T046|AB|719.05|ICD9CM|Joint effusion-pelvis|Joint effusion-pelvis
C0158155|T046|PT|719.06|ICD9CM|Effusion of joint, lower leg|Effusion of joint, lower leg
C0158155|T046|AB|719.06|ICD9CM|Joint effusion-l/leg|Joint effusion-l/leg
C0158156|T046|PT|719.07|ICD9CM|Effusion of joint, ankle and foot|Effusion of joint, ankle and foot
C0158156|T046|AB|719.07|ICD9CM|Joint effusion-ankle|Joint effusion-ankle
C0158157|T184|PT|719.08|ICD9CM|Effusion of joint, other specified sites|Effusion of joint, other specified sites
C0158157|T184|AB|719.08|ICD9CM|Joint effusion-jt NEC|Joint effusion-jt NEC
C0158158|T046|PT|719.09|ICD9CM|Effusion of joint, multiple sites|Effusion of joint, multiple sites
C0158158|T046|AB|719.09|ICD9CM|Joint effusion-mult jts|Joint effusion-mult jts
C0018924|T046|HT|719.1|ICD9CM|Hemarthrosis|Hemarthrosis
C0018924|T046|AB|719.10|ICD9CM|Hemarthrosis-unspec|Hemarthrosis-unspec
C0018924|T046|PT|719.10|ICD9CM|Hemarthrosis, site unspecified|Hemarthrosis, site unspecified
C0158159|T047|AB|719.11|ICD9CM|Hemarthrosis-shlder|Hemarthrosis-shlder
C0158159|T047|PT|719.11|ICD9CM|Hemarthrosis, shoulder region|Hemarthrosis, shoulder region
C0263836|T047|AB|719.12|ICD9CM|Hemarthrosis-up/arm|Hemarthrosis-up/arm
C0263836|T047|PT|719.12|ICD9CM|Hemarthrosis, upper arm|Hemarthrosis, upper arm
C0263837|T047|AB|719.13|ICD9CM|Hemarthrosis-forearm|Hemarthrosis-forearm
C0263837|T047|PT|719.13|ICD9CM|Hemarthrosis, forearm|Hemarthrosis, forearm
C0158162|T047|AB|719.14|ICD9CM|Hemarthrosis-hand|Hemarthrosis-hand
C0158162|T047|PT|719.14|ICD9CM|Hemarthrosis, hand|Hemarthrosis, hand
C0263838|T046|AB|719.15|ICD9CM|Hemarthrosis-pelvis|Hemarthrosis-pelvis
C0263838|T046|PT|719.15|ICD9CM|Hemarthrosis, pelvic region and thigh|Hemarthrosis, pelvic region and thigh
C0263840|T047|AB|719.16|ICD9CM|Hemarthrosis-l/leg|Hemarthrosis-l/leg
C0263840|T047|PT|719.16|ICD9CM|Hemarthrosis, lower leg|Hemarthrosis, lower leg
C0263841|T033|AB|719.17|ICD9CM|Hemarthrosis-ankle|Hemarthrosis-ankle
C0263841|T033|PT|719.17|ICD9CM|Hemarthrosis, ankle and foot|Hemarthrosis, ankle and foot
C0473719|T046|AB|719.18|ICD9CM|Hemarthrosis-jt NEC|Hemarthrosis-jt NEC
C0473719|T046|PT|719.18|ICD9CM|Hemarthrosis, other specified sites|Hemarthrosis, other specified sites
C0158167|T046|AB|719.19|ICD9CM|Hemarthrosis-mult jts|Hemarthrosis-mult jts
C0158167|T046|PT|719.19|ICD9CM|Hemarthrosis, multiple sites|Hemarthrosis, multiple sites
C0158168|T047|HT|719.2|ICD9CM|Villonodular synovitis|Villonodular synovitis
C0158168|T047|AB|719.20|ICD9CM|Villonod synovit-unspec|Villonod synovit-unspec
C0158168|T047|PT|719.20|ICD9CM|Villonodular synovitis, site unspecified|Villonodular synovitis, site unspecified
C0158169|T047|AB|719.21|ICD9CM|Villonod synovit-shlder|Villonod synovit-shlder
C0158169|T047|PT|719.21|ICD9CM|Villonodular synovitis, shoulder region|Villonodular synovitis, shoulder region
C0409787|T047|AB|719.22|ICD9CM|Villonod synovit-up/arm|Villonod synovit-up/arm
C0409787|T047|PT|719.22|ICD9CM|Villonodular synovitis, upper arm|Villonodular synovitis, upper arm
C0409784|T047|AB|719.23|ICD9CM|Villonod synovit-forearm|Villonod synovit-forearm
C0409784|T047|PT|719.23|ICD9CM|Villonodular synovitis, forearm|Villonodular synovitis, forearm
C0409780|T191|AB|719.24|ICD9CM|Villonod synovit-hand|Villonod synovit-hand
C0409780|T191|PT|719.24|ICD9CM|Villonodular synovitis, hand|Villonodular synovitis, hand
C0409775|T047|AB|719.25|ICD9CM|Villonod synovit-pelvis|Villonod synovit-pelvis
C0409775|T047|PT|719.25|ICD9CM|Villonodular synovitis, pelvic region and thigh|Villonodular synovitis, pelvic region and thigh
C0409774|T047|AB|719.26|ICD9CM|Villonod synovit-l/leg|Villonod synovit-l/leg
C0409774|T047|PT|719.26|ICD9CM|Villonodular synovitis, lower leg|Villonodular synovitis, lower leg
C0158175|T047|AB|719.27|ICD9CM|Villonod synovit-ankle|Villonod synovit-ankle
C0158175|T047|PT|719.27|ICD9CM|Villonodular synovitis, ankle and foot|Villonodular synovitis, ankle and foot
C0409765|T047|AB|719.28|ICD9CM|Villonod synovit-jt NEC|Villonod synovit-jt NEC
C0409765|T047|PT|719.28|ICD9CM|Villonodular synovitis, other specified sites|Villonodular synovitis, other specified sites
C0837909|T191|AB|719.29|ICD9CM|Villonod synovit-mult jt|Villonod synovit-mult jt
C0837909|T191|PT|719.29|ICD9CM|Villonodular synovitis, multiple sites|Villonodular synovitis, multiple sites
C0085574|T047|HT|719.3|ICD9CM|Palindromic rheumatism|Palindromic rheumatism
C0085574|T047|AB|719.30|ICD9CM|Palindrom rheum-unspec|Palindrom rheum-unspec
C0085574|T047|PT|719.30|ICD9CM|Palindromic rheumatism, site unspecified|Palindromic rheumatism, site unspecified
C0158178|T046|AB|719.31|ICD9CM|Palindrom rheum-shlder|Palindrom rheum-shlder
C0158178|T046|PT|719.31|ICD9CM|Palindromic rheumatism, shoulder region|Palindromic rheumatism, shoulder region
C0409663|T047|AB|719.32|ICD9CM|Palindrom rheum-up/arm|Palindrom rheum-up/arm
C0409663|T047|PT|719.32|ICD9CM|Palindromic rheumatism, upper arm|Palindromic rheumatism, upper arm
C0409662|T047|AB|719.33|ICD9CM|Palindrom rheum-forearm|Palindrom rheum-forearm
C0409662|T047|PT|719.33|ICD9CM|Palindromic rheumatism, forearm|Palindromic rheumatism, forearm
C0158181|T047|AB|719.34|ICD9CM|Palindrom rheum-hand|Palindrom rheum-hand
C0158181|T047|PT|719.34|ICD9CM|Palindromic rheumatism, hand|Palindromic rheumatism, hand
C0409661|T047|AB|719.35|ICD9CM|Palindrom rheum-pelvis|Palindrom rheum-pelvis
C0409661|T047|PT|719.35|ICD9CM|Palindromic rheumatism, pelvic region and thigh|Palindromic rheumatism, pelvic region and thigh
C0409660|T047|AB|719.36|ICD9CM|Palindrom rheum-l/leg|Palindrom rheum-l/leg
C0409660|T047|PT|719.36|ICD9CM|Palindromic rheumatism, lower leg|Palindromic rheumatism, lower leg
C0409659|T047|AB|719.37|ICD9CM|Palindrom rheum-ankle|Palindrom rheum-ankle
C0409659|T047|PT|719.37|ICD9CM|Palindromic rheumatism, ankle and foot|Palindromic rheumatism, ankle and foot
C0409658|T047|AB|719.38|ICD9CM|Palindrom rheum-jt NEC|Palindrom rheum-jt NEC
C0409658|T047|PT|719.38|ICD9CM|Palindromic rheumatism, other specified sites|Palindromic rheumatism, other specified sites
C0158186|T047|AB|719.39|ICD9CM|Palindrom rheum-mult jts|Palindrom rheum-mult jts
C0158186|T047|PT|719.39|ICD9CM|Palindromic rheumatism, multiple sites|Palindromic rheumatism, multiple sites
C0003862|T184|HT|719.4|ICD9CM|Pain in joint|Pain in joint
C0003862|T184|AB|719.40|ICD9CM|Joint pain-unspec|Joint pain-unspec
C0003862|T184|PT|719.40|ICD9CM|Pain in joint, site unspecified|Pain in joint, site unspecified
C0838222|T184|AB|719.41|ICD9CM|Joint pain-shlder|Joint pain-shlder
C0838222|T184|PT|719.41|ICD9CM|Pain in joint, shoulder region|Pain in joint, shoulder region
C0838223|T184|AB|719.42|ICD9CM|Joint pain-up/arm|Joint pain-up/arm
C0838223|T184|PT|719.42|ICD9CM|Pain in joint, upper arm|Pain in joint, upper arm
C0838224|T184|AB|719.43|ICD9CM|Joint pain-forearm|Joint pain-forearm
C0838224|T184|PT|719.43|ICD9CM|Pain in joint, forearm|Pain in joint, forearm
C0423665|T184|AB|719.44|ICD9CM|Joint pain-hand|Joint pain-hand
C0423665|T184|PT|719.44|ICD9CM|Pain in joint, hand|Pain in joint, hand
C0838226|T184|AB|719.45|ICD9CM|Joint pain-pelvis|Joint pain-pelvis
C0838226|T184|PT|719.45|ICD9CM|Pain in joint, pelvic region and thigh|Pain in joint, pelvic region and thigh
C0838227|T184|AB|719.46|ICD9CM|Joint pain-l/leg|Joint pain-l/leg
C0838227|T184|PT|719.46|ICD9CM|Pain in joint, lower leg|Pain in joint, lower leg
C2919460|T184|AB|719.47|ICD9CM|Joint pain-ankle|Joint pain-ankle
C2919460|T184|PT|719.47|ICD9CM|Pain in joint, ankle and foot|Pain in joint, ankle and foot
C0158194|T184|AB|719.48|ICD9CM|Joint pain-jt NEC|Joint pain-jt NEC
C0158194|T184|PT|719.48|ICD9CM|Pain in joint, other specified sites|Pain in joint, other specified sites
C0162296|T047|AB|719.49|ICD9CM|Joint pain-mult jts|Joint pain-mult jts
C0162296|T047|PT|719.49|ICD9CM|Pain in joint, multiple sites|Pain in joint, multiple sites
C0869450|T184|HT|719.5|ICD9CM|Stiffness of joint, not elsewhere classified|Stiffness of joint, not elsewhere classified
C0158195|T047|AB|719.50|ICD9CM|Jt stiffness NEC-unspec|Jt stiffness NEC-unspec
C0158195|T047|PT|719.50|ICD9CM|Stiffness of joint, not elsewhere classified, site unspecified|Stiffness of joint, not elsewhere classified, site unspecified
C0158196|T047|AB|719.51|ICD9CM|Jt stiffness NEC-shlder|Jt stiffness NEC-shlder
C0158196|T047|PT|719.51|ICD9CM|Stiffness of joint, not elsewhere classified, shoulder region|Stiffness of joint, not elsewhere classified, shoulder region
C0158197|T047|AB|719.52|ICD9CM|Jt stiffness NEC-up/arm|Jt stiffness NEC-up/arm
C0158197|T047|PT|719.52|ICD9CM|Stiffness of joint, not elsewhere classified, upper arm|Stiffness of joint, not elsewhere classified, upper arm
C0158198|T047|AB|719.53|ICD9CM|Jt stiffnes NEC-forearm|Jt stiffnes NEC-forearm
C0158198|T047|PT|719.53|ICD9CM|Stiffness of joint, not elsewhere classified, forearm|Stiffness of joint, not elsewhere classified, forearm
C0158199|T047|AB|719.54|ICD9CM|Jt stiffness NEC-hand|Jt stiffness NEC-hand
C0158199|T047|PT|719.54|ICD9CM|Stiffness of joint, not elsewhere classified, hand|Stiffness of joint, not elsewhere classified, hand
C0158200|T047|AB|719.55|ICD9CM|Jt stiffness NEC-pelvis|Jt stiffness NEC-pelvis
C0158200|T047|PT|719.55|ICD9CM|Stiffness of joint, not elsewhere classified, pelvic region and thigh|Stiffness of joint, not elsewhere classified, pelvic region and thigh
C0158201|T047|AB|719.56|ICD9CM|Jt stiffness NEC-l/leg|Jt stiffness NEC-l/leg
C0158201|T047|PT|719.56|ICD9CM|Stiffness of joint, not elsewhere classified, lower leg|Stiffness of joint, not elsewhere classified, lower leg
C0158202|T047|AB|719.57|ICD9CM|Jt stiffness NEC-ankle|Jt stiffness NEC-ankle
C0158202|T047|PT|719.57|ICD9CM|Stiffness of joint, not elsewhere classified, ankle and foot|Stiffness of joint, not elsewhere classified, ankle and foot
C0158203|T047|AB|719.58|ICD9CM|Jt stiffness NEC-oth jt|Jt stiffness NEC-oth jt
C0158203|T047|PT|719.58|ICD9CM|Stiffness of joint, not elsewhere classified, other specified sites|Stiffness of joint, not elsewhere classified, other specified sites
C0158204|T047|AB|719.59|ICD9CM|Jt stiffness NEC-mult jt|Jt stiffness NEC-mult jt
C0158204|T047|PT|719.59|ICD9CM|Stiffness of joint, not elsewhere classified, multiple sites|Stiffness of joint, not elsewhere classified, multiple sites
C0158205|T184|HT|719.6|ICD9CM|Other symptoms referable to joint|Other symptoms referable to joint
C0375492|T184|AB|719.60|ICD9CM|Joint sympt NEC-unsp jt|Joint sympt NEC-unsp jt
C0375492|T184|PT|719.60|ICD9CM|Other symptoms referable to joint, site unspecified|Other symptoms referable to joint, site unspecified
C0158206|T184|AB|719.61|ICD9CM|Joint symptom NEC-shlder|Joint symptom NEC-shlder
C0158206|T184|PT|719.61|ICD9CM|Other symptoms referable to joint, shoulder region|Other symptoms referable to joint, shoulder region
C0158207|T184|AB|719.62|ICD9CM|Joint symptom NEC-up/arm|Joint symptom NEC-up/arm
C0158207|T184|PT|719.62|ICD9CM|Other symptoms referable to joint, upper arm|Other symptoms referable to joint, upper arm
C0158208|T184|AB|719.63|ICD9CM|Joint sympt NEC-forearm|Joint sympt NEC-forearm
C0158208|T184|PT|719.63|ICD9CM|Other symptoms referable to joint, forearm|Other symptoms referable to joint, forearm
C0158209|T184|AB|719.64|ICD9CM|Joint symptom NEC-hand|Joint symptom NEC-hand
C0158209|T184|PT|719.64|ICD9CM|Other symptoms referable to joint, hand|Other symptoms referable to joint, hand
C0158210|T184|AB|719.65|ICD9CM|Joint symptom NEC-pelvis|Joint symptom NEC-pelvis
C0158210|T184|PT|719.65|ICD9CM|Other symptoms referable to joint, pelvic region and thigh|Other symptoms referable to joint, pelvic region and thigh
C0158211|T184|AB|719.66|ICD9CM|Joint symptom NEC-l/leg|Joint symptom NEC-l/leg
C0158211|T184|PT|719.66|ICD9CM|Other symptoms referable to joint, lower leg|Other symptoms referable to joint, lower leg
C0158212|T184|AB|719.67|ICD9CM|Joint symptom NEC-ankle|Joint symptom NEC-ankle
C0158212|T184|PT|719.67|ICD9CM|Other symptoms referable to joint, ankle and foot|Other symptoms referable to joint, ankle and foot
C0158213|T184|AB|719.68|ICD9CM|Joint symptom NEC-oth jt|Joint symptom NEC-oth jt
C0158213|T184|PT|719.68|ICD9CM|Other symptoms referable to joint, other specified sites|Other symptoms referable to joint, other specified sites
C0158214|T184|AB|719.69|ICD9CM|Joint sympt NEC-mult jts|Joint sympt NEC-mult jts
C0158214|T184|PT|719.69|ICD9CM|Other symptoms referable to joint, multiple sites|Other symptoms referable to joint, multiple sites
C0311394|T033|AB|719.7|ICD9CM|Difficulty in walking|Difficulty in walking
C0311394|T033|PT|719.7|ICD9CM|Difficulty in walking|Difficulty in walking
C0029746|T047|HT|719.8|ICD9CM|Other specified disorders of joint|Other specified disorders of joint
C0869062|T047|AB|719.80|ICD9CM|Joint dis NEC-unspec|Joint dis NEC-unspec
C0869062|T047|PT|719.80|ICD9CM|Other specified disorders of joint, site unspecified|Other specified disorders of joint, site unspecified
C0158222|T047|AB|719.81|ICD9CM|Joint dis NEC-shlder|Joint dis NEC-shlder
C0158222|T047|PT|719.81|ICD9CM|Other specified disorders of joint, shoulder region|Other specified disorders of joint, shoulder region
C0158223|T047|AB|719.82|ICD9CM|Joint dis NEC-up/arm|Joint dis NEC-up/arm
C0158223|T047|PT|719.82|ICD9CM|Other specified disorders of joint, upper arm|Other specified disorders of joint, upper arm
C0158224|T047|AB|719.83|ICD9CM|Joint dis NEC-forearm|Joint dis NEC-forearm
C0158224|T047|PT|719.83|ICD9CM|Other specified disorders of joint, forearm|Other specified disorders of joint, forearm
C0158225|T047|AB|719.84|ICD9CM|Joint dis NEC-hand|Joint dis NEC-hand
C0158225|T047|PT|719.84|ICD9CM|Other specified disorders of joint, hand|Other specified disorders of joint, hand
C0158226|T047|AB|719.85|ICD9CM|Joint dis NEC-pelvis|Joint dis NEC-pelvis
C0158226|T047|PT|719.85|ICD9CM|Other specified disorders of joint, pelvic region and thigh|Other specified disorders of joint, pelvic region and thigh
C0158227|T047|AB|719.86|ICD9CM|Joint dis NEC-l/leg|Joint dis NEC-l/leg
C0158227|T047|PT|719.86|ICD9CM|Other specified disorders of joint, lower leg|Other specified disorders of joint, lower leg
C0158228|T047|AB|719.87|ICD9CM|Joint dis NEC-ankle|Joint dis NEC-ankle
C0158228|T047|PT|719.87|ICD9CM|Other specified disorders of joint, ankle and foot|Other specified disorders of joint, ankle and foot
C0158229|T047|AB|719.88|ICD9CM|Joint dis NEC-oth jt|Joint dis NEC-oth jt
C0158229|T047|PT|719.88|ICD9CM|Other specified disorders of joint, other specified sites|Other specified disorders of joint, other specified sites
C0158230|T047|AB|719.89|ICD9CM|Joint dis NEC-mult jts|Joint dis NEC-mult jts
C0158230|T047|PT|719.89|ICD9CM|Other specified disorders of joint, multiple sites|Other specified disorders of joint, multiple sites
C0022408|T047|HT|719.9|ICD9CM|Unspecified disorder of joint|Unspecified disorder of joint
C0022408|T047|AB|719.90|ICD9CM|Joint dis NOS-unspec jt|Joint dis NOS-unspec jt
C0022408|T047|PT|719.90|ICD9CM|Unspecified disorder of joint, site unspecified|Unspecified disorder of joint, site unspecified
C0158231|T047|AB|719.91|ICD9CM|Joint dis NOS-shlder|Joint dis NOS-shlder
C0158231|T047|PT|719.91|ICD9CM|Unspecified disorder of joint, shoulder region|Unspecified disorder of joint, shoulder region
C0158232|T047|AB|719.92|ICD9CM|Joint dis NOS-up/arm|Joint dis NOS-up/arm
C0158232|T047|PT|719.92|ICD9CM|Unspecified disorder of joint, upper arm|Unspecified disorder of joint, upper arm
C0158233|T047|AB|719.93|ICD9CM|Joint dis NOS-forearm|Joint dis NOS-forearm
C0158233|T047|PT|719.93|ICD9CM|Unspecified disorder of joint, forearm|Unspecified disorder of joint, forearm
C0158234|T047|AB|719.94|ICD9CM|Joint dis NOS-hand|Joint dis NOS-hand
C0158234|T047|PT|719.94|ICD9CM|Unspecified disorder of joint, hand|Unspecified disorder of joint, hand
C0158235|T047|AB|719.95|ICD9CM|Joint dis NOS-pelvis|Joint dis NOS-pelvis
C0158235|T047|PT|719.95|ICD9CM|Unspecified disorder of joint, pelvic region and thigh|Unspecified disorder of joint, pelvic region and thigh
C0158236|T047|AB|719.96|ICD9CM|Joint dis NOS-l/leg|Joint dis NOS-l/leg
C0158236|T047|PT|719.96|ICD9CM|Unspecified disorder of joint, lower leg|Unspecified disorder of joint, lower leg
C0409264|T047|AB|719.97|ICD9CM|Joint dis NOS-ankle|Joint dis NOS-ankle
C0409264|T047|PT|719.97|ICD9CM|Unspecified disorder of joint, ankle and foot|Unspecified disorder of joint, ankle and foot
C0489969|T047|AB|719.98|ICD9CM|Joint dis NOS-oth jt|Joint dis NOS-oth jt
C0489969|T047|PT|719.98|ICD9CM|Unspecified disorder of joint, other specified sites|Unspecified disorder of joint, other specified sites
C0158239|T047|AB|719.99|ICD9CM|Joint dis NOS-mult jts|Joint dis NOS-mult jts
C0158239|T047|PT|719.99|ICD9CM|Unspecified disorder of joint, multiple sites|Unspecified disorder of joint, multiple sites
C0003089|T047|HT|720|ICD9CM|Ankylosing spondylitis and other inflammatory spondylopathies|Ankylosing spondylitis and other inflammatory spondylopathies
C3241938|T047|HT|720-724.99|ICD9CM|DORSOPATHIES|DORSOPATHIES
C0038013|T047|AB|720.0|ICD9CM|Ankylosing spondylitis|Ankylosing spondylitis
C0038013|T047|PT|720.0|ICD9CM|Ankylosing spondylitis|Ankylosing spondylitis
C0152090|T047|AB|720.1|ICD9CM|Spinal enthesopathy|Spinal enthesopathy
C0152090|T047|PT|720.1|ICD9CM|Spinal enthesopathy|Spinal enthesopathy
C0868862|T047|AB|720.2|ICD9CM|Sacroiliitis NEC|Sacroiliitis NEC
C0868862|T047|PT|720.2|ICD9CM|Sacroiliitis, not elsewhere classified|Sacroiliitis, not elsewhere classified
C0029644|T047|HT|720.8|ICD9CM|Other inflammatory spondylopathies|Other inflammatory spondylopathies
C0021396|T047|PT|720.81|ICD9CM|Inflammatory spondylopathies in diseases classified elsewhere|Inflammatory spondylopathies in diseases classified elsewhere
C0021396|T047|AB|720.81|ICD9CM|Spondylopathy in oth dis|Spondylopathy in oth dis
C0029644|T047|AB|720.89|ICD9CM|Inflam spondylopathy NEC|Inflam spondylopathy NEC
C0029644|T047|PT|720.89|ICD9CM|Other inflammatory spondylopathies|Other inflammatory spondylopathies
C0038012|T047|AB|720.9|ICD9CM|Inflam spondylopathy NOS|Inflam spondylopathy NOS
C0038012|T047|PT|720.9|ICD9CM|Unspecified inflammatory spondylopathy|Unspecified inflammatory spondylopathy
C0158240|T047|HT|721|ICD9CM|Spondylosis and allied disorders|Spondylosis and allied disorders
C0158241|T047|AB|721.0|ICD9CM|Cervical spondylosis|Cervical spondylosis
C0158241|T047|PT|721.0|ICD9CM|Cervical spondylosis without myelopathy|Cervical spondylosis without myelopathy
C0158242|T047|AB|721.1|ICD9CM|Cerv spondyl w myelopath|Cerv spondyl w myelopath
C0158242|T047|PT|721.1|ICD9CM|Cervical spondylosis with myelopathy|Cervical spondylosis with myelopathy
C0158243|T047|AB|721.2|ICD9CM|Thoracic spondylosis|Thoracic spondylosis
C0158243|T047|PT|721.2|ICD9CM|Thoracic spondylosis without myelopathy|Thoracic spondylosis without myelopathy
C0158244|T047|AB|721.3|ICD9CM|Lumbosacral spondylosis|Lumbosacral spondylosis
C0158244|T047|PT|721.3|ICD9CM|Lumbosacral spondylosis without myelopathy|Lumbosacral spondylosis without myelopathy
C0158245|T047|HT|721.4|ICD9CM|Thoracic or lumbar spondylosis with myelopathy|Thoracic or lumbar spondylosis with myelopathy
C0158246|T047|AB|721.41|ICD9CM|Spond compr thor sp cord|Spond compr thor sp cord
C0158246|T047|PT|721.41|ICD9CM|Spondylosis with myelopathy, thoracic region|Spondylosis with myelopathy, thoracic region
C0158247|T047|AB|721.42|ICD9CM|Spond compr lumb sp cord|Spond compr lumb sp cord
C0158247|T047|PT|721.42|ICD9CM|Spondylosis with myelopathy, lumbar region|Spondylosis with myelopathy, lumbar region
C0158248|T047|AB|721.5|ICD9CM|Kissing spine|Kissing spine
C0158248|T047|PT|721.5|ICD9CM|Kissing spine|Kissing spine
C0020498|T047|AB|721.6|ICD9CM|Ankyl vert hyperostosis|Ankyl vert hyperostosis
C0020498|T047|PT|721.6|ICD9CM|Ankylosing vertebral hyperostosis|Ankylosing vertebral hyperostosis
C0152088|T047|AB|721.7|ICD9CM|Traumatic spondylopathy|Traumatic spondylopathy
C0152088|T047|PT|721.7|ICD9CM|Traumatic spondylopathy|Traumatic spondylopathy
C0158249|T047|PT|721.8|ICD9CM|Other allied disorders of spine|Other allied disorders of spine
C0158249|T047|AB|721.8|ICD9CM|Spinal disorders NEC|Spinal disorders NEC
C0038019|T047|HT|721.9|ICD9CM|Spondylosis of unspecified site|Spondylosis of unspecified site
C0263851|T047|AB|721.90|ICD9CM|Spondylos NOS w/o myelop|Spondylos NOS w/o myelop
C0263851|T047|PT|721.90|ICD9CM|Spondylosis of unspecified site, without mention of myelopathy|Spondylosis of unspecified site, without mention of myelopathy
C0263853|T047|AB|721.91|ICD9CM|Spondylosis NOS w myelop|Spondylosis NOS w myelop
C0263853|T047|PT|721.91|ICD9CM|Spondylosis of unspecified site, with myelopathy|Spondylosis of unspecified site, with myelopathy
C0158252|T047|HT|722|ICD9CM|Intervertebral disc disorders|Intervertebral disc disorders
C0158253|T047|AB|722.0|ICD9CM|Cervical disc displacmnt|Cervical disc displacmnt
C0158253|T047|PT|722.0|ICD9CM|Displacement of cervical intervertebral disc without myelopathy|Displacement of cervical intervertebral disc without myelopathy
C0158254|T047|HT|722.1|ICD9CM|Displacement of thoracic or lumbar intervertebral disc without myelopathy|Displacement of thoracic or lumbar intervertebral disc without myelopathy
C0158255|T047|PT|722.10|ICD9CM|Displacement of lumbar intervertebral disc without myelopathy|Displacement of lumbar intervertebral disc without myelopathy
C0158255|T047|AB|722.10|ICD9CM|Lumbar disc displacement|Lumbar disc displacement
C0158256|T047|PT|722.11|ICD9CM|Displacement of thoracic intervertebral disc without myelopathy|Displacement of thoracic intervertebral disc without myelopathy
C0158256|T047|AB|722.11|ICD9CM|Thoracic disc displacmnt|Thoracic disc displacmnt
C1328971|T047|AB|722.2|ICD9CM|Disc displacement NOS|Disc displacement NOS
C1328971|T047|PT|722.2|ICD9CM|Displacement of intervertebral disc, site unspecified, without myelopathy|Displacement of intervertebral disc, site unspecified, without myelopathy
C0410632|T047|HT|722.3|ICD9CM|Schmorl's nodes|Schmorl's nodes
C0410632|T047|AB|722.30|ICD9CM|Schmorl's nodes NOS|Schmorl's nodes NOS
C0410632|T047|PT|722.30|ICD9CM|Schmorl's nodes, unspecified region|Schmorl's nodes, unspecified region
C0158259|T047|PT|722.31|ICD9CM|Schmorl's nodes, thoracic region|Schmorl's nodes, thoracic region
C0158259|T047|AB|722.31|ICD9CM|Schmorls node-thoracic|Schmorls node-thoracic
C0158260|T047|PT|722.32|ICD9CM|Schmorl's nodes, lumbar region|Schmorl's nodes, lumbar region
C0158260|T047|AB|722.32|ICD9CM|Schmorls node-lumbar|Schmorls node-lumbar
C0158261|T047|PT|722.39|ICD9CM|Schmorl's nodes, other region|Schmorl's nodes, other region
C0158261|T047|AB|722.39|ICD9CM|Schmorls node-region NEC|Schmorls node-region NEC
C0158262|T047|AB|722.4|ICD9CM|Cervical disc degen|Cervical disc degen
C0158262|T047|PT|722.4|ICD9CM|Degeneration of cervical intervertebral disc|Degeneration of cervical intervertebral disc
C0158263|T047|HT|722.5|ICD9CM|Degeneration of thoracic or lumbar intervertebral disc|Degeneration of thoracic or lumbar intervertebral disc
C0158264|T047|PT|722.51|ICD9CM|Degeneration of thoracic or thoracolumbar intervertebral disc|Degeneration of thoracic or thoracolumbar intervertebral disc
C0158264|T047|AB|722.51|ICD9CM|Thoracic disc degen|Thoracic disc degen
C0158265|T047|PT|722.52|ICD9CM|Degeneration of lumbar or lumbosacral intervertebral disc|Degeneration of lumbar or lumbosacral intervertebral disc
C0158265|T047|AB|722.52|ICD9CM|Lumb/lumbosac disc degen|Lumb/lumbosac disc degen
C0158266|T047|PT|722.6|ICD9CM|Degeneration of intervertebral disc, site unspecified|Degeneration of intervertebral disc, site unspecified
C0158266|T047|AB|722.6|ICD9CM|Disc degeneration NOS|Disc degeneration NOS
C0158267|T047|HT|722.7|ICD9CM|Intervertebral disc disorder with myelopathy|Intervertebral disc disorder with myelopathy
C0375497|T047|AB|722.70|ICD9CM|Disc dis w myelopath NOS|Disc dis w myelopath NOS
C0375497|T047|PT|722.70|ICD9CM|Intervertebral disc disorder with myelopathy, unspecified region|Intervertebral disc disorder with myelopathy, unspecified region
C0158268|T047|AB|722.71|ICD9CM|Cerv disc dis w myelopat|Cerv disc dis w myelopat
C0158268|T047|PT|722.71|ICD9CM|Intervertebral disc disorder with myelopathy, cervical region|Intervertebral disc disorder with myelopathy, cervical region
C0158269|T047|PT|722.72|ICD9CM|Intervertebral disc disorder with myelopathy, thoracic region|Intervertebral disc disorder with myelopathy, thoracic region
C0158269|T047|AB|722.72|ICD9CM|Thor disc dis w myelopat|Thor disc dis w myelopat
C0158270|T047|PT|722.73|ICD9CM|Intervertebral disc disorder with myelopathy, lumbar region|Intervertebral disc disorder with myelopathy, lumbar region
C0158270|T047|AB|722.73|ICD9CM|Lumb disc dis w myelopat|Lumb disc dis w myelopat
C0152089|T047|HT|722.8|ICD9CM|Postlaminectomy syndrome|Postlaminectomy syndrome
C0152089|T047|AB|722.80|ICD9CM|Postlaminectomy synd NOS|Postlaminectomy synd NOS
C0152089|T047|PT|722.80|ICD9CM|Postlaminectomy syndrome, unspecified region|Postlaminectomy syndrome, unspecified region
C0158272|T047|AB|722.81|ICD9CM|Postlaminect synd-cerv|Postlaminect synd-cerv
C0158272|T047|PT|722.81|ICD9CM|Postlaminectomy syndrome, cervical region|Postlaminectomy syndrome, cervical region
C0158273|T047|AB|722.82|ICD9CM|Postlaminect synd-thorac|Postlaminect synd-thorac
C0158273|T047|PT|722.82|ICD9CM|Postlaminectomy syndrome, thoracic region|Postlaminectomy syndrome, thoracic region
C0158274|T047|AB|722.83|ICD9CM|Postlaminect synd-lumbar|Postlaminect synd-lumbar
C0158274|T047|PT|722.83|ICD9CM|Postlaminectomy syndrome, lumbar region|Postlaminectomy syndrome, lumbar region
C0158275|T047|HT|722.9|ICD9CM|Other and unspecified disc disorder|Other and unspecified disc disorder
C0029497|T047|AB|722.90|ICD9CM|Disc dis NEC/NOS-unspec|Disc dis NEC/NOS-unspec
C0029497|T047|PT|722.90|ICD9CM|Other and unspecified disc disorder, unspecified region|Other and unspecified disc disorder, unspecified region
C0158276|T047|AB|722.91|ICD9CM|Disc dis NEC/NOS-cerv|Disc dis NEC/NOS-cerv
C0158276|T047|PT|722.91|ICD9CM|Other and unspecified disc disorder, cervical region|Other and unspecified disc disorder, cervical region
C0158277|T047|AB|722.92|ICD9CM|Disc dis NEC/NOS-thorac|Disc dis NEC/NOS-thorac
C0158277|T047|PT|722.92|ICD9CM|Other and unspecified disc disorder, thoracic region|Other and unspecified disc disorder, thoracic region
C0158278|T047|AB|722.93|ICD9CM|Disc dis NEC/NOS-lumbar|Disc dis NEC/NOS-lumbar
C0158278|T047|PT|722.93|ICD9CM|Other and unspecified disc disorder, lumbar region|Other and unspecified disc disorder, lumbar region
C0158279|T047|HT|723|ICD9CM|Other disorders of cervical region|Other disorders of cervical region
C0158280|T047|AB|723.0|ICD9CM|Cervical spinal stenosis|Cervical spinal stenosis
C0158280|T047|PT|723.0|ICD9CM|Spinal stenosis in cervical region|Spinal stenosis in cervical region
C0007859|T184|AB|723.1|ICD9CM|Cervicalgia|Cervicalgia
C0007859|T184|PT|723.1|ICD9CM|Cervicalgia|Cervicalgia
C2355645|T047|AB|723.2|ICD9CM|Cervicocranial syndrome|Cervicocranial syndrome
C2355645|T047|PT|723.2|ICD9CM|Cervicocranial syndrome|Cervicocranial syndrome
C0158281|T047|AB|723.3|ICD9CM|Cervicobrachial syndrome|Cervicobrachial syndrome
C0158281|T047|PT|723.3|ICD9CM|Cervicobrachial syndrome (diffuse)|Cervicobrachial syndrome (diffuse)
C1442952|T047|AB|723.4|ICD9CM|Brachial neuritis NOS|Brachial neuritis NOS
C1442952|T047|PT|723.4|ICD9CM|Brachial neuritis or radiculitis NOS|Brachial neuritis or radiculitis NOS
C0040485|T184|AB|723.5|ICD9CM|Torticollis NOS|Torticollis NOS
C0040485|T184|PT|723.5|ICD9CM|Torticollis, unspecified|Torticollis, unspecified
C0263013|T047|AB|723.6|ICD9CM|Panniculitis of neck|Panniculitis of neck
C0263013|T047|PT|723.6|ICD9CM|Panniculitis specified as affecting neck|Panniculitis specified as affecting neck
C0699899|T046|AB|723.7|ICD9CM|Ossification cerv lig|Ossification cerv lig
C0699899|T046|PT|723.7|ICD9CM|Ossification of posterior longitudinal ligament in cervical region|Ossification of posterior longitudinal ligament in cervical region
C0158284|T047|AB|723.8|ICD9CM|Cervical syndrome NEC|Cervical syndrome NEC
C0158284|T047|PT|723.8|ICD9CM|Other syndromes affecting cervical region|Other syndromes affecting cervical region
C0158285|T047|AB|723.9|ICD9CM|Neck disorder/sympt NOS|Neck disorder/sympt NOS
C0158285|T047|PT|723.9|ICD9CM|Unspecified musculoskeletal disorders and symptoms referable to neck|Unspecified musculoskeletal disorders and symptoms referable to neck
C0158298|T047|HT|724|ICD9CM|Other and unspecified disorders of back|Other and unspecified disorders of back
C0037947|T190|HT|724.0|ICD9CM|Spinal stenosis, other than cervical|Spinal stenosis, other than cervical
C0037944|T020|AB|724.00|ICD9CM|Spinal stenosis NOS|Spinal stenosis NOS
C0037944|T020|PT|724.00|ICD9CM|Spinal stenosis, unspecified region|Spinal stenosis, unspecified region
C0158287|T047|AB|724.01|ICD9CM|Spinal stenosis-thoracic|Spinal stenosis-thoracic
C0158287|T047|PT|724.01|ICD9CM|Spinal stenosis, thoracic region|Spinal stenosis, thoracic region
C2921108|T047|AB|724.02|ICD9CM|Spin sten,lumbr wo claud|Spin sten,lumbr wo claud
C2921108|T047|PT|724.02|ICD9CM|Spinal stenosis, lumbar region, without neurogenic claudication|Spinal stenosis, lumbar region, without neurogenic claudication
C2921109|T047|AB|724.03|ICD9CM|Spin sten,lumbr w claud|Spin sten,lumbr w claud
C2921109|T047|PT|724.03|ICD9CM|Spinal stenosis, lumbar region, with neurogenic claudication|Spinal stenosis, lumbar region, with neurogenic claudication
C0158289|T190|AB|724.09|ICD9CM|Spinal stenosis-oth site|Spinal stenosis-oth site
C0158289|T190|PT|724.09|ICD9CM|Spinal stenosis, other region|Spinal stenosis, other region
C0677061|T184|AB|724.1|ICD9CM|Pain in thoracic spine|Pain in thoracic spine
C0677061|T184|PT|724.1|ICD9CM|Pain in thoracic spine|Pain in thoracic spine
C0024031|T184|AB|724.2|ICD9CM|Lumbago|Lumbago
C0024031|T184|PT|724.2|ICD9CM|Lumbago|Lumbago
C0036396|T184|AB|724.3|ICD9CM|Sciatica|Sciatica
C0036396|T184|PT|724.3|ICD9CM|Sciatica|Sciatica
C0158291|T047|AB|724.4|ICD9CM|Lumbosacral neuritis NOS|Lumbosacral neuritis NOS
C0158291|T047|PT|724.4|ICD9CM|Thoracic or lumbosacral neuritis or radiculitis, unspecified|Thoracic or lumbosacral neuritis or radiculitis, unspecified
C0004604|T184|AB|724.5|ICD9CM|Backache NOS|Backache NOS
C0004604|T184|PT|724.5|ICD9CM|Backache, unspecified|Backache, unspecified
C0158292|T047|AB|724.6|ICD9CM|Disorders of sacrum|Disorders of sacrum
C0158292|T047|PT|724.6|ICD9CM|Disorders of sacrum|Disorders of sacrum
C0158293|T047|HT|724.7|ICD9CM|Disorders of coccyx|Disorders of coccyx
C0158293|T047|AB|724.70|ICD9CM|Disorder of coccyx NOS|Disorder of coccyx NOS
C0158293|T047|PT|724.70|ICD9CM|Unspecified disorder of coccyx|Unspecified disorder of coccyx
C0158295|T047|AB|724.71|ICD9CM|Hypermobility of coccyx|Hypermobility of coccyx
C0158295|T047|PT|724.71|ICD9CM|Hypermobility of coccyx|Hypermobility of coccyx
C0158296|T047|AB|724.79|ICD9CM|Disorder of coccyx NEC|Disorder of coccyx NEC
C0158296|T047|PT|724.79|ICD9CM|Other disorders of coccyx|Other disorders of coccyx
C0158297|T184|AB|724.8|ICD9CM|Other back symptoms|Other back symptoms
C0158297|T184|PT|724.8|ICD9CM|Other symptoms referable to back|Other symptoms referable to back
C0158298|T047|AB|724.9|ICD9CM|Back disorder NOS|Back disorder NOS
C0158298|T047|PT|724.9|ICD9CM|Other unspecified back disorders|Other unspecified back disorders
C0032533|T047|AB|725|ICD9CM|Polymyalgia rheumatica|Polymyalgia rheumatica
C0032533|T047|PT|725|ICD9CM|Polymyalgia rheumatica|Polymyalgia rheumatica
C0178305|T047|HT|725-729.99|ICD9CM|RHEUMATISM, EXCLUDING THE BACK|RHEUMATISM, EXCLUDING THE BACK
C1442902|T047|HT|726|ICD9CM|Peripheral enthesopathies and allied syndromes|Peripheral enthesopathies and allied syndromes
C0311223|T047|AB|726.0|ICD9CM|Adhesive capsulit shlder|Adhesive capsulit shlder
C0311223|T047|PT|726.0|ICD9CM|Adhesive capsulitis of shoulder|Adhesive capsulitis of shoulder
C0158301|T047|HT|726.1|ICD9CM|Rotator cuff syndrome of shoulder and allied disorders|Rotator cuff syndrome of shoulder and allied disorders
C0158302|T047|PT|726.10|ICD9CM|Disorders of bursae and tendons in shoulder region, unspecified|Disorders of bursae and tendons in shoulder region, unspecified
C0158302|T047|AB|726.10|ICD9CM|Rotator cuff synd NOS|Rotator cuff synd NOS
C0158303|T047|AB|726.11|ICD9CM|Calcif tendinitis shlder|Calcif tendinitis shlder
C0158303|T047|PT|726.11|ICD9CM|Calcifying tendinitis of shoulder|Calcifying tendinitis of shoulder
C0158304|T047|AB|726.12|ICD9CM|Bicipital tenosynovitis|Bicipital tenosynovitis
C0158304|T047|PT|726.12|ICD9CM|Bicipital tenosynovitis|Bicipital tenosynovitis
C3161123|T037|PT|726.13|ICD9CM|Partial tear of rotator cuff|Partial tear of rotator cuff
C3161123|T037|AB|726.13|ICD9CM|Partial tear rotatr cuff|Partial tear rotatr cuff
C0158305|T047|PT|726.19|ICD9CM|Other specified disorders of bursae and tendons in shoulder region|Other specified disorders of bursae and tendons in shoulder region
C0158305|T047|AB|726.19|ICD9CM|Rotator cuff dis NEC|Rotator cuff dis NEC
C0869438|T047|PT|726.2|ICD9CM|Other affections of shoulder region, not elsewhere classified|Other affections of shoulder region, not elsewhere classified
C0869438|T047|AB|726.2|ICD9CM|Shoulder region dis NEC|Shoulder region dis NEC
C0158307|T046|HT|726.3|ICD9CM|Enthesopathy of elbow region|Enthesopathy of elbow region
C0158307|T046|AB|726.30|ICD9CM|Elbow enthesopathy NOS|Elbow enthesopathy NOS
C0158307|T046|PT|726.30|ICD9CM|Enthesopathy of elbow, unspecified|Enthesopathy of elbow, unspecified
C0158309|T020|AB|726.31|ICD9CM|Medial epicondylitis|Medial epicondylitis
C0158309|T020|PT|726.31|ICD9CM|Medial epicondylitis|Medial epicondylitis
C0039516|T047|AB|726.32|ICD9CM|Lateral epicondylitis|Lateral epicondylitis
C0039516|T047|PT|726.32|ICD9CM|Lateral epicondylitis|Lateral epicondylitis
C0263962|T047|AB|726.33|ICD9CM|Olecranon bursitis|Olecranon bursitis
C0263962|T047|PT|726.33|ICD9CM|Olecranon bursitis|Olecranon bursitis
C0158310|T047|AB|726.39|ICD9CM|Elbow enthesopathy NEC|Elbow enthesopathy NEC
C0158310|T047|PT|726.39|ICD9CM|Other enthesopathy of elbow region|Other enthesopathy of elbow region
C0158311|T047|AB|726.4|ICD9CM|Enthesopathy of wrist|Enthesopathy of wrist
C0158311|T047|PT|726.4|ICD9CM|Enthesopathy of wrist and carpus|Enthesopathy of wrist and carpus
C0158312|T047|AB|726.5|ICD9CM|Enthesopathy of hip|Enthesopathy of hip
C0158312|T047|PT|726.5|ICD9CM|Enthesopathy of hip region|Enthesopathy of hip region
C0158313|T047|HT|726.6|ICD9CM|Enthesopathy of knee|Enthesopathy of knee
C0158313|T047|AB|726.60|ICD9CM|Enthesopathy of knee NOS|Enthesopathy of knee NOS
C0158313|T047|PT|726.60|ICD9CM|Enthesopathy of knee, unspecified|Enthesopathy of knee, unspecified
C0158314|T047|AB|726.61|ICD9CM|Pes anserinus tendinitis|Pes anserinus tendinitis
C0158314|T047|PT|726.61|ICD9CM|Pes anserinus tendinitis or bursitis|Pes anserinus tendinitis or bursitis
C0158315|T047|AB|726.62|ICD9CM|Tibial coll lig bursitis|Tibial coll lig bursitis
C0158315|T047|PT|726.62|ICD9CM|Tibial collateral ligament bursitis|Tibial collateral ligament bursitis
C0158316|T047|AB|726.63|ICD9CM|Fibula coll lig bursitis|Fibula coll lig bursitis
C0158316|T047|PT|726.63|ICD9CM|Fibular collateral ligament bursitis|Fibular collateral ligament bursitis
C0158317|T047|AB|726.64|ICD9CM|Patellar tendinitis|Patellar tendinitis
C0158317|T047|PT|726.64|ICD9CM|Patellar tendinitis|Patellar tendinitis
C0851258|T047|AB|726.65|ICD9CM|Prepatellar bursitis|Prepatellar bursitis
C0851258|T047|PT|726.65|ICD9CM|Prepatellar bursitis|Prepatellar bursitis
C0158318|T047|AB|726.69|ICD9CM|Enthesopathy of knee NEC|Enthesopathy of knee NEC
C0158318|T047|PT|726.69|ICD9CM|Other enthesopathy of knee|Other enthesopathy of knee
C0158319|T047|HT|726.7|ICD9CM|Enthesopathy of ankle and tarsus|Enthesopathy of ankle and tarsus
C0158319|T047|AB|726.70|ICD9CM|Ankle enthesopathy NOS|Ankle enthesopathy NOS
C0158319|T047|PT|726.70|ICD9CM|Enthesopathy of ankle and tarsus, unspecified|Enthesopathy of ankle and tarsus, unspecified
C0263933|T047|PT|726.71|ICD9CM|Achilles bursitis or tendinitis|Achilles bursitis or tendinitis
C0263933|T047|AB|726.71|ICD9CM|Achilles tendinitis|Achilles tendinitis
C0158321|T047|AB|726.72|ICD9CM|Tibialis tendinitis|Tibialis tendinitis
C0158321|T047|PT|726.72|ICD9CM|Tibialis tendinitis|Tibialis tendinitis
C0158322|T047|AB|726.73|ICD9CM|Calcaneal spur|Calcaneal spur
C0158322|T047|PT|726.73|ICD9CM|Calcaneal spur|Calcaneal spur
C0158323|T047|AB|726.79|ICD9CM|Ankle enthesopathy NEC|Ankle enthesopathy NEC
C0158323|T047|PT|726.79|ICD9CM|Other enthesopathy of ankle and tarsus|Other enthesopathy of ankle and tarsus
C0158324|T047|PT|726.8|ICD9CM|Other peripheral enthesopathies|Other peripheral enthesopathies
C0158324|T047|AB|726.8|ICD9CM|Periph enthesopathy NEC|Periph enthesopathy NEC
C0242490|T047|HT|726.9|ICD9CM|Unspecified enthesopathy|Unspecified enthesopathy
C0242490|T047|PT|726.90|ICD9CM|Enthesopathy of unspecified site|Enthesopathy of unspecified site
C0242490|T047|AB|726.90|ICD9CM|Enthesopathy, site NOS|Enthesopathy, site NOS
C1442903|T047|PT|726.91|ICD9CM|Exostosis of unspecified site|Exostosis of unspecified site
C1442903|T047|AB|726.91|ICD9CM|Exostosis, site NOS|Exostosis, site NOS
C0158326|T047|HT|727|ICD9CM|Other disorders of synovium, tendon, and bursa|Other disorders of synovium, tendon, and bursa
C0039104|T047|HT|727.0|ICD9CM|Synovitis and tenosynovitis|Synovitis and tenosynovitis
C0039104|T047|PT|727.00|ICD9CM|Synovitis and tenosynovitis, unspecified|Synovitis and tenosynovitis, unspecified
C0039104|T047|AB|727.00|ICD9CM|Synovitis NOS|Synovitis NOS
C0158327|T047|PT|727.01|ICD9CM|Synovitis and tenosynovitis in diseases classified elsewhere|Synovitis and tenosynovitis in diseases classified elsewhere
C0158327|T047|AB|727.01|ICD9CM|Synovitis in oth dis|Synovitis in oth dis
C1318543|T191|PT|727.02|ICD9CM|Giant cell tumor of tendon sheath|Giant cell tumor of tendon sheath
C1318543|T191|AB|727.02|ICD9CM|Giant cell tumor tendon|Giant cell tumor tendon
C3887597|T020|AB|727.03|ICD9CM|Trigger finger|Trigger finger
C3887597|T020|PT|727.03|ICD9CM|Trigger finger (acquired)|Trigger finger (acquired)
C0149870|T047|AB|727.04|ICD9CM|Radial styloid tenosynov|Radial styloid tenosynov
C0149870|T047|PT|727.04|ICD9CM|Radial styloid tenosynovitis|Radial styloid tenosynovitis
C2004376|T047|PT|727.05|ICD9CM|Other tenosynovitis of hand and wrist|Other tenosynovitis of hand and wrist
C2004376|T047|AB|727.05|ICD9CM|Tenosynov hand/wrist NEC|Tenosynov hand/wrist NEC
C0158331|T047|AB|727.06|ICD9CM|Tenosynovitis foot/ankle|Tenosynovitis foot/ankle
C0158331|T047|PT|727.06|ICD9CM|Tenosynovitis of foot and ankle|Tenosynovitis of foot and ankle
C0029856|T047|PT|727.09|ICD9CM|Other synovitis and tenosynovitis|Other synovitis and tenosynovitis
C0029856|T047|AB|727.09|ICD9CM|Synovitis NEC|Synovitis NEC
C0006386|T020|AB|727.1|ICD9CM|Bunion|Bunion
C0006386|T020|PT|727.1|ICD9CM|Bunion|Bunion
C0158332|T047|AB|727.2|ICD9CM|Occupational bursitis|Occupational bursitis
C0158332|T047|PT|727.2|ICD9CM|Specific bursitides often of occupational origin|Specific bursitides often of occupational origin
C0029528|T047|AB|727.3|ICD9CM|Bursitis NEC|Bursitis NEC
C0029528|T047|PT|727.3|ICD9CM|Other bursitis|Other bursitis
C0349693|T047|HT|727.4|ICD9CM|Ganglion and cyst of synovium, tendon, and bursa|Ganglion and cyst of synovium, tendon, and bursa
C0085648|T047|AB|727.40|ICD9CM|Synovial cyst NOS|Synovial cyst NOS
C0085648|T047|PT|727.40|ICD9CM|Synovial cyst, unspecified|Synovial cyst, unspecified
C0158334|T047|AB|727.41|ICD9CM|Ganglion of joint|Ganglion of joint
C0158334|T047|PT|727.41|ICD9CM|Ganglion of joint|Ganglion of joint
C0158335|T020|AB|727.42|ICD9CM|Ganglion of tendon|Ganglion of tendon
C0158335|T020|PT|727.42|ICD9CM|Ganglion of tendon sheath|Ganglion of tendon sheath
C1258666|T047|AB|727.43|ICD9CM|Ganglion NOS|Ganglion NOS
C1258666|T047|PT|727.43|ICD9CM|Ganglion, unspecified|Ganglion, unspecified
C0158336|T047|AB|727.49|ICD9CM|Bursal cyst NEC|Bursal cyst NEC
C0158336|T047|PT|727.49|ICD9CM|Other ganglion and cyst of synovium, tendon, and bursa|Other ganglion and cyst of synovium, tendon, and bursa
C0158337|T046|HT|727.5|ICD9CM|Rupture of synovium|Rupture of synovium
C0158337|T046|AB|727.50|ICD9CM|Rupture of synovium NOS|Rupture of synovium NOS
C0158337|T046|PT|727.50|ICD9CM|Rupture of synovium, unspecified|Rupture of synovium, unspecified
C0032650|T020|AB|727.51|ICD9CM|Popliteal synovial cyst|Popliteal synovial cyst
C0032650|T020|PT|727.51|ICD9CM|Synovial cyst of popliteal space|Synovial cyst of popliteal space
C0158338|T047|PT|727.59|ICD9CM|Other rupture of synovium|Other rupture of synovium
C0158338|T047|AB|727.59|ICD9CM|Rupture of synovium NEC|Rupture of synovium NEC
C0158339|T047|HT|727.6|ICD9CM|Rupture of tendon, nontraumatic|Rupture of tendon, nontraumatic
C0158339|T047|AB|727.60|ICD9CM|Nontraum tendon rupt NOS|Nontraum tendon rupt NOS
C0158339|T047|PT|727.60|ICD9CM|Nontraumatic rupture of unspecified tendon|Nontraumatic rupture of unspecified tendon
C0410017|T037|PT|727.61|ICD9CM|Complete rupture of rotator cuff|Complete rupture of rotator cuff
C0410017|T037|AB|727.61|ICD9CM|Rotator cuff rupture|Rotator cuff rupture
C0158342|T037|AB|727.62|ICD9CM|Biceps tendon rupture|Biceps tendon rupture
C0158342|T037|PT|727.62|ICD9CM|Nontraumatic rupture of tendons of biceps (long head)|Nontraumatic rupture of tendons of biceps (long head)
C4076694|T046|PT|727.63|ICD9CM|Nontraumatic rupture of extensor tendons of hand and wrist|Nontraumatic rupture of extensor tendons of hand and wrist
C4076694|T046|AB|727.63|ICD9CM|Rupt exten tendon hand|Rupt exten tendon hand
C0158344|T047|PT|727.64|ICD9CM|Nontraumatic rupture of flexor tendons of hand and wrist|Nontraumatic rupture of flexor tendons of hand and wrist
C0158344|T047|AB|727.64|ICD9CM|Rupt flexor tendon hand|Rupt flexor tendon hand
C0158345|T037|PT|727.65|ICD9CM|Nontraumatic rupture of quadriceps tendon|Nontraumatic rupture of quadriceps tendon
C0158345|T037|AB|727.65|ICD9CM|Rupture quadricep tendon|Rupture quadricep tendon
C0158346|T037|PT|727.66|ICD9CM|Nontraumatic rupture of patellar tendon|Nontraumatic rupture of patellar tendon
C0158346|T037|AB|727.66|ICD9CM|Rupture patellar tendon|Rupture patellar tendon
C0158347|T037|PT|727.67|ICD9CM|Nontraumatic rupture of achilles tendon|Nontraumatic rupture of achilles tendon
C0158347|T037|AB|727.67|ICD9CM|Rupture achilles tendon|Rupture achilles tendon
C0158348|T047|PT|727.68|ICD9CM|Nontraumatic rupture of other tendons of foot and ankle|Nontraumatic rupture of other tendons of foot and ankle
C0158348|T047|AB|727.68|ICD9CM|Rupture tendon foot NEC|Rupture tendon foot NEC
C0158349|T047|AB|727.69|ICD9CM|Nontraum tendon rupt NEC|Nontraum tendon rupt NEC
C0158349|T047|PT|727.69|ICD9CM|Nontraumatic rupture of other tendon|Nontraumatic rupture of other tendon
C0158326|T047|HT|727.8|ICD9CM|Other disorders of synovium, tendon, and bursa|Other disorders of synovium, tendon, and bursa
C0158350|T046|AB|727.81|ICD9CM|Contracture of tendon|Contracture of tendon
C0158350|T046|PT|727.81|ICD9CM|Contracture of tendon (sheath)|Contracture of tendon (sheath)
C0006690|T033|AB|727.82|ICD9CM|Calcium deposit tendon|Calcium deposit tendon
C0006690|T033|PT|727.82|ICD9CM|Calcium deposits in tendon and bursa|Calcium deposits in tendon and bursa
C0878705|T047|AB|727.83|ICD9CM|Plica syndrome|Plica syndrome
C0878705|T047|PT|727.83|ICD9CM|Plica syndrome|Plica syndrome
C0158326|T047|PT|727.89|ICD9CM|Other disorders of synovium, tendon, and bursa|Other disorders of synovium, tendon, and bursa
C0158326|T047|AB|727.89|ICD9CM|Synov/tend/bursa dis NEC|Synov/tend/bursa dis NEC
C0158351|T047|AB|727.9|ICD9CM|Synov/tend/bursa dis NOS|Synov/tend/bursa dis NOS
C0158351|T047|PT|727.9|ICD9CM|Unspecified disorder of synovium, tendon, and bursa|Unspecified disorder of synovium, tendon, and bursa
C0158352|T047|HT|728|ICD9CM|Disorders of muscle, ligament, and fascia|Disorders of muscle, ligament, and fascia
C0158353|T047|AB|728.0|ICD9CM|Infective myositis|Infective myositis
C0158353|T047|PT|728.0|ICD9CM|Infective myositis|Infective myositis
C0343251|T047|HT|728.1|ICD9CM|Muscular calcification and ossification|Muscular calcification and ossification
C0158355|T047|PT|728.10|ICD9CM|Calcification and ossification, unspecified|Calcification and ossification, unspecified
C0158355|T047|AB|728.10|ICD9CM|Muscular calcificat NOS|Muscular calcificat NOS
C0016037|T047|AB|728.11|ICD9CM|Prog myositis ossificans|Prog myositis ossificans
C0016037|T047|PT|728.11|ICD9CM|Progressive myositis ossificans|Progressive myositis ossificans
C0040798|T047|AB|728.12|ICD9CM|Traum myositis ossifican|Traum myositis ossifican
C0040798|T047|PT|728.12|ICD9CM|Traumatic myositis ossificans|Traumatic myositis ossificans
C0158357|T046|AB|728.13|ICD9CM|Postop heterotopic calc|Postop heterotopic calc
C0158357|T046|PT|728.13|ICD9CM|Postoperative heterotopic calcification|Postoperative heterotopic calcification
C0158358|T047|AB|728.19|ICD9CM|Muscular calcificat NEC|Muscular calcificat NEC
C0158358|T047|PT|728.19|ICD9CM|Other muscular calcification and ossification|Other muscular calcification and ossification
C0868752|T046|AB|728.2|ICD9CM|Musc disuse atrophy NEC|Musc disuse atrophy NEC
C0868752|T046|PT|728.2|ICD9CM|Muscular wasting and disuse atrophy, not elsewhere classified|Muscular wasting and disuse atrophy, not elsewhere classified
C0029741|T047|AB|728.3|ICD9CM|Muscle disorders NEC|Muscle disorders NEC
C0029741|T047|PT|728.3|ICD9CM|Other specific muscle disorders|Other specific muscle disorders
C0158359|T046|AB|728.4|ICD9CM|Laxity of ligament|Laxity of ligament
C0158359|T046|PT|728.4|ICD9CM|Laxity of ligament|Laxity of ligament
C0152093|T047|AB|728.5|ICD9CM|Hypermobility syndrome|Hypermobility syndrome
C0152093|T047|PT|728.5|ICD9CM|Hypermobility syndrome|Hypermobility syndrome
C0013312|T047|AB|728.6|ICD9CM|Contracted palmar fascia|Contracted palmar fascia
C0013312|T047|PT|728.6|ICD9CM|Contracture of palmar fascia|Contracture of palmar fascia
C0079954|T047|HT|728.7|ICD9CM|Other fibromatoses of muscle, ligament, and fascia|Other fibromatoses of muscle, ligament, and fascia
C0158360|T047|PT|728.71|ICD9CM|Plantar fascial fibromatosis|Plantar fascial fibromatosis
C0158360|T047|AB|728.71|ICD9CM|Plantar fibromatosis|Plantar fibromatosis
C0079954|T047|AB|728.79|ICD9CM|Fibromatoses NEC|Fibromatoses NEC
C0079954|T047|PT|728.79|ICD9CM|Other fibromatoses of muscle, ligament, and fascia|Other fibromatoses of muscle, ligament, and fascia
C0158361|T047|HT|728.8|ICD9CM|Other disorders of muscle, ligament, and fascia|Other disorders of muscle, ligament, and fascia
C0158362|T047|AB|728.81|ICD9CM|Interstitial myositis|Interstitial myositis
C0158362|T047|PT|728.81|ICD9CM|Interstitial myositis|Interstitial myositis
C0016545|T047|AB|728.82|ICD9CM|FB granuloma of muscle|FB granuloma of muscle
C0016545|T047|PT|728.82|ICD9CM|Foreign body granuloma of muscle|Foreign body granuloma of muscle
C0158363|T037|AB|728.83|ICD9CM|Nontraum muscle rupture|Nontraum muscle rupture
C0158363|T037|PT|728.83|ICD9CM|Rupture of muscle, nontraumatic|Rupture of muscle, nontraumatic
C0158364|T190|AB|728.84|ICD9CM|Diastasis of muscle|Diastasis of muscle
C0158364|T190|PT|728.84|ICD9CM|Diastasis of muscle|Diastasis of muscle
C0037763|T184|AB|728.85|ICD9CM|Spasm of muscle|Spasm of muscle
C0037763|T184|PT|728.85|ICD9CM|Spasm of muscle|Spasm of muscle
C0238124|T047|AB|728.86|ICD9CM|Necrotizing fasciitis|Necrotizing fasciitis
C0238124|T047|PT|728.86|ICD9CM|Necrotizing fasciitis|Necrotizing fasciitis
C0746674|T184|PT|728.87|ICD9CM|Muscle weakness (generalized)|Muscle weakness (generalized)
C0746674|T184|AB|728.87|ICD9CM|Muscle weakness-general|Muscle weakness-general
C0035410|T046|AB|728.88|ICD9CM|Rhabdomyolysis|Rhabdomyolysis
C0035410|T046|PT|728.88|ICD9CM|Rhabdomyolysis|Rhabdomyolysis
C0158361|T047|AB|728.89|ICD9CM|Muscle/ligament dis NEC|Muscle/ligament dis NEC
C0158361|T047|PT|728.89|ICD9CM|Other disorders of muscle, ligament, and fascia|Other disorders of muscle, ligament, and fascia
C0158352|T047|AB|728.9|ICD9CM|Muscle/ligament dis NOS|Muscle/ligament dis NOS
C0158352|T047|PT|728.9|ICD9CM|Unspecified disorder of muscle, ligament, and fascia|Unspecified disorder of muscle, ligament, and fascia
C0158370|T047|HT|729|ICD9CM|Other disorders of soft tissues|Other disorders of soft tissues
C0035445|T047|AB|729.0|ICD9CM|Rheumatism NOS|Rheumatism NOS
C0035445|T047|PT|729.0|ICD9CM|Rheumatism, unspecified and fibrositis|Rheumatism, unspecified and fibrositis
C0026893|T047|AB|729.1|ICD9CM|Myalgia and myositis NOS|Myalgia and myositis NOS
C0026893|T047|PT|729.1|ICD9CM|Myalgia and myositis, unspecified|Myalgia and myositis, unspecified
C0347894|T047|PT|729.2|ICD9CM|Neuralgia, neuritis, and radiculitis, unspecified|Neuralgia, neuritis, and radiculitis, unspecified
C0347894|T047|AB|729.2|ICD9CM|Neuralgia/neuritis NOS|Neuralgia/neuritis NOS
C0030326|T047|HT|729.3|ICD9CM|Panniculitis, unspecified|Panniculitis, unspecified
C0030326|T047|AB|729.30|ICD9CM|Panniculitis, unsp site|Panniculitis, unsp site
C0030326|T047|PT|729.30|ICD9CM|Panniculitis, unspecified site|Panniculitis, unspecified site
C0158366|T033|AB|729.31|ICD9CM|Hypertrophy of fat pad|Hypertrophy of fat pad
C0158366|T033|PT|729.31|ICD9CM|Hypertrophy of fat pad, knee|Hypertrophy of fat pad, knee
C0158367|T047|PT|729.39|ICD9CM|Panniculitis, other site|Panniculitis, other site
C0158367|T047|AB|729.39|ICD9CM|Panniculitis, site NEC|Panniculitis, site NEC
C0015645|T047|AB|729.4|ICD9CM|Fasciitis NOS|Fasciitis NOS
C0015645|T047|PT|729.4|ICD9CM|Fasciitis, unspecified|Fasciitis, unspecified
C0030196|T184|AB|729.5|ICD9CM|Pain in limb|Pain in limb
C0030196|T184|PT|729.5|ICD9CM|Pain in limb|Pain in limb
C0158368|T020|AB|729.6|ICD9CM|Old FB in soft tissue|Old FB in soft tissue
C0158368|T020|PT|729.6|ICD9CM|Residual foreign body in soft tissue|Residual foreign body in soft tissue
C1719623|T047|HT|729.7|ICD9CM|Nontraumatic compartment syndrome|Nontraumatic compartment syndrome
C1719618|T047|AB|729.71|ICD9CM|Nontraum comp syn-up ext|Nontraum comp syn-up ext
C1719618|T047|PT|729.71|ICD9CM|Nontraumatic compartment syndrome of upper extremity|Nontraumatic compartment syndrome of upper extremity
C1719620|T047|AB|729.72|ICD9CM|Nontraum comp syn-low ex|Nontraum comp syn-low ex
C1719620|T047|PT|729.72|ICD9CM|Nontraumatic compartment syndrome of lower extremity|Nontraumatic compartment syndrome of lower extremity
C1719621|T047|AB|729.73|ICD9CM|Nontrauma comp syn-abd|Nontrauma comp syn-abd
C1719621|T047|PT|729.73|ICD9CM|Nontraumatic compartment syndrome of abdomen|Nontraumatic compartment syndrome of abdomen
C1719622|T047|AB|729.79|ICD9CM|Nontrauma comp syn NEC|Nontrauma comp syn NEC
C1719622|T047|PT|729.79|ICD9CM|Nontraumatic compartment syndrome of other sites|Nontraumatic compartment syndrome of other sites
C0029669|T184|HT|729.8|ICD9CM|Other musculoskeletal symptoms referable to limbs|Other musculoskeletal symptoms referable to limbs
C0158369|T184|AB|729.81|ICD9CM|Swelling of limb|Swelling of limb
C0158369|T184|PT|729.81|ICD9CM|Swelling of limb|Swelling of limb
C0010263|T184|AB|729.82|ICD9CM|Cramp in limb|Cramp in limb
C0010263|T184|PT|729.82|ICD9CM|Cramp of limb|Cramp of limb
C0029669|T184|AB|729.89|ICD9CM|Muscskel sympt limb NEC|Muscskel sympt limb NEC
C0029669|T184|PT|729.89|ICD9CM|Other musculoskeletal symptoms referable to limbs|Other musculoskeletal symptoms referable to limbs
C0158370|T047|HT|729.9|ICD9CM|Other and unspecified disorders of soft tissue|Other and unspecified disorders of soft tissue
C0263978|T047|PT|729.90|ICD9CM|Disorders of soft tissue, unspecified|Disorders of soft tissue, unspecified
C0263978|T047|AB|729.90|ICD9CM|Soft tissue disord NOS|Soft tissue disord NOS
C2349647|T047|AB|729.91|ICD9CM|Post-traumatic seroma|Post-traumatic seroma
C2349647|T047|PT|729.91|ICD9CM|Post-traumatic seroma|Post-traumatic seroma
C2349648|T047|AB|729.92|ICD9CM|Nontrauma hema soft tiss|Nontrauma hema soft tiss
C2349648|T047|PT|729.92|ICD9CM|Nontraumatic hematoma of soft tissue|Nontraumatic hematoma of soft tissue
C0158370|T047|PT|729.99|ICD9CM|Other disorders of soft tissue|Other disorders of soft tissue
C0158370|T047|AB|729.99|ICD9CM|Soft tissue disorder NEC|Soft tissue disorder NEC
C0195720|T033|AB|73.3|ICD9CM|Failed forceps|Failed forceps
C0195720|T033|PT|73.3|ICD9CM|Failed forceps|Failed forceps
C0343139|T047|HT|730|ICD9CM|Osteomyelitis, periostitis, and other infections involving bone|Osteomyelitis, periostitis, and other infections involving bone
C0178306|T047|HT|730-739.99|ICD9CM|OSTEOPATHIES, CHONDROPATHIES, AND ACQUIRED MUSCULOSKELETAL DEFORMITIES|OSTEOPATHIES, CHONDROPATHIES, AND ACQUIRED MUSCULOSKELETAL DEFORMITIES
C0158371|T047|HT|730.0|ICD9CM|Acute osteomyelitis|Acute osteomyelitis
C0158371|T047|AB|730.00|ICD9CM|Ac osteomyelitis-unspec|Ac osteomyelitis-unspec
C0158371|T047|PT|730.00|ICD9CM|Acute osteomyelitis, site unspecified|Acute osteomyelitis, site unspecified
C0158372|T047|AB|730.01|ICD9CM|Ac osteomyelitis-shlder|Ac osteomyelitis-shlder
C0158372|T047|PT|730.01|ICD9CM|Acute osteomyelitis, shoulder region|Acute osteomyelitis, shoulder region
C0158373|T047|AB|730.02|ICD9CM|Ac osteomyelitis-up/arm|Ac osteomyelitis-up/arm
C0158373|T047|PT|730.02|ICD9CM|Acute osteomyelitis, upper arm|Acute osteomyelitis, upper arm
C0158374|T047|AB|730.03|ICD9CM|Ac osteomyelitis-forearm|Ac osteomyelitis-forearm
C0158374|T047|PT|730.03|ICD9CM|Acute osteomyelitis, forearm|Acute osteomyelitis, forearm
C0158375|T047|AB|730.04|ICD9CM|Ac osteomyelitis-hand|Ac osteomyelitis-hand
C0158375|T047|PT|730.04|ICD9CM|Acute osteomyelitis, hand|Acute osteomyelitis, hand
C1963552|T047|AB|730.05|ICD9CM|Ac osteomyelitis-pelvis|Ac osteomyelitis-pelvis
C1963552|T047|PT|730.05|ICD9CM|Acute osteomyelitis, pelvic region and thigh|Acute osteomyelitis, pelvic region and thigh
C0158377|T047|AB|730.06|ICD9CM|Ac osteomyelitis-l/leg|Ac osteomyelitis-l/leg
C0158377|T047|PT|730.06|ICD9CM|Acute osteomyelitis, lower leg|Acute osteomyelitis, lower leg
C0264039|T047|AB|730.07|ICD9CM|Ac osteomyelitis-ankle|Ac osteomyelitis-ankle
C0264039|T047|PT|730.07|ICD9CM|Acute osteomyelitis, ankle and foot|Acute osteomyelitis, ankle and foot
C0410385|T047|AB|730.08|ICD9CM|Ac osteomyelitis NEC|Ac osteomyelitis NEC
C0410385|T047|PT|730.08|ICD9CM|Acute osteomyelitis, other specified sites|Acute osteomyelitis, other specified sites
C0158380|T047|AB|730.09|ICD9CM|Ac osteomyelitis-mult|Ac osteomyelitis-mult
C0158380|T047|PT|730.09|ICD9CM|Acute osteomyelitis, multiple sites|Acute osteomyelitis, multiple sites
C0008707|T047|HT|730.1|ICD9CM|Chronic osteomyelitis|Chronic osteomyelitis
C0008707|T047|AB|730.10|ICD9CM|Chr osteomyelitis-unsp|Chr osteomyelitis-unsp
C0008707|T047|PT|730.10|ICD9CM|Chronic osteomyelitis, site unspecified|Chronic osteomyelitis, site unspecified
C0158381|T047|AB|730.11|ICD9CM|Chr osteomyelit-shlder|Chr osteomyelit-shlder
C0158381|T047|PT|730.11|ICD9CM|Chronic osteomyelitis, shoulder region|Chronic osteomyelitis, shoulder region
C0158382|T047|AB|730.12|ICD9CM|Chr osteomyelit-up/arm|Chr osteomyelit-up/arm
C0158382|T047|PT|730.12|ICD9CM|Chronic osteomyelitis, upper arm|Chronic osteomyelitis, upper arm
C0158383|T047|AB|730.13|ICD9CM|Chr osteomyelit-forearm|Chr osteomyelit-forearm
C0158383|T047|PT|730.13|ICD9CM|Chronic osteomyelitis, forearm|Chronic osteomyelitis, forearm
C0158384|T047|AB|730.14|ICD9CM|Chr osteomyelit-hand|Chr osteomyelit-hand
C0158384|T047|PT|730.14|ICD9CM|Chronic osteomyelitis, hand|Chronic osteomyelitis, hand
C0410420|T047|AB|730.15|ICD9CM|Chr osteomyelit-pelvis|Chr osteomyelit-pelvis
C0410420|T047|PT|730.15|ICD9CM|Chronic osteomyelitis, pelvic region and thigh|Chronic osteomyelitis, pelvic region and thigh
C0158386|T047|AB|730.16|ICD9CM|Chr osteomyelit-l/leg|Chr osteomyelit-l/leg
C0158386|T047|PT|730.16|ICD9CM|Chronic osteomyelitis, lower leg|Chronic osteomyelitis, lower leg
C0264049|T047|AB|730.17|ICD9CM|Chr osteomyelit-ankle|Chr osteomyelit-ankle
C0264049|T047|PT|730.17|ICD9CM|Chronic osteomyelitis, ankle and foot|Chronic osteomyelitis, ankle and foot
C0410417|T047|AB|730.18|ICD9CM|Chr osteomyelit NEC|Chr osteomyelit NEC
C0410417|T047|PT|730.18|ICD9CM|Chronic osteomyelitis, other specified sites|Chronic osteomyelitis, other specified sites
C0264051|T047|AB|730.19|ICD9CM|Chr osteomyelit-mult|Chr osteomyelit-mult
C0264051|T047|PT|730.19|ICD9CM|Chronic osteomyelitis, multiple sites|Chronic osteomyelitis, multiple sites
C0029443|T047|HT|730.2|ICD9CM|Unspecified osteomyelitis|Unspecified osteomyelitis
C0029443|T047|AB|730.20|ICD9CM|Osteomyelitis NOS-unspec|Osteomyelitis NOS-unspec
C0029443|T047|PT|730.20|ICD9CM|Unspecified osteomyelitis, site unspecified|Unspecified osteomyelitis, site unspecified
C0264022|T047|AB|730.21|ICD9CM|Osteomyelitis NOS-shlder|Osteomyelitis NOS-shlder
C0264022|T047|PT|730.21|ICD9CM|Unspecified osteomyelitis, shoulder region|Unspecified osteomyelitis, shoulder region
C0264023|T047|AB|730.22|ICD9CM|Osteomyelitis NOS-up/arm|Osteomyelitis NOS-up/arm
C0264023|T047|PT|730.22|ICD9CM|Unspecified osteomyelitis, upper arm|Unspecified osteomyelitis, upper arm
C0264024|T047|AB|730.23|ICD9CM|Osteomyelit NOS-forearm|Osteomyelit NOS-forearm
C0264024|T047|PT|730.23|ICD9CM|Unspecified osteomyelitis, forearm|Unspecified osteomyelitis, forearm
C0264025|T047|AB|730.24|ICD9CM|Osteomyelitis NOS-hand|Osteomyelitis NOS-hand
C0264025|T047|PT|730.24|ICD9CM|Unspecified osteomyelitis, hand|Unspecified osteomyelitis, hand
C0158434|T047|AB|730.25|ICD9CM|Osteomyelitis NOS-pelvis|Osteomyelitis NOS-pelvis
C0158434|T047|PT|730.25|ICD9CM|Unspecified osteomyelitis, pelvic region and thigh|Unspecified osteomyelitis, pelvic region and thigh
C0158395|T047|AB|730.26|ICD9CM|Osteomyelitis NOS-l/leg|Osteomyelitis NOS-l/leg
C0158395|T047|PT|730.26|ICD9CM|Unspecified osteomyelitis, lower leg|Unspecified osteomyelitis, lower leg
C0158396|T047|AB|730.27|ICD9CM|Osteomyelitis NOS-ankle|Osteomyelitis NOS-ankle
C0158396|T047|PT|730.27|ICD9CM|Unspecified osteomyelitis, ankle and foot|Unspecified osteomyelitis, ankle and foot
C0410376|T047|AB|730.28|ICD9CM|Osteomyelit NOS-oth site|Osteomyelit NOS-oth site
C0410376|T047|PT|730.28|ICD9CM|Unspecified osteomyelitis, other specified sites|Unspecified osteomyelitis, other specified sites
C0264031|T047|AB|730.29|ICD9CM|Osteomyelitis NOS-mult|Osteomyelitis NOS-mult
C0264031|T047|PT|730.29|ICD9CM|Unspecified osteomyelitis, multiple sites|Unspecified osteomyelitis, multiple sites
C0264069|T047|HT|730.3|ICD9CM|Periostitis without mention of osteomyelitis|Periostitis without mention of osteomyelitis
C0410437|T047|AB|730.30|ICD9CM|Periostitis-unspec|Periostitis-unspec
C0410437|T047|PT|730.30|ICD9CM|Periostitis, without mention of osteomyelitis, site unspecified|Periostitis, without mention of osteomyelitis, site unspecified
C0410436|T047|AB|730.31|ICD9CM|Periostitis-shlder|Periostitis-shlder
C0410436|T047|PT|730.31|ICD9CM|Periostitis, without mention of osteomyelitis, shoulder region|Periostitis, without mention of osteomyelitis, shoulder region
C0158401|T047|AB|730.32|ICD9CM|Periostitis-up/arm|Periostitis-up/arm
C0158401|T047|PT|730.32|ICD9CM|Periostitis, without mention of osteomyelitis, upper arm|Periostitis, without mention of osteomyelitis, upper arm
C0158402|T047|AB|730.33|ICD9CM|Periostitis-forearm|Periostitis-forearm
C0158402|T047|PT|730.33|ICD9CM|Periostitis, without mention of osteomyelitis, forearm|Periostitis, without mention of osteomyelitis, forearm
C0158403|T047|AB|730.34|ICD9CM|Periostitis-hand|Periostitis-hand
C0158403|T047|PT|730.34|ICD9CM|Periostitis, without mention of osteomyelitis, hand|Periostitis, without mention of osteomyelitis, hand
C0410435|T047|AB|730.35|ICD9CM|Periostitis-pelvis|Periostitis-pelvis
C0410435|T047|PT|730.35|ICD9CM|Periostitis, without mention of osteomyelitis, pelvic region and thigh|Periostitis, without mention of osteomyelitis, pelvic region and thigh
C0158405|T047|AB|730.36|ICD9CM|Periostitis-l/leg|Periostitis-l/leg
C0158405|T047|PT|730.36|ICD9CM|Periostitis, without mention of osteomyelitis, lower leg|Periostitis, without mention of osteomyelitis, lower leg
C0158406|T047|AB|730.37|ICD9CM|Periostitis-ankle|Periostitis-ankle
C0158406|T047|PT|730.37|ICD9CM|Periostitis, without mention of osteomyelitis, ankle and foot|Periostitis, without mention of osteomyelitis, ankle and foot
C0410434|T047|AB|730.38|ICD9CM|Periostitis NEC|Periostitis NEC
C0410434|T047|PT|730.38|ICD9CM|Periostitis, without mention of osteomyelitis, other specified sites|Periostitis, without mention of osteomyelitis, other specified sites
C0158407|T047|AB|730.39|ICD9CM|Periostitis-mult|Periostitis-mult
C0158407|T047|PT|730.39|ICD9CM|Periostitis, without mention of osteomyelitis, multiple sites|Periostitis, without mention of osteomyelitis, multiple sites
C0158408|T047|HT|730.7|ICD9CM|Osteopathy resulting from poliomyelitis|Osteopathy resulting from poliomyelitis
C0158408|T047|PT|730.70|ICD9CM|Osteopathy resulting from poliomyelitis, site unspecified|Osteopathy resulting from poliomyelitis, site unspecified
C0158408|T047|AB|730.70|ICD9CM|Polio osteopathy-unspec|Polio osteopathy-unspec
C0410326|T047|PT|730.71|ICD9CM|Osteopathy resulting from poliomyelitis, shoulder region|Osteopathy resulting from poliomyelitis, shoulder region
C0410326|T047|AB|730.71|ICD9CM|Polio osteopathy-shlder|Polio osteopathy-shlder
C0410325|T047|PT|730.72|ICD9CM|Osteopathy resulting from poliomyelitis, upper arm|Osteopathy resulting from poliomyelitis, upper arm
C0410325|T047|AB|730.72|ICD9CM|Polio osteopathy-up/arm|Polio osteopathy-up/arm
C0410324|T047|PT|730.73|ICD9CM|Osteopathy resulting from poliomyelitis, forearm|Osteopathy resulting from poliomyelitis, forearm
C0410324|T047|AB|730.73|ICD9CM|Polio osteopathy-forearm|Polio osteopathy-forearm
C0410323|T047|PT|730.74|ICD9CM|Osteopathy resulting from poliomyelitis, hand|Osteopathy resulting from poliomyelitis, hand
C0410323|T047|AB|730.74|ICD9CM|Polio osteopathy-hand|Polio osteopathy-hand
C0410322|T047|PT|730.75|ICD9CM|Osteopathy resulting from poliomyelitis, pelvic region and thigh|Osteopathy resulting from poliomyelitis, pelvic region and thigh
C0410322|T047|AB|730.75|ICD9CM|Polio osteopathy-pelvis|Polio osteopathy-pelvis
C0410321|T047|PT|730.76|ICD9CM|Osteopathy resulting from poliomyelitis, lower leg|Osteopathy resulting from poliomyelitis, lower leg
C0410321|T047|AB|730.76|ICD9CM|Polio osteopathy-l/leg|Polio osteopathy-l/leg
C0410320|T047|PT|730.77|ICD9CM|Osteopathy resulting from poliomyelitis, ankle and foot|Osteopathy resulting from poliomyelitis, ankle and foot
C0410320|T047|AB|730.77|ICD9CM|Polio osteopathy-ankle|Polio osteopathy-ankle
C0410319|T047|PT|730.78|ICD9CM|Osteopathy resulting from poliomyelitis, other specified sites|Osteopathy resulting from poliomyelitis, other specified sites
C0410319|T047|AB|730.78|ICD9CM|Polio osteopathy NEC|Polio osteopathy NEC
C0410318|T047|PT|730.79|ICD9CM|Osteopathy resulting from poliomyelitis, multiple sites|Osteopathy resulting from poliomyelitis, multiple sites
C0410318|T047|AB|730.79|ICD9CM|Polio osteopathy-mult|Polio osteopathy-mult
C0264070|T047|HT|730.8|ICD9CM|Other infections involving bone in disease classified elsewhere|Other infections involving bone in disease classified elsewhere
C0264070|T047|AB|730.80|ICD9CM|Bone infect NEC-unspec|Bone infect NEC-unspec
C0264070|T047|PT|730.80|ICD9CM|Other infections involving bone in diseases classified elsewhere, site unspecified|Other infections involving bone in diseases classified elsewhere, site unspecified
C0158420|T047|AB|730.81|ICD9CM|Bone infect NEC-shlder|Bone infect NEC-shlder
C0158420|T047|PT|730.81|ICD9CM|Other infections involving bone in diseases classified elsewhere, shoulder region|Other infections involving bone in diseases classified elsewhere, shoulder region
C0158421|T047|AB|730.82|ICD9CM|Bone infect NEC-up/arm|Bone infect NEC-up/arm
C0158421|T047|PT|730.82|ICD9CM|Other infections involving bone in diseases classified elsewhere, upper arm|Other infections involving bone in diseases classified elsewhere, upper arm
C0158422|T047|AB|730.83|ICD9CM|Bone infect NEC-forearm|Bone infect NEC-forearm
C0158422|T047|PT|730.83|ICD9CM|Other infections involving bone in diseases classified elsewhere, forearm|Other infections involving bone in diseases classified elsewhere, forearm
C0158423|T047|AB|730.84|ICD9CM|Bone infect NEC-hand|Bone infect NEC-hand
C0158423|T047|PT|730.84|ICD9CM|Other infections involving bone in diseases classified elsewhere, hand|Other infections involving bone in diseases classified elsewhere, hand
C0158424|T047|AB|730.85|ICD9CM|Bone infect NEC-pelvis|Bone infect NEC-pelvis
C0158424|T047|PT|730.85|ICD9CM|Other infections involving bone in diseases classified elsewhere, pelvic region and thigh|Other infections involving bone in diseases classified elsewhere, pelvic region and thigh
C0158425|T047|AB|730.86|ICD9CM|Bone infect NEC-l/leg|Bone infect NEC-l/leg
C0158425|T047|PT|730.86|ICD9CM|Other infections involving bone in diseases classified elsewhere, lower leg|Other infections involving bone in diseases classified elsewhere, lower leg
C0158426|T047|AB|730.87|ICD9CM|Bone infect NEC-ankle|Bone infect NEC-ankle
C0158426|T047|PT|730.87|ICD9CM|Other infections involving bone in diseases classified elsewhere, ankle and foot|Other infections involving bone in diseases classified elsewhere, ankle and foot
C0158427|T047|AB|730.88|ICD9CM|Bone infect NEC-oth site|Bone infect NEC-oth site
C0158427|T047|PT|730.88|ICD9CM|Other infections involving bone in diseases classified elsewhere, other specified sites|Other infections involving bone in diseases classified elsewhere, other specified sites
C0158428|T047|AB|730.89|ICD9CM|Bone infect NEC-mult|Bone infect NEC-mult
C0158428|T047|PT|730.89|ICD9CM|Other infections involving bone in diseases classified elsewhere, multiple sites|Other infections involving bone in diseases classified elsewhere, multiple sites
C2242472|T047|HT|730.9|ICD9CM|Unspecified infection of bone|Unspecified infection of bone
C2242472|T047|AB|730.90|ICD9CM|Bone infec NOS-unsp site|Bone infec NOS-unsp site
C2242472|T047|PT|730.90|ICD9CM|Unspecified infection of bone, site unspecified|Unspecified infection of bone, site unspecified
C0264022|T047|AB|730.91|ICD9CM|Bone infect NOS-shlder|Bone infect NOS-shlder
C0264022|T047|PT|730.91|ICD9CM|Unspecified infection of bone, shoulder region|Unspecified infection of bone, shoulder region
C0264023|T047|AB|730.92|ICD9CM|Bone infect NOS-up/arm|Bone infect NOS-up/arm
C0264023|T047|PT|730.92|ICD9CM|Unspecified infection of bone, upper arm|Unspecified infection of bone, upper arm
C0264024|T047|AB|730.93|ICD9CM|Bone infect NOS-forearm|Bone infect NOS-forearm
C0264024|T047|PT|730.93|ICD9CM|Unspecified infection of bone, forearm|Unspecified infection of bone, forearm
C2242475|T047|AB|730.94|ICD9CM|Bone infect NOS-hand|Bone infect NOS-hand
C2242475|T047|PT|730.94|ICD9CM|Unspecified infection of bone, hand|Unspecified infection of bone, hand
C0158434|T047|AB|730.95|ICD9CM|Bone infect NOS-pelvis|Bone infect NOS-pelvis
C0158434|T047|PT|730.95|ICD9CM|Unspecified infection of bone, pelvic region and thigh|Unspecified infection of bone, pelvic region and thigh
C0264028|T047|AB|730.96|ICD9CM|Bone infect NOS-l/leg|Bone infect NOS-l/leg
C0264028|T047|PT|730.96|ICD9CM|Unspecified infection of bone, lower leg|Unspecified infection of bone, lower leg
C0264029|T047|AB|730.97|ICD9CM|Bone infect NOS-ankle|Bone infect NOS-ankle
C0264029|T047|PT|730.97|ICD9CM|Unspecified infection of bone, ankle and foot|Unspecified infection of bone, ankle and foot
C0158437|T047|AB|730.98|ICD9CM|Bone infect NOS-oth site|Bone infect NOS-oth site
C0158437|T047|PT|730.98|ICD9CM|Unspecified infection of bone, other specified sites|Unspecified infection of bone, other specified sites
C0158438|T047|AB|730.99|ICD9CM|Bone infect NOS-mult|Bone infect NOS-mult
C0158438|T047|PT|730.99|ICD9CM|Unspecified infection of bone, multiple sites|Unspecified infection of bone, multiple sites
C0029402|T047|HT|731|ICD9CM|Osteitis deformans and osteopathies associated with other disorders classified elsewhere|Osteitis deformans and osteopathies associated with other disorders classified elsewhere
C0029403|T047|AB|731.0|ICD9CM|Osteitis deformans NOS|Osteitis deformans NOS
C0029403|T047|PT|731.0|ICD9CM|Osteitis deformans without mention of bone tumor|Osteitis deformans without mention of bone tumor
C0158439|T047|AB|731.1|ICD9CM|Osteitis def in oth dis|Osteitis def in oth dis
C0158439|T047|PT|731.1|ICD9CM|Osteitis deformans in diseases classified elsewhere|Osteitis deformans in diseases classified elsewhere
C0029412|T047|AB|731.2|ICD9CM|Hypertroph osteoarthrop|Hypertroph osteoarthrop
C0029412|T047|PT|731.2|ICD9CM|Hypertrophic pulmonary osteoarthropathy|Hypertrophic pulmonary osteoarthropathy
C1719624|T047|AB|731.3|ICD9CM|Major osseous defects|Major osseous defects
C1719624|T047|PT|731.3|ICD9CM|Major osseous defects|Major osseous defects
C0158440|T047|AB|731.8|ICD9CM|Bone involv in oth dis|Bone involv in oth dis
C0158440|T047|PT|731.8|ICD9CM|Other bone involvement in diseases classified elsewhere|Other bone involvement in diseases classified elsewhere
C0152091|T047|HT|732|ICD9CM|Osteochondropathies|Osteochondropathies
C0036310|T047|AB|732.0|ICD9CM|Juv osteochondros spine|Juv osteochondros spine
C0036310|T047|PT|732.0|ICD9CM|Juvenile osteochondrosis of spine|Juvenile osteochondrosis of spine
C0410502|T047|AB|732.1|ICD9CM|Juv osteochondros pelvis|Juv osteochondros pelvis
C0410502|T047|PT|732.1|ICD9CM|Juvenile osteochondrosis of hip and pelvis|Juvenile osteochondrosis of hip and pelvis
C0158441|T037|AB|732.2|ICD9CM|Femoral epiphysiolysis|Femoral epiphysiolysis
C0158441|T037|PT|732.2|ICD9CM|Nontraumatic slipped upper femoral epiphysis|Nontraumatic slipped upper femoral epiphysis
C0158442|T047|AB|732.3|ICD9CM|Juv osteochondrosis arm|Juv osteochondrosis arm
C0158442|T047|PT|732.3|ICD9CM|Juvenile osteochondrosis of upper extremity|Juvenile osteochondrosis of upper extremity
C1282912|T047|AB|732.4|ICD9CM|Juv osteochondrosis leg|Juv osteochondrosis leg
C1282912|T047|PT|732.4|ICD9CM|Juvenile osteochondrosis of lower extremity, excluding foot|Juvenile osteochondrosis of lower extremity, excluding foot
C0158444|T047|AB|732.5|ICD9CM|Juv osteochondrosis foot|Juv osteochondrosis foot
C0158444|T047|PT|732.5|ICD9CM|Juvenile osteochondrosis of foot|Juvenile osteochondrosis of foot
C0158445|T047|AB|732.6|ICD9CM|Juv osteochondrosis NEC|Juv osteochondrosis NEC
C0158445|T047|PT|732.6|ICD9CM|Other juvenile osteochondrosis|Other juvenile osteochondrosis
C0029421|T047|AB|732.7|ICD9CM|Osteochondrit dissecans|Osteochondrit dissecans
C0029421|T047|PT|732.7|ICD9CM|Osteochondritis dissecans|Osteochondritis dissecans
C0451640|T047|AB|732.8|ICD9CM|Osteochondropathy NEC|Osteochondropathy NEC
C0451640|T047|PT|732.8|ICD9CM|Other specified forms of osteochondropathy|Other specified forms of osteochondropathy
C0152091|T047|AB|732.9|ICD9CM|Osteochondropathy NOS|Osteochondropathy NOS
C0152091|T047|PT|732.9|ICD9CM|Unspecified osteochondropathy|Unspecified osteochondropathy
C0029586|T047|HT|733|ICD9CM|Other disorders of bone and cartilage|Other disorders of bone and cartilage
C0029456|T047|HT|733.0|ICD9CM|Osteoporosis|Osteoporosis
C0029456|T047|AB|733.00|ICD9CM|Osteoporosis NOS|Osteoporosis NOS
C0029456|T047|PT|733.00|ICD9CM|Osteoporosis, unspecified|Osteoporosis, unspecified
C0029459|T047|AB|733.01|ICD9CM|Senile osteoporosis|Senile osteoporosis
C0029459|T047|PT|733.01|ICD9CM|Senile osteoporosis|Senile osteoporosis
C0158447|T047|AB|733.02|ICD9CM|Idiopathic osteoporosis|Idiopathic osteoporosis
C0158447|T047|PT|733.02|ICD9CM|Idiopathic osteoporosis|Idiopathic osteoporosis
C0152256|T047|AB|733.03|ICD9CM|Disuse osteoporosis|Disuse osteoporosis
C0152256|T047|PT|733.03|ICD9CM|Disuse osteoporosis|Disuse osteoporosis
C0029694|T047|AB|733.09|ICD9CM|Osteoporosis NEC|Osteoporosis NEC
C0029694|T047|PT|733.09|ICD9CM|Other osteoporosis|Other osteoporosis
C0016663|T046|HT|733.1|ICD9CM|Pathologic fracture|Pathologic fracture
C0016663|T046|AB|733.10|ICD9CM|Path fx unspecified site|Path fx unspecified site
C0016663|T046|PT|733.10|ICD9CM|Pathologic fracture, unspecified site|Pathologic fracture, unspecified site
C0375504|T046|AB|733.11|ICD9CM|Path fx humerus|Path fx humerus
C0375504|T046|PT|733.11|ICD9CM|Pathologic fracture of humerus|Pathologic fracture of humerus
C0375505|T046|AB|733.12|ICD9CM|Path fx dstl radius ulna|Path fx dstl radius ulna
C0375505|T046|PT|733.12|ICD9CM|Pathologic fracture of distal radius and ulna|Pathologic fracture of distal radius and ulna
C0302491|T046|AB|733.13|ICD9CM|Path fx vertebrae|Path fx vertebrae
C0302491|T046|PT|733.13|ICD9CM|Pathologic fracture of vertebrae|Pathologic fracture of vertebrae
C1443978|T046|AB|733.14|ICD9CM|Path fx neck of femur|Path fx neck of femur
C1443978|T046|PT|733.14|ICD9CM|Pathologic fracture of neck of femur|Pathologic fracture of neck of femur
C0375507|T046|AB|733.15|ICD9CM|Path fx oth spcf prt fmr|Path fx oth spcf prt fmr
C0375507|T046|PT|733.15|ICD9CM|Pathologic fracture of other specified part of femur|Pathologic fracture of other specified part of femur
C0375508|T046|AB|733.16|ICD9CM|Path fx tibia fibula|Path fx tibia fibula
C0375508|T046|PT|733.16|ICD9CM|Pathologic fracture of tibia or fibula|Pathologic fracture of tibia or fibula
C0375509|T046|AB|733.19|ICD9CM|Path fx oth specif site|Path fx oth specif site
C0375509|T046|PT|733.19|ICD9CM|Pathologic fracture of other specified site|Pathologic fracture of other specified site
C0005937|T190|HT|733.2|ICD9CM|Cyst of bone|Cyst of bone
C0005937|T190|PT|733.20|ICD9CM|Cyst of bone (localized), unspecified|Cyst of bone (localized), unspecified
C0005937|T190|AB|733.20|ICD9CM|Cyst of bone NOS|Cyst of bone NOS
C0005937|T190|AB|733.21|ICD9CM|Solitary bone cyst|Solitary bone cyst
C0005937|T190|PT|733.21|ICD9CM|Solitary bone cyst|Solitary bone cyst
C0152244|T047|AB|733.22|ICD9CM|Aneurysmal bone cyst|Aneurysmal bone cyst
C0152244|T047|PT|733.22|ICD9CM|Aneurysmal bone cyst|Aneurysmal bone cyst
C0029525|T047|AB|733.29|ICD9CM|Bone cyst NEC|Bone cyst NEC
C0029525|T047|PT|733.29|ICD9CM|Other bone cyst|Other bone cyst
C0020496|T047|AB|733.3|ICD9CM|Hyperostosis of skull|Hyperostosis of skull
C0020496|T047|PT|733.3|ICD9CM|Hyperostosis of skull|Hyperostosis of skull
C0520474|T046|HT|733.4|ICD9CM|Aseptic necrosis of bone|Aseptic necrosis of bone
C0520474|T046|AB|733.40|ICD9CM|Asept necrosis bone NOS|Asept necrosis bone NOS
C0520474|T046|PT|733.40|ICD9CM|Aseptic necrosis of bone, site unspecified|Aseptic necrosis of bone, site unspecified
C0158449|T047|AB|733.41|ICD9CM|Aseptic necrosis humerus|Aseptic necrosis humerus
C0158449|T047|PT|733.41|ICD9CM|Aseptic necrosis of head of humerus|Aseptic necrosis of head of humerus
C0003977|T047|AB|733.42|ICD9CM|Aseptic necrosis femur|Aseptic necrosis femur
C0003977|T047|PT|733.42|ICD9CM|Aseptic necrosis of head and neck of femur|Aseptic necrosis of head and neck of femur
C0158450|T047|AB|733.43|ICD9CM|Asept necro femur condyl|Asept necro femur condyl
C0158450|T047|PT|733.43|ICD9CM|Aseptic necrosis of medial femoral condyle|Aseptic necrosis of medial femoral condyle
C0158451|T047|PT|733.44|ICD9CM|Aseptic necrosis of talus|Aseptic necrosis of talus
C0158451|T047|AB|733.44|ICD9CM|Aseptic necrosis talus|Aseptic necrosis talus
C1611734|T047|PT|733.45|ICD9CM|Aseptic necrosis of bone, jaw|Aseptic necrosis of bone, jaw
C1611734|T047|AB|733.45|ICD9CM|Aseptic necrosis of jaw|Aseptic necrosis of jaw
C0158452|T047|AB|733.49|ICD9CM|Asept necrosis bone NEC|Asept necrosis bone NEC
C0158452|T047|PT|733.49|ICD9CM|Aseptic necrosis of bone, other|Aseptic necrosis of bone, other
C0152263|T047|AB|733.5|ICD9CM|Osteitis condensans|Osteitis condensans
C0152263|T047|PT|733.5|ICD9CM|Osteitis condensans|Osteitis condensans
C0040213|T047|AB|733.6|ICD9CM|Tietze's disease|Tietze's disease
C0040213|T047|PT|733.6|ICD9CM|Tietze's disease|Tietze's disease
C0205930|T047|AB|733.7|ICD9CM|Algoneurodystrophy|Algoneurodystrophy
C0205930|T047|PT|733.7|ICD9CM|Algoneurodystrophy|Algoneurodystrophy
C0158453|T046|HT|733.8|ICD9CM|Malunion and nonunion of fracture|Malunion and nonunion of fracture
C0158454|T046|AB|733.81|ICD9CM|Malunion of fracture|Malunion of fracture
C0158454|T046|PT|733.81|ICD9CM|Malunion of fracture|Malunion of fracture
C0016665|T046|AB|733.82|ICD9CM|Nonunion of fracture|Nonunion of fracture
C0016665|T046|PT|733.82|ICD9CM|Nonunion of fracture|Nonunion of fracture
C0029586|T047|HT|733.9|ICD9CM|Other and unspecified disorders of bone and cartilage|Other and unspecified disorders of bone and cartilage
C0152091|T047|AB|733.90|ICD9CM|Bone & cartilage dis NOS|Bone & cartilage dis NOS
C0152091|T047|PT|733.90|ICD9CM|Disorder of bone and cartilage, unspecified|Disorder of bone and cartilage, unspecified
C0158456|T047|PT|733.91|ICD9CM|Arrest of bone development or growth|Arrest of bone development or growth
C0158456|T047|AB|733.91|ICD9CM|Arrest of bone growth|Arrest of bone growth
C0085700|T047|AB|733.92|ICD9CM|Chondromalacia|Chondromalacia
C0085700|T047|PT|733.92|ICD9CM|Chondromalacia|Chondromalacia
C0949138|T047|PT|733.93|ICD9CM|Stress fracture of tibia or fibula|Stress fracture of tibia or fibula
C0949138|T047|AB|733.93|ICD9CM|Stress fx tibia/fibula|Stress fx tibia/fibula
C0949139|T047|PT|733.94|ICD9CM|Stress fracture of the metatarsals|Stress fracture of the metatarsals
C0949139|T047|AB|733.94|ICD9CM|Stress fx metatarsals|Stress fx metatarsals
C0949140|T047|AB|733.95|ICD9CM|Stress fracture bone NEC|Stress fracture bone NEC
C0949140|T047|PT|733.95|ICD9CM|Stress fracture of other bone|Stress fracture of other bone
C2349651|T046|PT|733.96|ICD9CM|Stress fracture of femoral neck|Stress fracture of femoral neck
C2349651|T046|AB|733.96|ICD9CM|Stress fx femoral neck|Stress fx femoral neck
C2349653|T047|PT|733.97|ICD9CM|Stress fracture of shaft of femur|Stress fracture of shaft of femur
C2349653|T047|AB|733.97|ICD9CM|Stress fx shaft femur|Stress fx shaft femur
C2317110|T037|PT|733.98|ICD9CM|Stress fracture of pelvis|Stress fracture of pelvis
C2317110|T037|AB|733.98|ICD9CM|Stress fx pelvis|Stress fx pelvis
C0029586|T047|AB|733.99|ICD9CM|Bone & cartilage dis NEC|Bone & cartilage dis NEC
C0029586|T047|PT|733.99|ICD9CM|Other disorders of bone and cartilage|Other disorders of bone and cartilage
C0264133|T020|AB|734|ICD9CM|Flat foot|Flat foot
C0264133|T020|PT|734|ICD9CM|Flat foot|Flat foot
C0158457|T020|HT|735|ICD9CM|Acquired deformities of toe|Acquired deformities of toe
C0158458|T020|AB|735.0|ICD9CM|Hallux valgus|Hallux valgus
C0158458|T020|PT|735.0|ICD9CM|Hallux valgus (acquired)|Hallux valgus (acquired)
C0866710|T020|AB|735.1|ICD9CM|Hallux varus|Hallux varus
C0866710|T020|PT|735.1|ICD9CM|Hallux varus (acquired)|Hallux varus (acquired)
C0264134|T047|AB|735.2|ICD9CM|Hallux rigidus|Hallux rigidus
C0264134|T047|PT|735.2|ICD9CM|Hallux rigidus|Hallux rigidus
C0410779|T020|AB|735.3|ICD9CM|Hallux malleus|Hallux malleus
C0410779|T020|PT|735.3|ICD9CM|Hallux malleus|Hallux malleus
C0477572|T020|AB|735.4|ICD9CM|Other hammer toe|Other hammer toe
C0477572|T020|PT|735.4|ICD9CM|Other hammer toe (acquired)|Other hammer toe (acquired)
C0158461|T020|AB|735.5|ICD9CM|Claw toe|Claw toe
C0158461|T020|PT|735.5|ICD9CM|Claw toe (acquired)|Claw toe (acquired)
C0477573|T020|AB|735.8|ICD9CM|Acq deformity of toe NEC|Acq deformity of toe NEC
C0477573|T020|PT|735.8|ICD9CM|Other acquired deformities of toe|Other acquired deformities of toe
C0158457|T020|AB|735.9|ICD9CM|Acq deformity of toe NOS|Acq deformity of toe NOS
C0158457|T020|PT|735.9|ICD9CM|Unspecified acquired deformity of toe|Unspecified acquired deformity of toe
C0158463|T020|HT|736|ICD9CM|Other acquired deformities of limbs|Other acquired deformities of limbs
C0158464|T020|HT|736.0|ICD9CM|Acquired deformities of forearm, excluding fingers|Acquired deformities of forearm, excluding fingers
C0041784|T190|AB|736.00|ICD9CM|Forearm deformity NOS|Forearm deformity NOS
C0041784|T190|PT|736.00|ICD9CM|Unspecified deformity of forearm, excluding fingers|Unspecified deformity of forearm, excluding fingers
C0158465|T020|AB|736.01|ICD9CM|Cubitus valgus|Cubitus valgus
C0158465|T020|PT|736.01|ICD9CM|Cubitus valgus (acquired)|Cubitus valgus (acquired)
C0158466|T020|AB|736.02|ICD9CM|Cubitus varus|Cubitus varus
C0158466|T020|PT|736.02|ICD9CM|Cubitus varus (acquired)|Cubitus varus (acquired)
C0158467|T020|PT|736.03|ICD9CM|Valgus deformity of wrist (acquired)|Valgus deformity of wrist (acquired)
C0158467|T020|AB|736.03|ICD9CM|Valgus deformity wrist|Valgus deformity wrist
C0158468|T020|PT|736.04|ICD9CM|Varus deformity of wrist (acquired)|Varus deformity of wrist (acquired)
C0158468|T020|AB|736.04|ICD9CM|Varus deformity wrist|Varus deformity wrist
C0231666|T033|AB|736.05|ICD9CM|Wrist drop|Wrist drop
C0231666|T033|PT|736.05|ICD9CM|Wrist drop (acquired)|Wrist drop (acquired)
C0158470|T020|AB|736.06|ICD9CM|Claw hand|Claw hand
C0158470|T020|PT|736.06|ICD9CM|Claw hand (acquired)|Claw hand (acquired)
C0158471|T020|AB|736.07|ICD9CM|Club hand, acquired|Club hand, acquired
C0158471|T020|PT|736.07|ICD9CM|Club hand, acquired|Club hand, acquired
C0158472|T020|AB|736.09|ICD9CM|Forearm deformity NEC|Forearm deformity NEC
C0158472|T020|PT|736.09|ICD9CM|Other acquired deformities of forearm, excluding fingers|Other acquired deformities of forearm, excluding fingers
C0158473|T020|AB|736.1|ICD9CM|Mallet finger|Mallet finger
C0158473|T020|PT|736.1|ICD9CM|Mallet finger|Mallet finger
C0158474|T020|HT|736.2|ICD9CM|Other acquired deformities of finger|Other acquired deformities of finger
C0410740|T020|AB|736.20|ICD9CM|Acq finger deformity NOS|Acq finger deformity NOS
C0410740|T020|PT|736.20|ICD9CM|Unspecified deformity of finger|Unspecified deformity of finger
C0158476|T020|AB|736.21|ICD9CM|Boutonniere deformity|Boutonniere deformity
C0158476|T020|PT|736.21|ICD9CM|Boutonniere deformity|Boutonniere deformity
C0158477|T020|AB|736.22|ICD9CM|Swan-neck deformity|Swan-neck deformity
C0158477|T020|PT|736.22|ICD9CM|Swan-neck deformity|Swan-neck deformity
C0158474|T020|AB|736.29|ICD9CM|Acq finger deformity NEC|Acq finger deformity NEC
C0158474|T020|PT|736.29|ICD9CM|Other acquired deformities of finger|Other acquired deformities of finger
C0158478|T020|HT|736.3|ICD9CM|Acquired deformities of hip|Acquired deformities of hip
C0158478|T020|AB|736.30|ICD9CM|Acq hip deformity NOS|Acq hip deformity NOS
C0158478|T020|PT|736.30|ICD9CM|Unspecified acquired deformity of hip|Unspecified acquired deformity of hip
C0158480|T020|AB|736.31|ICD9CM|Coxa valga|Coxa valga
C0158480|T020|PT|736.31|ICD9CM|Coxa valga (acquired)|Coxa valga (acquired)
C0158481|T020|AB|736.32|ICD9CM|Coxa vara|Coxa vara
C0158481|T020|PT|736.32|ICD9CM|Coxa vara (acquired)|Coxa vara (acquired)
C0158482|T020|AB|736.39|ICD9CM|Acq hip deformity NEC|Acq hip deformity NEC
C0158482|T020|PT|736.39|ICD9CM|Other acquired deformities of hip|Other acquired deformities of hip
C0158483|T020|HT|736.4|ICD9CM|Genu valgum or varum (acquired)|Genu valgum or varum (acquired)
C0158484|T020|AB|736.41|ICD9CM|Genu valgum|Genu valgum
C0158484|T020|PT|736.41|ICD9CM|Genu valgum (acquired)|Genu valgum (acquired)
C0158485|T020|AB|736.42|ICD9CM|Genu varum|Genu varum
C0158485|T020|PT|736.42|ICD9CM|Genu varum (acquired)|Genu varum (acquired)
C0158486|T020|AB|736.5|ICD9CM|Genu recurvatum|Genu recurvatum
C0158486|T020|PT|736.5|ICD9CM|Genu recurvatum (acquired)|Genu recurvatum (acquired)
C0158487|T020|AB|736.6|ICD9CM|Acq knee deformity NEC|Acq knee deformity NEC
C0158487|T020|PT|736.6|ICD9CM|Other acquired deformities of knee|Other acquired deformities of knee
C0158488|T020|HT|736.7|ICD9CM|Other acquired deformities of ankle and foot|Other acquired deformities of ankle and foot
C0264150|T020|AB|736.70|ICD9CM|Acq ankle-foot def NOS|Acq ankle-foot def NOS
C0264150|T020|PT|736.70|ICD9CM|Unspecified deformity of ankle and foot, acquired|Unspecified deformity of ankle and foot, acquired
C0158489|T020|AB|736.71|ICD9CM|Acq equinovarus|Acq equinovarus
C0158489|T020|PT|736.71|ICD9CM|Acquired equinovarus deformity|Acquired equinovarus deformity
C0158490|T020|AB|736.72|ICD9CM|Acq equinus deformity|Acq equinus deformity
C0158490|T020|PT|736.72|ICD9CM|Equinus deformity of foot, acquired|Equinus deformity of foot, acquired
C2239098|T047|AB|736.73|ICD9CM|Cavus deformity of foot|Cavus deformity of foot
C2239098|T047|PT|736.73|ICD9CM|Cavus deformity of foot, acquired|Cavus deformity of foot, acquired
C0158461|T020|AB|736.74|ICD9CM|Claw foot, acquired|Claw foot, acquired
C0158461|T020|PT|736.74|ICD9CM|Claw foot, acquired|Claw foot, acquired
C0158493|T020|AB|736.75|ICD9CM|Acq cavovarus deformity|Acq cavovarus deformity
C0158493|T020|PT|736.75|ICD9CM|Cavovarus deformity of foot, acquired|Cavovarus deformity of foot, acquired
C0158494|T020|AB|736.76|ICD9CM|Calcaneus deformity NEC|Calcaneus deformity NEC
C0158494|T020|PT|736.76|ICD9CM|Other acquired calcaneus deformity|Other acquired calcaneus deformity
C0158488|T020|AB|736.79|ICD9CM|Acq ankle-foot def NEC|Acq ankle-foot def NEC
C0158488|T020|PT|736.79|ICD9CM|Other acquired deformities of ankle and foot|Other acquired deformities of ankle and foot
C0158495|T020|HT|736.8|ICD9CM|Acquired deformities of other parts of limbs|Acquired deformities of other parts of limbs
C0264156|T020|AB|736.81|ICD9CM|Unequal leg length|Unequal leg length
C0264156|T020|PT|736.81|ICD9CM|Unequal leg length (acquired)|Unequal leg length (acquired)
C0029486|T020|AB|736.89|ICD9CM|Oth acq limb deformity|Oth acq limb deformity
C0029486|T020|PT|736.89|ICD9CM|Other acquired deformity of other parts of limb|Other acquired deformity of other parts of limb
C0264155|T020|AB|736.9|ICD9CM|Acq limb deformity NOS|Acq limb deformity NOS
C0264155|T020|PT|736.9|ICD9CM|Acquired deformity of limb, site unspecified|Acquired deformity of limb, site unspecified
C0037932|T033|HT|737|ICD9CM|Curvature of spine|Curvature of spine
C0158497|T020|AB|737.0|ICD9CM|Adoles postural kyphosis|Adoles postural kyphosis
C0158497|T020|PT|737.0|ICD9CM|Adolescent postural kyphosis|Adolescent postural kyphosis
C0022822|T020|HT|737.1|ICD9CM|Kyphosis (acquired)|Kyphosis (acquired)
C0022823|T020|PT|737.10|ICD9CM|Kyphosis (acquired) (postural)|Kyphosis (acquired) (postural)
C0022823|T020|AB|737.10|ICD9CM|Kyphosis NOS|Kyphosis NOS
C0158498|T046|PT|737.11|ICD9CM|Kyphosis due to radiation|Kyphosis due to radiation
C0158498|T046|AB|737.11|ICD9CM|Radiation kyphosis|Radiation kyphosis
C0158499|T020|PT|737.12|ICD9CM|Kyphosis, postlaminectomy|Kyphosis, postlaminectomy
C0158499|T020|AB|737.12|ICD9CM|Postlaminectomy kyphosis|Postlaminectomy kyphosis
C0029653|T020|AB|737.19|ICD9CM|Kyphosis NEC|Kyphosis NEC
C0029653|T020|PT|737.19|ICD9CM|Other kyphosis (acquired)|Other kyphosis (acquired)
C0024004|T020|HT|737.2|ICD9CM|Lordosis (acquired)|Lordosis (acquired)
C0024005|T020|PT|737.20|ICD9CM|Lordosis (acquired) (postural)|Lordosis (acquired) (postural)
C0024005|T020|AB|737.20|ICD9CM|Lordosis NOS|Lordosis NOS
C0158500|T020|PT|737.21|ICD9CM|Lordosis, postlaminectomy|Lordosis, postlaminectomy
C0158500|T020|AB|737.21|ICD9CM|Postlaminectomy lordosis|Postlaminectomy lordosis
C0158501|T020|AB|737.22|ICD9CM|Oth postsurgery lordosis|Oth postsurgery lordosis
C0158501|T020|PT|737.22|ICD9CM|Other postsurgical lordosis|Other postsurgical lordosis
C0029658|T020|AB|737.29|ICD9CM|Lordosis NEC|Lordosis NEC
C0029658|T020|PT|737.29|ICD9CM|Other lordosis (acquired)|Other lordosis (acquired)
C0022820|T190|HT|737.3|ICD9CM|Kyphoscoliosis and scoliosis|Kyphoscoliosis and scoliosis
C0036440|T190|AB|737.30|ICD9CM|Idiopathic scoliosis|Idiopathic scoliosis
C0036440|T190|PT|737.30|ICD9CM|Scoliosis [and kyphoscoliosis], idiopathic|Scoliosis [and kyphoscoliosis], idiopathic
C0158502|T020|AB|737.31|ICD9CM|Resolv idiopath scolios|Resolv idiopath scolios
C0158502|T020|PT|737.31|ICD9CM|Resolving infantile idiopathic scoliosis|Resolving infantile idiopathic scoliosis
C0158503|T047|AB|737.32|ICD9CM|Progr idiopath scoliosis|Progr idiopath scoliosis
C0158503|T047|PT|737.32|ICD9CM|Progressive infantile idiopathic scoliosis|Progressive infantile idiopathic scoliosis
C0158504|T046|AB|737.33|ICD9CM|Radiation scoliosis|Radiation scoliosis
C0158504|T046|PT|737.33|ICD9CM|Scoliosis due to radiation|Scoliosis due to radiation
C0158505|T047|AB|737.34|ICD9CM|Thoracogenic scoliosis|Thoracogenic scoliosis
C0158505|T047|PT|737.34|ICD9CM|Thoracogenic scoliosis|Thoracogenic scoliosis
C0029652|T047|PT|737.39|ICD9CM|Other kyphoscoliosis and scoliosis|Other kyphoscoliosis and scoliosis
C0029652|T047|AB|737.39|ICD9CM|Scoliosis NEC|Scoliosis NEC
C0158506|T190|HT|737.4|ICD9CM|Curvature of spine associated with other conditions|Curvature of spine associated with other conditions
C0158506|T190|PT|737.40|ICD9CM|Curvature of spine, unspecified, associated with other conditions|Curvature of spine, unspecified, associated with other conditions
C0158506|T190|AB|737.40|ICD9CM|Spin curv NOS in oth dis|Spin curv NOS in oth dis
C0158507|T047|PT|737.41|ICD9CM|Kyphosis associated with other conditions|Kyphosis associated with other conditions
C0158507|T047|AB|737.41|ICD9CM|Kyphosis in oth dis|Kyphosis in oth dis
C0158508|T047|PT|737.42|ICD9CM|Lordosis associated with other conditions|Lordosis associated with other conditions
C0158508|T047|AB|737.42|ICD9CM|Lordosis in oth dis|Lordosis in oth dis
C0158509|T047|PT|737.43|ICD9CM|Scoliosis associated with other conditions|Scoliosis associated with other conditions
C0158509|T047|AB|737.43|ICD9CM|Scoliosis in oth dis|Scoliosis in oth dis
C0410693|T020|AB|737.8|ICD9CM|Curvature of spine NEC|Curvature of spine NEC
C0410693|T020|PT|737.8|ICD9CM|Other curvatures of spine|Other curvatures of spine
C0158506|T190|AB|737.9|ICD9CM|Curvature of spine NOS|Curvature of spine NOS
C0158506|T190|PT|737.9|ICD9CM|Unspecified curvature of spine|Unspecified curvature of spine
C0158510|T020|HT|738|ICD9CM|Other acquired musculoskeletal deformity|Other acquired musculoskeletal deformity
C0028431|T020|AB|738.0|ICD9CM|Acq nose deformity|Acq nose deformity
C0028431|T020|PT|738.0|ICD9CM|Acquired deformity of nose|Acquired deformity of nose
C0158511|T020|HT|738.1|ICD9CM|Other acquired deformity of head|Other acquired deformity of head
C1290220|T020|PT|738.10|ICD9CM|Unspecified acquired deformity of head|Unspecified acquired deformity of head
C1290220|T020|AB|738.10|ICD9CM|Unspf acq deformity head|Unspf acq deformity head
C4082244|T047|AB|738.11|ICD9CM|Zygomatic hyperplasia|Zygomatic hyperplasia
C4082244|T047|PT|738.11|ICD9CM|Zygomatic hyperplasia|Zygomatic hyperplasia
C0375512|T020|AB|738.12|ICD9CM|Zygomatic hypoplasia|Zygomatic hypoplasia
C0375512|T020|PT|738.12|ICD9CM|Zygomatic hypoplasia|Zygomatic hypoplasia
C0375513|T020|AB|738.19|ICD9CM|Oth spcf deformity head|Oth spcf deformity head
C0375513|T020|PT|738.19|ICD9CM|Other specified acquired deformity of head|Other specified acquired deformity of head
C0158512|T020|AB|738.2|ICD9CM|Acq neck deformity|Acq neck deformity
C0158512|T020|PT|738.2|ICD9CM|Acquired deformity of neck|Acquired deformity of neck
C0001171|T020|AB|738.3|ICD9CM|Acq chest deformity|Acq chest deformity
C0001171|T020|PT|738.3|ICD9CM|Acquired deformity of chest and rib|Acquired deformity of chest and rib
C2242765|T020|AB|738.4|ICD9CM|Acq spondylolisthesis|Acq spondylolisthesis
C2242765|T020|PT|738.4|ICD9CM|Acquired spondylolisthesis|Acquired spondylolisthesis
C0158514|T020|AB|738.5|ICD9CM|Other acq back deformity|Other acq back deformity
C0158514|T020|PT|738.5|ICD9CM|Other acquired deformity of back or spine|Other acquired deformity of back or spine
C0158515|T020|AB|738.6|ICD9CM|Acq pelvic deformity|Acq pelvic deformity
C0158515|T020|PT|738.6|ICD9CM|Acquired deformity of pelvis|Acquired deformity of pelvis
C0158516|T020|AB|738.7|ICD9CM|Cauliflower ear|Cauliflower ear
C0158516|T020|PT|738.7|ICD9CM|Cauliflower ear|Cauliflower ear
C0158517|T020|AB|738.8|ICD9CM|Acq deformity NEC|Acq deformity NEC
C0158517|T020|PT|738.8|ICD9CM|Acquired deformity of other specified site|Acquired deformity of other specified site
C0264132|T020|AB|738.9|ICD9CM|Acq deformity NOS|Acq deformity NOS
C0264132|T020|PT|738.9|ICD9CM|Acquired deformity of unspecified site|Acquired deformity of unspecified site
C0869269|T047|HT|739|ICD9CM|Nonallopathic lesions, not elsewhere classified|Nonallopathic lesions, not elsewhere classified
C0877720|T047|PT|739.0|ICD9CM|Nonallopathic lesions, head region|Nonallopathic lesions, head region
C0877720|T047|AB|739.0|ICD9CM|Somat dys head region|Somat dys head region
C0877722|T047|PT|739.1|ICD9CM|Nonallopathic lesions, cervical region|Nonallopathic lesions, cervical region
C0877722|T047|AB|739.1|ICD9CM|Somat dysfunc cervic reg|Somat dysfunc cervic reg
C0877724|T047|PT|739.2|ICD9CM|Nonallopathic lesions, thoracic region|Nonallopathic lesions, thoracic region
C0877724|T047|AB|739.2|ICD9CM|Somat dysfunc thorac reg|Somat dysfunc thorac reg
C0877726|T047|PT|739.3|ICD9CM|Nonallopathic lesions, lumbar region|Nonallopathic lesions, lumbar region
C0877726|T047|AB|739.3|ICD9CM|Somat dysfunc lumbar reg|Somat dysfunc lumbar reg
C0877728|T047|PT|739.4|ICD9CM|Nonallopathic lesions, sacral region|Nonallopathic lesions, sacral region
C0877728|T047|AB|739.4|ICD9CM|Somat dysfunc sacral reg|Somat dysfunc sacral reg
C0877730|T047|PT|739.5|ICD9CM|Nonallopathic lesions, pelvic region|Nonallopathic lesions, pelvic region
C0877730|T047|AB|739.5|ICD9CM|Somat dysfunc pelvic reg|Somat dysfunc pelvic reg
C0877732|T047|PT|739.6|ICD9CM|Nonallopathic lesions, lower extremities|Nonallopathic lesions, lower extremities
C0877732|T047|AB|739.6|ICD9CM|Somat dysfunc lower extr|Somat dysfunc lower extr
C0877734|T047|PT|739.7|ICD9CM|Nonallopathic lesions, upper extremities|Nonallopathic lesions, upper extremities
C0877734|T047|AB|739.7|ICD9CM|Somat dysfunc upper extr|Somat dysfunc upper extr
C0877736|T047|PT|739.8|ICD9CM|Nonallopathic lesions, rib cage|Nonallopathic lesions, rib cage
C0877736|T047|AB|739.8|ICD9CM|Somat dysfunc rib cage|Somat dysfunc rib cage
C0302396|T047|PT|739.9|ICD9CM|Nonallopathic lesions, abdomen and other sites|Nonallopathic lesions, abdomen and other sites
C0302396|T047|AB|739.9|ICD9CM|Somatic dysfunction NEC|Somatic dysfunction NEC
C0158530|T019|HT|740|ICD9CM|Anencephalus and similar anomalies|Anencephalus and similar anomalies
C0000768|T019|HT|740-759.99|ICD9CM|CONGENITAL ANOMALIES|CONGENITAL ANOMALIES
C0002902|T019|AB|740.0|ICD9CM|Anencephalus|Anencephalus
C0002902|T019|PT|740.0|ICD9CM|Anencephalus|Anencephalus
C0152426|T019|AB|740.1|ICD9CM|Craniorachischisis|Craniorachischisis
C0152426|T019|PT|740.1|ICD9CM|Craniorachischisis|Craniorachischisis
C0152234|T019|AB|740.2|ICD9CM|Iniencephaly|Iniencephaly
C0152234|T019|PT|740.2|ICD9CM|Iniencephaly|Iniencephaly
C0080178|T019|HT|741|ICD9CM|Spina bifida|Spina bifida
C0477973|T019|HT|741.0|ICD9CM|Spina bifida with hydrocephalus|Spina bifida with hydrocephalus
C0477973|T019|AB|741.00|ICD9CM|Spin bif w hydroceph NOS|Spin bif w hydroceph NOS
C0477973|T019|PT|741.00|ICD9CM|Spina bifida with hydrocephalus, unspecified region|Spina bifida with hydrocephalus, unspecified region
C0431321|T019|AB|741.01|ICD9CM|Spin bif w hydrceph-cerv|Spin bif w hydrceph-cerv
C0431321|T019|PT|741.01|ICD9CM|Spina bifida with hydrocephalus, cervical region|Spina bifida with hydrocephalus, cervical region
C0431320|T019|AB|741.02|ICD9CM|Spin bif w hydrceph-dors|Spin bif w hydrceph-dors
C0431320|T019|PT|741.02|ICD9CM|Spina bifida with hydrocephalus, dorsal (thoracic) region|Spina bifida with hydrocephalus, dorsal (thoracic) region
C0431319|T019|AB|741.03|ICD9CM|Spin bif w hydrceph-lumb|Spin bif w hydrceph-lumb
C0431319|T019|PT|741.03|ICD9CM|Spina bifida with hydrocephalus, lumbar region|Spina bifida with hydrocephalus, lumbar region
C0158534|T019|HT|741.9|ICD9CM|Spina bifida without mention of hydrocephalus|Spina bifida without mention of hydrocephalus
C0158534|T019|AB|741.90|ICD9CM|Spina bifida|Spina bifida
C0158534|T019|PT|741.90|ICD9CM|Spina bifida without mention of hydrocephalus, unspecified region|Spina bifida without mention of hydrocephalus, unspecified region
C0158535|T019|PT|741.91|ICD9CM|Spina bifida without mention of hydrocephalus, cervical region|Spina bifida without mention of hydrocephalus, cervical region
C0158535|T019|AB|741.91|ICD9CM|Spina bifida-cerv|Spina bifida-cerv
C0158536|T019|PT|741.92|ICD9CM|Spina bifida without mention of hydrocephalus, dorsal (thoracic) region|Spina bifida without mention of hydrocephalus, dorsal (thoracic) region
C0158536|T019|AB|741.92|ICD9CM|Spina bifida-dorsal|Spina bifida-dorsal
C0158537|T019|PT|741.93|ICD9CM|Spina bifida without mention of hydrocephalus, lumbar region|Spina bifida without mention of hydrocephalus, lumbar region
C0158537|T019|AB|741.93|ICD9CM|Spina bifida-lumbar|Spina bifida-lumbar
C0158538|T019|HT|742|ICD9CM|Other congenital anomalies of nervous system|Other congenital anomalies of nervous system
C4551722|T019|AB|742.0|ICD9CM|Encephalocele|Encephalocele
C4551722|T019|PT|742.0|ICD9CM|Encephalocele|Encephalocele
C0025958|T019|AB|742.1|ICD9CM|Microcephalus|Microcephalus
C0025958|T019|PT|742.1|ICD9CM|Microcephalus|Microcephalus
C0079157|T019|PT|742.2|ICD9CM|Congenital reduction deformities of brain|Congenital reduction deformities of brain
C0079157|T019|AB|742.2|ICD9CM|Reduction deform, brain|Reduction deform, brain
C0020256|T019|AB|742.3|ICD9CM|Congenital hydrocephalus|Congenital hydrocephalus
C0020256|T019|PT|742.3|ICD9CM|Congenital hydrocephalus|Congenital hydrocephalus
C0477972|T019|AB|742.4|ICD9CM|Brain anomaly NEC|Brain anomaly NEC
C0477972|T019|PT|742.4|ICD9CM|Other specified congenital anomalies of brain|Other specified congenital anomalies of brain
C0477975|T019|HT|742.5|ICD9CM|Other specified congenital anomalies of spinal cord|Other specified congenital anomalies of spinal cord
C0011999|T019|AB|742.51|ICD9CM|Diastematomyelia|Diastematomyelia
C0011999|T019|PT|742.51|ICD9CM|Diastematomyelia|Diastematomyelia
C0152444|T047|AB|742.53|ICD9CM|Hydromyelia|Hydromyelia
C0152444|T047|PT|742.53|ICD9CM|Hydromyelia|Hydromyelia
C0477975|T019|PT|742.59|ICD9CM|Other specified congenital anomalies of spinal cord|Other specified congenital anomalies of spinal cord
C0477975|T019|AB|742.59|ICD9CM|Spinal cord anomaly NEC|Spinal cord anomaly NEC
C0477976|T019|AB|742.8|ICD9CM|Nervous system anom NEC|Nervous system anom NEC
C0477976|T019|PT|742.8|ICD9CM|Other specified congenital anomalies of nervous system|Other specified congenital anomalies of nervous system
C0497552|T019|AB|742.9|ICD9CM|Nervous system anom NOS|Nervous system anom NOS
C0497552|T019|PT|742.9|ICD9CM|Unspecified congenital anomaly of brain, spinal cord, and nervous system|Unspecified congenital anomaly of brain, spinal cord, and nervous system
C0015393|T019|HT|743|ICD9CM|Congenital anomalies of eye|Congenital anomalies of eye
C0003119|T019|HT|743.0|ICD9CM|Anophthalmos|Anophthalmos
C0003119|T019|AB|743.00|ICD9CM|Clinic anophthalmos NOS|Clinic anophthalmos NOS
C0003119|T019|PT|743.00|ICD9CM|Clinical anophthalmos, unspecified|Clinical anophthalmos, unspecified
C0158543|T019|AB|743.03|ICD9CM|Congen cystic eyeball|Congen cystic eyeball
C0158543|T019|PT|743.03|ICD9CM|Cystic eyeball, congenital|Cystic eyeball, congenital
C0311249|T019|AB|743.06|ICD9CM|Cryptophthalmos|Cryptophthalmos
C0311249|T019|PT|743.06|ICD9CM|Cryptophthalmos|Cryptophthalmos
C0026010|T019|HT|743.1|ICD9CM|Microphthalmos|Microphthalmos
C0026010|T019|AB|743.10|ICD9CM|Microphthalmos NOS|Microphthalmos NOS
C0026010|T019|PT|743.10|ICD9CM|Microphthalmos, unspecified|Microphthalmos, unspecified
C0026010|T019|AB|743.11|ICD9CM|Simple microphthalmos|Simple microphthalmos
C0026010|T019|PT|743.11|ICD9CM|Simple microphthalmos|Simple microphthalmos
C0158545|T019|AB|743.12|ICD9CM|Microphth w oth eye anom|Microphth w oth eye anom
C0158545|T019|PT|743.12|ICD9CM|Microphthalmos associated with other anomalies of eye and adnexa|Microphthalmos associated with other anomalies of eye and adnexa
C4551507|T019|HT|743.2|ICD9CM|Buphthalmos|Buphthalmos
C4551507|T019|AB|743.20|ICD9CM|Buphthalmos NOS|Buphthalmos NOS
C4551507|T019|PT|743.20|ICD9CM|Buphthalmos, unspecified|Buphthalmos, unspecified
C0311251|T019|AB|743.21|ICD9CM|Simple buphthalmos|Simple buphthalmos
C0311251|T019|PT|743.21|ICD9CM|Simple buphthalmos|Simple buphthalmos
C0158547|T019|AB|743.22|ICD9CM|Buphthal w oth eye anom|Buphthal w oth eye anom
C0158547|T019|PT|743.22|ICD9CM|Buphthalmos associated with other ocular anomalies|Buphthalmos associated with other ocular anomalies
C0158548|T019|HT|743.3|ICD9CM|Congenital cataract and lens anomalies|Congenital cataract and lens anomalies
C0009691|T019|AB|743.30|ICD9CM|Congenital cataract NOS|Congenital cataract NOS
C0009691|T019|PT|743.30|ICD9CM|Congenital cataract, unspecified|Congenital cataract, unspecified
C0158549|T019|AB|743.31|ICD9CM|Capsular cataract|Capsular cataract
C0158549|T019|PT|743.31|ICD9CM|Congenital capsular and subcapsular cataract|Congenital capsular and subcapsular cataract
C0489970|T019|PT|743.32|ICD9CM|Congenital cortical and zonular cataract|Congenital cortical and zonular cataract
C0489970|T019|AB|743.32|ICD9CM|Cortical/zonular catarac|Cortical/zonular catarac
C0158551|T019|PT|743.33|ICD9CM|Congenital nuclear cataract|Congenital nuclear cataract
C0158551|T019|AB|743.33|ICD9CM|Nuclear cataract|Nuclear cataract
C0158552|T019|AB|743.34|ICD9CM|Cong tot/subtot cataract|Cong tot/subtot cataract
C0158552|T019|PT|743.34|ICD9CM|Total and subtotal cataract, congenital|Total and subtotal cataract, congenital
C0152422|T019|AB|743.35|ICD9CM|Congenital aphakia|Congenital aphakia
C0152422|T019|PT|743.35|ICD9CM|Congenital aphakia|Congenital aphakia
C0158553|T019|AB|743.36|ICD9CM|Anomalies of lens shape|Anomalies of lens shape
C0158553|T019|PT|743.36|ICD9CM|Congenital anomalies of lens shape|Congenital anomalies of lens shape
C0013581|T019|PT|743.37|ICD9CM|Congenital ectopic lens|Congenital ectopic lens
C0013581|T019|AB|743.37|ICD9CM|Congenital ectopic lens|Congenital ectopic lens
C0158554|T019|AB|743.39|ICD9CM|Cong catar/lens anom NEC|Cong catar/lens anom NEC
C0158554|T019|PT|743.39|ICD9CM|Other congenital cataract and lens anomalies|Other congenital cataract and lens anomalies
C0158555|T019|HT|743.4|ICD9CM|Coloboma and other anomalies of anterior segment|Coloboma and other anomalies of anterior segment
C0344528|T019|AB|743.41|ICD9CM|Anom corneal size/shape|Anom corneal size/shape
C0344528|T019|PT|743.41|ICD9CM|Congenital anomalies of corneal size and shape|Congenital anomalies of corneal size and shape
C0158557|T019|AB|743.42|ICD9CM|Cong cornea opac aff vis|Cong cornea opac aff vis
C0158557|T019|PT|743.42|ICD9CM|Corneal opacities, interfering with vision, congenital|Corneal opacities, interfering with vision, congenital
C0158558|T019|AB|743.43|ICD9CM|Cong corneal opacit NEC|Cong corneal opacit NEC
C0158558|T019|PT|743.43|ICD9CM|Other corneal opacities, congenital|Other corneal opacities, congenital
C0701146|T019|AB|743.44|ICD9CM|Anom anter chamber-eye|Anom anter chamber-eye
C0701146|T019|PT|743.44|ICD9CM|Specified congenital anomalies of anterior chamber, chamber angle, and related structures|Specified congenital anomalies of anterior chamber, chamber angle, and related structures
C0003076|T019|AB|743.45|ICD9CM|Aniridia|Aniridia
C0003076|T019|PT|743.45|ICD9CM|Aniridia|Aniridia
C0158560|T047|AB|743.46|ICD9CM|Anom iris & cil body NEC|Anom iris & cil body NEC
C0158560|T047|PT|743.46|ICD9CM|Other specified congenital anomalies of iris and ciliary body|Other specified congenital anomalies of iris and ciliary body
C0344538|T019|AB|743.47|ICD9CM|Anomalies of sclera|Anomalies of sclera
C0344538|T019|PT|743.47|ICD9CM|Specified congenital anomalies of sclera|Specified congenital anomalies of sclera
C0158562|T019|AB|743.48|ICD9CM|Mult anom anter seg-eye|Mult anom anter seg-eye
C0158562|T019|PT|743.48|ICD9CM|Multiple and combined congenital anomalies of anterior segment|Multiple and combined congenital anomalies of anterior segment
C0029552|T019|AB|743.49|ICD9CM|Anom anter seg NEC-eye|Anom anter seg NEC-eye
C0029552|T019|PT|743.49|ICD9CM|Other congenital anomalies of anterior segment|Other congenital anomalies of anterior segment
C0439001|T019|HT|743.5|ICD9CM|Congenital anomalies of posterior segment|Congenital anomalies of posterior segment
C0158564|T019|AB|743.51|ICD9CM|Vitreous anomalies|Vitreous anomalies
C0158564|T019|PT|743.51|ICD9CM|Vitreous anomalies|Vitreous anomalies
C0240896|T019|AB|743.52|ICD9CM|Fundus coloboma|Fundus coloboma
C0240896|T019|PT|743.52|ICD9CM|Fundus coloboma|Fundus coloboma
C0158566|T047|PT|743.53|ICD9CM|Chorioretinal degeneration, congenital|Chorioretinal degeneration, congenital
C0158566|T047|AB|743.53|ICD9CM|Cong chorioretinal degen|Cong chorioretinal degen
C0158567|T019|AB|743.54|ICD9CM|Cong fold/cyst post eye|Cong fold/cyst post eye
C0158567|T019|PT|743.54|ICD9CM|Congenital folds and cysts of posterior segment|Congenital folds and cysts of posterior segment
C0158568|T047|AB|743.55|ICD9CM|Cong macular change-eye|Cong macular change-eye
C0158568|T047|PT|743.55|ICD9CM|Congenital macular changes|Congenital macular changes
C0029729|T047|AB|743.56|ICD9CM|Cong retinal changes NEC|Cong retinal changes NEC
C0029729|T047|PT|743.56|ICD9CM|Other retinal changes, congenital|Other retinal changes, congenital
C0344553|T019|AB|743.57|ICD9CM|Optic disc anomalies|Optic disc anomalies
C0344553|T019|PT|743.57|ICD9CM|Specified congenital anomalies of optic disc|Specified congenital anomalies of optic disc
C1961121|T019|AB|743.58|ICD9CM|Vascular anom post eye|Vascular anom post eye
C1961121|T019|PT|743.58|ICD9CM|Vascular anomalies|Vascular anomalies
C0158571|T019|PT|743.59|ICD9CM|Other congenital anomalies of posterior segment|Other congenital anomalies of posterior segment
C0158571|T019|AB|743.59|ICD9CM|Post segmnt anom NEC-eye|Post segmnt anom NEC-eye
C0158572|T019|HT|743.6|ICD9CM|Congenital anomalies of eyelids, lacrimal system, and orbit|Congenital anomalies of eyelids, lacrimal system, and orbit
C0266573|T019|AB|743.61|ICD9CM|Congenital ptosis|Congenital ptosis
C0266573|T019|PT|743.61|ICD9CM|Congenital ptosis|Congenital ptosis
C0266572|T019|PT|743.62|ICD9CM|Congenital deformities of eyelids|Congenital deformities of eyelids
C0266572|T019|AB|743.62|ICD9CM|Congenital eyelid deform|Congenital eyelid deform
C0158575|T019|PT|743.63|ICD9CM|Other specified congenital anomalies of eyelid|Other specified congenital anomalies of eyelid
C0158575|T019|AB|743.63|ICD9CM|Spec anom of eyelid NEC|Spec anom of eyelid NEC
C0158576|T019|AB|743.64|ICD9CM|Spec lacrimal gland anom|Spec lacrimal gland anom
C0158576|T019|PT|743.64|ICD9CM|Specified congenital anomalies of lacrimal gland|Specified congenital anomalies of lacrimal gland
C0158577|T019|AB|743.65|ICD9CM|Spec lacrimal pass anom|Spec lacrimal pass anom
C0158577|T019|PT|743.65|ICD9CM|Specified congenital anomalies of lacrimal passages|Specified congenital anomalies of lacrimal passages
C0266587|T019|AB|743.66|ICD9CM|Spec anomaly of orbit|Spec anomaly of orbit
C0266587|T019|PT|743.66|ICD9CM|Specified congenital anomalies of orbit|Specified congenital anomalies of orbit
C0158579|T047|AB|743.69|ICD9CM|Anom eyelid/lacr/orb NEC|Anom eyelid/lacr/orb NEC
C0158579|T047|PT|743.69|ICD9CM|Other congenital anomalies of eyelids, lacrimal system, and orbit|Other congenital anomalies of eyelids, lacrimal system, and orbit
C0477986|T019|AB|743.8|ICD9CM|Eye anomalies NEC|Eye anomalies NEC
C0477986|T019|PT|743.8|ICD9CM|Other specified anomalies of eye|Other specified anomalies of eye
C0015393|T019|AB|743.9|ICD9CM|Eye anomaly NOS|Eye anomaly NOS
C0015393|T019|PT|743.9|ICD9CM|Unspecified anomaly of eye|Unspecified anomaly of eye
C0158581|T019|HT|744|ICD9CM|Congenital anomalies of ear, face, and neck|Congenital anomalies of ear, face, and neck
C0266592|T019|HT|744.0|ICD9CM|Congenital anomalies of ear causing impairment of hearing|Congenital anomalies of ear causing impairment of hearing
C0266592|T019|AB|744.00|ICD9CM|Ear anom NOS/impair hear|Ear anom NOS/impair hear
C0266592|T019|PT|744.00|ICD9CM|Unspecified anomaly of ear with impairment of hearing|Unspecified anomaly of ear with impairment of hearing
C0702139|T019|PT|744.01|ICD9CM|Absence of external ear|Absence of external ear
C0702139|T019|AB|744.01|ICD9CM|Cong absence ext ear|Cong absence ext ear
C0431467|T019|AB|744.02|ICD9CM|Ex ear anm NEC-impr hear|Ex ear anm NEC-impr hear
C0431467|T019|PT|744.02|ICD9CM|Other anomalies of external ear with impairment of hearing|Other anomalies of external ear with impairment of hearing
C0431468|T019|PT|744.03|ICD9CM|Anomaly of middle ear, except ossicles|Anomaly of middle ear, except ossicles
C0431468|T019|AB|744.03|ICD9CM|Middle ear anomaly NEC|Middle ear anomaly NEC
C0158587|T019|AB|744.04|ICD9CM|Anomalies ear ossicles|Anomalies ear ossicles
C0158587|T019|PT|744.04|ICD9CM|Anomalies of ear ossicles|Anomalies of ear ossicles
C0685874|T019|AB|744.05|ICD9CM|Anomalies of inner ear|Anomalies of inner ear
C0685874|T019|PT|744.05|ICD9CM|Anomalies of inner ear|Anomalies of inner ear
C0158589|T019|AB|744.09|ICD9CM|Ear anom NEC/impair hear|Ear anom NEC/impair hear
C0158589|T019|PT|744.09|ICD9CM|Other anomalies of ear causing impairment of hearing|Other anomalies of ear causing impairment of hearing
C0266611|T019|AB|744.1|ICD9CM|Accessory auricle|Accessory auricle
C0266611|T019|PT|744.1|ICD9CM|Accessory auricle|Accessory auricle
C0477990|T019|HT|744.2|ICD9CM|Other specified congenital anomalies of ear|Other specified congenital anomalies of ear
C0158591|T019|PT|744.21|ICD9CM|Absence of ear lobe, congenital|Absence of ear lobe, congenital
C0158591|T019|AB|744.21|ICD9CM|Cong absence of ear lobe|Cong absence of ear lobe
C0152421|T019|AB|744.22|ICD9CM|Macrotia|Macrotia
C0152421|T019|PT|744.22|ICD9CM|Macrotia|Macrotia
C0152423|T019|AB|744.23|ICD9CM|Microtia|Microtia
C0152423|T019|PT|744.23|ICD9CM|Microtia|Microtia
C0158592|T019|AB|744.24|ICD9CM|Eustachian tube anom NEC|Eustachian tube anom NEC
C0158592|T019|PT|744.24|ICD9CM|Specified anomalies of Eustachian tube|Specified anomalies of Eustachian tube
C0431479|T019|AB|744.29|ICD9CM|Ear anomalies NEC|Ear anomalies NEC
C0431479|T019|PT|744.29|ICD9CM|Other specified anomalies of ear|Other specified anomalies of ear
C0266589|T019|AB|744.3|ICD9CM|Ear anomaly NOS|Ear anomaly NOS
C0266589|T019|PT|744.3|ICD9CM|Unspecified anomaly of ear|Unspecified anomaly of ear
C0158595|T047|HT|744.4|ICD9CM|Branchial cleft cyst or fistula; preauricular sinus|Branchial cleft cyst or fistula; preauricular sinus
C0344572|T047|AB|744.41|ICD9CM|Branch cleft sinus/fistu|Branch cleft sinus/fistu
C0344572|T047|PT|744.41|ICD9CM|Branchial cleft sinus or fistula|Branchial cleft sinus or fistula
C0006131|T019|AB|744.42|ICD9CM|Branchial cleft cyst|Branchial cleft cyst
C0006131|T019|PT|744.42|ICD9CM|Branchial cleft cyst|Branchial cleft cyst
C2363280|T019|AB|744.43|ICD9CM|Cervical auricle|Cervical auricle
C2363280|T019|PT|744.43|ICD9CM|Cervical auricle|Cervical auricle
C0158598|T047|PT|744.46|ICD9CM|Preauricular sinus or fistula|Preauricular sinus or fistula
C0158598|T047|AB|744.46|ICD9CM|Preauricular sinus/fistu|Preauricular sinus/fistu
C0158599|T047|AB|744.47|ICD9CM|Preauricular cyst|Preauricular cyst
C0158599|T047|PT|744.47|ICD9CM|Preauricular cyst|Preauricular cyst
C0431491|T047|AB|744.49|ICD9CM|Branchial cleft anom NEC|Branchial cleft anom NEC
C0431491|T047|PT|744.49|ICD9CM|Other branchial cleft cyst or fistula; preauricular sinus|Other branchial cleft cyst or fistula; preauricular sinus
C0221217|T019|AB|744.5|ICD9CM|Webbing of neck|Webbing of neck
C0221217|T019|PT|744.5|ICD9CM|Webbing of neck|Webbing of neck
C0477992|T019|HT|744.8|ICD9CM|Other specified congenital anomalies of face and neck|Other specified congenital anomalies of face and neck
C0266094|T019|AB|744.81|ICD9CM|Macrocheilia|Macrocheilia
C0266094|T019|PT|744.81|ICD9CM|Macrocheilia|Macrocheilia
C0266095|T019|AB|744.82|ICD9CM|Microcheilia|Microcheilia
C0266095|T019|PT|744.82|ICD9CM|Microcheilia|Microcheilia
C0024433|T019|AB|744.83|ICD9CM|Macrostomia|Macrostomia
C0024433|T019|PT|744.83|ICD9CM|Macrostomia|Macrostomia
C0026034|T019|AB|744.84|ICD9CM|Microstomia|Microstomia
C0026034|T019|PT|744.84|ICD9CM|Microstomia|Microstomia
C0477992|T019|AB|744.89|ICD9CM|Cong face/neck anom NEC|Cong face/neck anom NEC
C0477992|T019|PT|744.89|ICD9CM|Other specified congenital anomalies of face and neck|Other specified congenital anomalies of face and neck
C0869095|T019|AB|744.9|ICD9CM|Cong face/neck anom NOS|Cong face/neck anom NOS
C0869095|T019|PT|744.9|ICD9CM|Unspecified congenital anomalies of face and neck|Unspecified congenital anomalies of face and neck
C0158606|T019|HT|745|ICD9CM|Bulbus cordis anomalies and anomalies of cardiac septal closure|Bulbus cordis anomalies and anomalies of cardiac septal closure
C0041207|T019|AB|745.0|ICD9CM|Common truncus|Common truncus
C0041207|T019|PT|745.0|ICD9CM|Common truncus|Common truncus
C0040761|T019|HT|745.1|ICD9CM|Transposition of great vessels|Transposition of great vessels
C0040761|T019|AB|745.10|ICD9CM|Compl transpos great ves|Compl transpos great ves
C0040761|T019|PT|745.10|ICD9CM|Complete transposition of great vessels|Complete transposition of great vessels
C0013069|T019|PT|745.11|ICD9CM|Double outlet right ventricle|Double outlet right ventricle
C0013069|T019|AB|745.11|ICD9CM|Double outlet rt ventric|Double outlet rt ventric
C0344616|T019|AB|745.12|ICD9CM|Correct transpos grt ves|Correct transpos grt ves
C0344616|T019|PT|745.12|ICD9CM|Corrected transposition of great vessels|Corrected transposition of great vessels
C0158608|T019|PT|745.19|ICD9CM|Other transposition of great vessels|Other transposition of great vessels
C0158608|T019|AB|745.19|ICD9CM|Transpos great vess NEC|Transpos great vess NEC
C0039685|T019|AB|745.2|ICD9CM|Tetralogy of fallot|Tetralogy of fallot
C0039685|T019|PT|745.2|ICD9CM|Tetralogy of fallot|Tetralogy of fallot
C0152424|T019|AB|745.3|ICD9CM|Common ventricle|Common ventricle
C0152424|T019|PT|745.3|ICD9CM|Common ventricle|Common ventricle
C0018818|T019|AB|745.4|ICD9CM|Ventricular sept defect|Ventricular sept defect
C0018818|T019|PT|745.4|ICD9CM|Ventricular septal defect|Ventricular septal defect
C0344724|T019|PT|745.5|ICD9CM|Ostium secundum type atrial septal defect|Ostium secundum type atrial septal defect
C0344724|T019|AB|745.5|ICD9CM|Secundum atrial sept def|Secundum atrial sept def
C0014116|T019|HT|745.6|ICD9CM|Endocardial cushion defects|Endocardial cushion defects
C0014116|T019|AB|745.60|ICD9CM|Endocard cushion def NOS|Endocard cushion def NOS
C0014116|T019|PT|745.60|ICD9CM|Endocardial cushion defect, unspecified type|Endocardial cushion defect, unspecified type
C0031192|T019|AB|745.61|ICD9CM|Ostium primum defect|Ostium primum defect
C0031192|T019|PT|745.61|ICD9CM|Ostium primum defect|Ostium primum defect
C0029608|T019|AB|745.69|ICD9CM|Endocard cushion def NEC|Endocard cushion def NEC
C0029608|T019|PT|745.69|ICD9CM|Other endocardial cushion defects|Other endocardial cushion defects
C0152238|T019|AB|745.7|ICD9CM|Cor biloculare|Cor biloculare
C0152238|T047|AB|745.7|ICD9CM|Cor biloculare|Cor biloculare
C0152238|T019|PT|745.7|ICD9CM|Cor biloculare|Cor biloculare
C0152238|T047|PT|745.7|ICD9CM|Cor biloculare|Cor biloculare
C0158609|T019|PT|745.8|ICD9CM|Other bulbus cordis anomalies and anomalies of cardiac septal closure|Other bulbus cordis anomalies and anomalies of cardiac septal closure
C0158609|T019|AB|745.8|ICD9CM|Septal closure anom NEC|Septal closure anom NEC
C0158610|T019|AB|745.9|ICD9CM|Septal closure anom NOS|Septal closure anom NOS
C0158610|T019|PT|745.9|ICD9CM|Unspecified defect of septal closure|Unspecified defect of septal closure
C0158611|T019|HT|746|ICD9CM|Other congenital anomalies of heart|Other congenital anomalies of heart
C0265830|T019|HT|746.0|ICD9CM|Anomalies of pulmonary valve, congenital|Anomalies of pulmonary valve, congenital
C0265830|T019|PT|746.00|ICD9CM|Congenital pulmonary valve anomaly, unspecified|Congenital pulmonary valve anomaly, unspecified
C0265830|T019|AB|746.00|ICD9CM|Pulmonary valve anom NOS|Pulmonary valve anom NOS
C0242855|T047|PT|746.01|ICD9CM|Atresia of pulmonary valve, congenital|Atresia of pulmonary valve, congenital
C0242855|T047|AB|746.01|ICD9CM|Cong pulmon valv atresia|Cong pulmon valv atresia
C0162164|T019|AB|746.02|ICD9CM|Cong pulmon valve stenos|Cong pulmon valve stenos
C0162164|T019|PT|746.02|ICD9CM|Stenosis of pulmonary valve, congenital|Stenosis of pulmonary valve, congenital
C0477996|T019|PT|746.09|ICD9CM|Other congenital anomalies of pulmonary valve|Other congenital anomalies of pulmonary valve
C0477996|T019|AB|746.09|ICD9CM|Pulmonary valve anom NEC|Pulmonary valve anom NEC
C0158616|T019|AB|746.1|ICD9CM|Cong tricusp atres/sten|Cong tricusp atres/sten
C0158616|T019|PT|746.1|ICD9CM|Tricuspid atresia and stenosis, congenital|Tricuspid atresia and stenosis, congenital
C0013481|T019|AB|746.2|ICD9CM|Ebstein's anomaly|Ebstein's anomaly
C0013481|T019|PT|746.2|ICD9CM|Ebstein's anomaly|Ebstein's anomaly
C0152417|T019|AB|746.3|ICD9CM|Cong aorta valv stenosis|Cong aorta valv stenosis
C0152417|T019|PT|746.3|ICD9CM|Congenital stenosis of aortic valve|Congenital stenosis of aortic valve
C0158617|T047|AB|746.4|ICD9CM|Cong aorta valv insuffic|Cong aorta valv insuffic
C0158617|T047|PT|746.4|ICD9CM|Congenital insufficiency of aortic valve|Congenital insufficiency of aortic valve
C0158618|T019|AB|746.5|ICD9CM|Congen mitral stenosis|Congen mitral stenosis
C0158618|T019|PT|746.5|ICD9CM|Congenital mitral stenosis|Congenital mitral stenosis
C0158619|T019|AB|746.6|ICD9CM|Cong mitral insufficienc|Cong mitral insufficienc
C0158619|T047|AB|746.6|ICD9CM|Cong mitral insufficienc|Cong mitral insufficienc
C0158619|T019|PT|746.6|ICD9CM|Congenital mitral insufficiency|Congenital mitral insufficiency
C0158619|T047|PT|746.6|ICD9CM|Congenital mitral insufficiency|Congenital mitral insufficiency
C0152101|T047|AB|746.7|ICD9CM|Hypoplas left heart synd|Hypoplas left heart synd
C0152101|T047|PT|746.7|ICD9CM|Hypoplastic left heart syndrome|Hypoplastic left heart syndrome
C0477999|T019|HT|746.8|ICD9CM|Other specified congenital anomalies of heart|Other specified congenital anomalies of heart
C0158621|T019|AB|746.81|ICD9CM|Cong subaortic stenosis|Cong subaortic stenosis
C0158621|T019|PT|746.81|ICD9CM|Subaortic stenosis|Subaortic stenosis
C0009995|T019|AB|746.82|ICD9CM|Cor triatriatum|Cor triatriatum
C0009995|T019|PT|746.82|ICD9CM|Cor triatriatum|Cor triatriatum
C0034084|T046|AB|746.83|ICD9CM|Infundib pulmon stenosis|Infundib pulmon stenosis
C0034084|T046|PT|746.83|ICD9CM|Infundibular pulmonic stenosis|Infundibular pulmonic stenosis
C0869419|T019|AB|746.84|ICD9CM|Obstruct heart anom NEC|Obstruct heart anom NEC
C0869419|T019|PT|746.84|ICD9CM|Obstructive anomalies of heart, not elsewhere classified|Obstructive anomalies of heart, not elsewhere classified
C0158623|T019|AB|746.85|ICD9CM|Coronary artery anomaly|Coronary artery anomaly
C0158623|T019|PT|746.85|ICD9CM|Coronary artery anomaly|Coronary artery anomaly
C0149530|T019|AB|746.86|ICD9CM|Congenital heart block|Congenital heart block
C0149530|T047|AB|746.86|ICD9CM|Congenital heart block|Congenital heart block
C0149530|T019|PT|746.86|ICD9CM|Congenital heart block|Congenital heart block
C0149530|T047|PT|746.86|ICD9CM|Congenital heart block|Congenital heart block
C0024649|T019|AB|746.87|ICD9CM|Malposition of heart|Malposition of heart
C0024649|T019|PT|746.87|ICD9CM|Malposition of heart and cardiac apex|Malposition of heart and cardiac apex
C0477999|T019|AB|746.89|ICD9CM|Cong heart anomaly NEC|Cong heart anomaly NEC
C0477999|T019|PT|746.89|ICD9CM|Other specified congenital anomalies of heart|Other specified congenital anomalies of heart
C0018798|T019|AB|746.9|ICD9CM|Cong heart anomaly NOS|Cong heart anomaly NOS
C0018798|T019|PT|746.9|ICD9CM|Unspecified congenital anomaly of heart|Unspecified congenital anomaly of heart
C0158625|T019|HT|747|ICD9CM|Other congenital anomalies of circulatory system|Other congenital anomalies of circulatory system
C0013274|T019|AB|747.0|ICD9CM|Patent ductus arteriosus|Patent ductus arteriosus
C0013274|T019|PT|747.0|ICD9CM|Patent ductus arteriosus|Patent ductus arteriosus
C0003492|T019|HT|747.1|ICD9CM|Coarctation of aorta|Coarctation of aorta
C0003492|T019|AB|747.10|ICD9CM|Coarctation of aorta|Coarctation of aorta
C0003492|T019|PT|747.10|ICD9CM|Coarctation of aorta (preductal) (postductal)|Coarctation of aorta (preductal) (postductal)
C0152419|T019|AB|747.11|ICD9CM|Interrupt of aortic arch|Interrupt of aortic arch
C0152419|T019|PT|747.11|ICD9CM|Interruption of aortic arch|Interruption of aortic arch
C0478000|T019|HT|747.2|ICD9CM|Other congenital anomalies of aorta|Other congenital anomalies of aorta
C0302467|T019|PT|747.20|ICD9CM|Anomaly of aorta, unspecified|Anomaly of aorta, unspecified
C0302467|T019|AB|747.20|ICD9CM|Cong anom of aorta NOS|Cong anom of aorta NOS
C0158629|T019|AB|747.21|ICD9CM|Anomalies of aortic arch|Anomalies of aortic arch
C0158629|T019|PT|747.21|ICD9CM|Anomalies of aortic arch|Anomalies of aortic arch
C0345010|T019|AB|747.22|ICD9CM|Aortic atresia/stenosis|Aortic atresia/stenosis
C0345010|T019|PT|747.22|ICD9CM|Atresia and stenosis of aorta|Atresia and stenosis of aorta
C0478000|T019|AB|747.29|ICD9CM|Cong anom of aorta NEC|Cong anom of aorta NEC
C0478000|T019|PT|747.29|ICD9CM|Other anomalies of aorta|Other anomalies of aorta
C0009681|T019|HT|747.3|ICD9CM|Anomalies of pulmonary artery, congenital|Anomalies of pulmonary artery, congenital
C3161124|T019|AB|747.31|ICD9CM|Pulmon art coarct/atres|Pulmon art coarct/atres
C3161124|T019|PT|747.31|ICD9CM|Pulmonary artery coarctation and atresia|Pulmonary artery coarctation and atresia
C0241790|T019|PT|747.32|ICD9CM|Pulmonary arteriovenous malformation|Pulmonary arteriovenous malformation
C0241790|T019|AB|747.32|ICD9CM|Pulmonary AV malformatn|Pulmonary AV malformatn
C3161125|T019|AB|747.39|ICD9CM|Oth anom pul artery/circ|Oth anom pul artery/circ
C3161125|T019|PT|747.39|ICD9CM|Other anomalies of pulmonary artery and pulmonary circulation|Other anomalies of pulmonary artery and pulmonary circulation
C0158632|T019|HT|747.4|ICD9CM|Anomalies of great veins, congenital|Anomalies of great veins, congenital
C0158632|T019|PT|747.40|ICD9CM|Anomaly of great veins, unspecified|Anomaly of great veins, unspecified
C0158632|T019|AB|747.40|ICD9CM|Great vein anomaly NOS|Great vein anomaly NOS
C4551903|T047|AB|747.41|ICD9CM|Tot anom pulm ven connec|Tot anom pulm ven connec
C4551903|T047|PT|747.41|ICD9CM|Total anomalous pulmonary venous connection|Total anomalous pulmonary venous connection
C0158634|T019|AB|747.42|ICD9CM|Part anom pulm ven conn|Part anom pulm ven conn
C0158634|T019|PT|747.42|ICD9CM|Partial anomalous pulmonary venous connection|Partial anomalous pulmonary venous connection
C0029520|T019|AB|747.49|ICD9CM|Great vein anomaly NEC|Great vein anomaly NEC
C0029520|T019|PT|747.49|ICD9CM|Other anomalies of great veins|Other anomalies of great veins
C0158635|T019|PT|747.5|ICD9CM|Absence or hypoplasia of umbilical artery|Absence or hypoplasia of umbilical artery
C0158635|T019|AB|747.5|ICD9CM|Umbilical artery absence|Umbilical artery absence
C1963536|T019|HT|747.6|ICD9CM|Other congenital anomalies of peripheral vascular system|Other congenital anomalies of peripheral vascular system
C0340797|T019|PT|747.60|ICD9CM|Anomaly of the peripheral vascular system, unspecified site|Anomaly of the peripheral vascular system, unspecified site
C0340797|T019|AB|747.60|ICD9CM|Unsp prpherl vasc anomal|Unsp prpherl vasc anomal
C0375518|T019|PT|747.61|ICD9CM|Gastrointestinal vessel anomaly|Gastrointestinal vessel anomaly
C0375518|T019|AB|747.61|ICD9CM|Gstrontest vesl anomaly|Gstrontest vesl anomaly
C0302468|T019|AB|747.62|ICD9CM|Renal vessel anomaly|Renal vessel anomaly
C0302468|T019|PT|747.62|ICD9CM|Renal vessel anomaly|Renal vessel anomaly
C0375519|T019|PT|747.63|ICD9CM|Upper limb vessel anomaly|Upper limb vessel anomaly
C0375519|T019|AB|747.63|ICD9CM|Upr limb vessel anomaly|Upr limb vessel anomaly
C0375520|T019|PT|747.64|ICD9CM|Lower limb vessel anomaly|Lower limb vessel anomaly
C0375520|T019|AB|747.64|ICD9CM|Lwr limb vessel anomaly|Lwr limb vessel anomaly
C0375521|T019|PT|747.69|ICD9CM|Anomalies of other specified sites of peripheral vascular system|Anomalies of other specified sites of peripheral vascular system
C0375521|T019|AB|747.69|ICD9CM|Oth spcf prph vscl anoml|Oth spcf prph vscl anoml
C0478008|T019|HT|747.8|ICD9CM|Other specified congenital anomalies of circulatory system|Other specified congenital anomalies of circulatory system
C0158638|T019|PT|747.81|ICD9CM|Anomalies of cerebrovascular system|Anomalies of cerebrovascular system
C0158638|T019|AB|747.81|ICD9CM|Cerebrovascular anomaly|Cerebrovascular anomaly
C0375522|T019|AB|747.82|ICD9CM|Spinal vessel anomaly|Spinal vessel anomaly
C0375522|T019|PT|747.82|ICD9CM|Spinal vessel anomaly|Spinal vessel anomaly
C0031190|T047|AB|747.83|ICD9CM|Persistent fetal circ|Persistent fetal circ
C0031190|T047|PT|747.83|ICD9CM|Persistent fetal circulation|Persistent fetal circulation
C0478008|T019|AB|747.89|ICD9CM|Circulatory anomaly NEC|Circulatory anomaly NEC
C0478008|T019|PT|747.89|ICD9CM|Other specified anomalies of circulatory system|Other specified anomalies of circulatory system
C0478013|T019|AB|747.9|ICD9CM|Circulatory anomaly NOS|Circulatory anomaly NOS
C0478013|T019|PT|747.9|ICD9CM|Unspecified anomaly of circulatory system|Unspecified anomaly of circulatory system
C0035238|T019|HT|748|ICD9CM|Anomalies of respiratory system, congenital|Anomalies of respiratory system, congenital
C0008297|T019|AB|748.0|ICD9CM|Choanal atresia|Choanal atresia
C0008297|T019|PT|748.0|ICD9CM|Choanal atresia|Choanal atresia
C0478014|T019|AB|748.1|ICD9CM|Nose anomaly NEC|Nose anomaly NEC
C0478014|T019|PT|748.1|ICD9CM|Other anomalies of nose|Other anomalies of nose
C0281890|T047|AB|748.2|ICD9CM|Laryngeal web|Laryngeal web
C0281890|T047|PT|748.2|ICD9CM|Web of larynx|Web of larynx
C0431510|T019|AB|748.3|ICD9CM|Laryngotrach anomaly NEC|Laryngotrach anomaly NEC
C0431510|T019|PT|748.3|ICD9CM|Other anomalies of larynx, trachea, and bronchus|Other anomalies of larynx, trachea, and bronchus
C0158641|T019|AB|748.4|ICD9CM|Congenital cystic lung|Congenital cystic lung
C0158641|T019|PT|748.4|ICD9CM|Congenital cystic lung|Congenital cystic lung
C0438699|T019|AB|748.5|ICD9CM|Agenesis of lung|Agenesis of lung
C0438699|T019|PT|748.5|ICD9CM|Agenesis, hypoplasia, and dysplasia of lung|Agenesis, hypoplasia, and dysplasia of lung
C0478018|T019|HT|748.6|ICD9CM|Congenital other anomalies of lung|Congenital other anomalies of lung
C0158644|T019|PT|748.60|ICD9CM|Anomaly of lung, unspecified|Anomaly of lung, unspecified
C0158644|T019|AB|748.60|ICD9CM|Lung anomaly NOS|Lung anomaly NOS
C0152239|T019|AB|748.61|ICD9CM|Congen bronchiectasis|Congen bronchiectasis
C0152239|T047|AB|748.61|ICD9CM|Congen bronchiectasis|Congen bronchiectasis
C0152239|T019|PT|748.61|ICD9CM|Congenital bronchiectasis|Congenital bronchiectasis
C0152239|T047|PT|748.61|ICD9CM|Congenital bronchiectasis|Congenital bronchiectasis
C0478018|T019|AB|748.69|ICD9CM|Lung anomaly NEC|Lung anomaly NEC
C0478018|T019|PT|748.69|ICD9CM|Other congenital anomalies of lung|Other congenital anomalies of lung
C0478019|T019|PT|748.8|ICD9CM|Other specified anomalies of respiratory system|Other specified anomalies of respiratory system
C0478019|T019|AB|748.8|ICD9CM|Respiratory anomaly NEC|Respiratory anomaly NEC
C0035238|T019|AB|748.9|ICD9CM|Respiratory anomaly NOS|Respiratory anomaly NOS
C0035238|T019|PT|748.9|ICD9CM|Unspecified anomaly of respiratory system|Unspecified anomaly of respiratory system
C0158646|T019|HT|749|ICD9CM|Cleft palate and cleft lip|Cleft palate and cleft lip
C0008925|T019|HT|749.0|ICD9CM|Cleft palate|Cleft palate
C0008925|T019|AB|749.00|ICD9CM|Cleft palate NOS|Cleft palate NOS
C0008925|T019|PT|749.00|ICD9CM|Cleft palate, unspecified|Cleft palate, unspecified
C0158647|T019|PT|749.01|ICD9CM|Cleft palate, unilateral, complete|Cleft palate, unilateral, complete
C0158647|T019|AB|749.01|ICD9CM|Unilat cleft palate-comp|Unilat cleft palate-comp
C0158648|T019|PT|749.02|ICD9CM|Cleft palate, unilateral, incomplete|Cleft palate, unilateral, incomplete
C0158648|T019|AB|749.02|ICD9CM|Unilat cleft palate-inc|Unilat cleft palate-inc
C0158649|T019|AB|749.03|ICD9CM|Bilat cleft palate-compl|Bilat cleft palate-compl
C0158649|T019|PT|749.03|ICD9CM|Cleft palate, bilateral, complete|Cleft palate, bilateral, complete
C0158650|T019|AB|749.04|ICD9CM|Bilat cleft palate-inc|Bilat cleft palate-inc
C0158650|T019|PT|749.04|ICD9CM|Cleft palate, bilateral, incomplete|Cleft palate, bilateral, incomplete
C0008924|T019|HT|749.1|ICD9CM|Cleft lip|Cleft lip
C0008924|T019|AB|749.10|ICD9CM|Cleft lip NOS|Cleft lip NOS
C0008924|T019|PT|749.10|ICD9CM|Cleft lip, unspecified|Cleft lip, unspecified
C0158651|T019|PT|749.11|ICD9CM|Cleft lip, unilateral, complete|Cleft lip, unilateral, complete
C0158651|T019|AB|749.11|ICD9CM|Unilat cleft lip-compl|Unilat cleft lip-compl
C0158652|T019|PT|749.12|ICD9CM|Cleft lip, unilateral, incomplete|Cleft lip, unilateral, incomplete
C0158652|T019|AB|749.12|ICD9CM|Unilat cleft lip-imcompl|Unilat cleft lip-imcompl
C0158653|T019|AB|749.13|ICD9CM|Bilat cleft lip-complete|Bilat cleft lip-complete
C0158653|T019|PT|749.13|ICD9CM|Cleft lip, bilateral, complete|Cleft lip, bilateral, complete
C0158654|T019|AB|749.14|ICD9CM|Bilat cleft lip-incompl|Bilat cleft lip-incompl
C0158654|T019|PT|749.14|ICD9CM|Cleft lip, bilateral, incomplete|Cleft lip, bilateral, incomplete
C0158646|T019|HT|749.2|ICD9CM|Cleft palate with cleft lip|Cleft palate with cleft lip
C0158646|T019|AB|749.20|ICD9CM|Cleft palate & lip NOS|Cleft palate & lip NOS
C0158646|T019|PT|749.20|ICD9CM|Cleft palate with cleft lip, unspecified|Cleft palate with cleft lip, unspecified
C0158655|T019|PT|749.21|ICD9CM|Cleft palate with cleft lip, unilateral, complete|Cleft palate with cleft lip, unilateral, complete
C0158655|T019|AB|749.21|ICD9CM|Unil cleft palat/lip-com|Unil cleft palat/lip-com
C0158656|T019|PT|749.22|ICD9CM|Cleft palate with cleft lip, unilateral, incomplete|Cleft palate with cleft lip, unilateral, incomplete
C0158656|T019|AB|749.22|ICD9CM|Unil cleft palat/lip-inc|Unil cleft palat/lip-inc
C0158657|T019|AB|749.23|ICD9CM|Bilat clft palat/lip-com|Bilat clft palat/lip-com
C0158657|T019|PT|749.23|ICD9CM|Cleft palate with cleft lip, bilateral, complete|Cleft palate with cleft lip, bilateral, complete
C0158658|T019|AB|749.24|ICD9CM|Bilat clft palat/lip-inc|Bilat clft palat/lip-inc
C0158658|T019|PT|749.24|ICD9CM|Cleft palate with cleft lip, bilateral, incomplete|Cleft palate with cleft lip, bilateral, incomplete
C0158659|T019|AB|749.25|ICD9CM|Cleft palate & lip NEC|Cleft palate & lip NEC
C0158659|T019|PT|749.25|ICD9CM|Other combinations of cleft palate with cleft lip|Other combinations of cleft palate with cleft lip
C2910173|T019|HT|750|ICD9CM|Other congenital anomalies of upper alimentary tract|Other congenital anomalies of upper alimentary tract
C0152415|T019|AB|750.0|ICD9CM|Tongue tie|Tongue tie
C0152415|T019|PT|750.0|ICD9CM|Tongue tie|Tongue tie
C0478024|T019|HT|750.1|ICD9CM|Other congenital anomalies of tongue|Other congenital anomalies of tongue
C0158662|T019|PT|750.10|ICD9CM|Congenital anomaly of tongue, unspecified|Congenital anomaly of tongue, unspecified
C0158662|T019|AB|750.10|ICD9CM|Tongue anomaly NOS|Tongue anomaly NOS
C0158663|T019|AB|750.11|ICD9CM|Aglossia|Aglossia
C0158663|T019|PT|750.11|ICD9CM|Aglossia|Aglossia
C0158664|T019|AB|750.12|ICD9CM|Cong adhesions of tongue|Cong adhesions of tongue
C0158664|T019|PT|750.12|ICD9CM|Congenital adhesions of tongue|Congenital adhesions of tongue
C2349953|T019|AB|750.13|ICD9CM|Cong fissure of tongue|Cong fissure of tongue
C2349953|T019|PT|750.13|ICD9CM|Fissure of tongue|Fissure of tongue
C0009677|T019|AB|750.15|ICD9CM|Cong macroglossia|Cong macroglossia
C0009677|T019|PT|750.15|ICD9CM|Macroglossia|Macroglossia
C0025988|T019|AB|750.16|ICD9CM|Microglossia|Microglossia
C0025988|T019|PT|750.16|ICD9CM|Microglossia|Microglossia
C0478024|T019|PT|750.19|ICD9CM|Other congenital anomalies of tongue|Other congenital anomalies of tongue
C0478024|T019|AB|750.19|ICD9CM|Tongue anomaly NEC|Tongue anomaly NEC
C0431553|T019|HT|750.2|ICD9CM|Other specified congenital anomalies of mouth and pharynx|Other specified congenital anomalies of mouth and pharynx
C0158667|T019|PT|750.21|ICD9CM|Absence of salivary gland|Absence of salivary gland
C0158667|T019|AB|750.21|ICD9CM|Salivary gland absence|Salivary gland absence
C0152429|T019|AB|750.22|ICD9CM|Accessory salivary gland|Accessory salivary gland
C0152429|T019|PT|750.22|ICD9CM|Accessory salivary gland|Accessory salivary gland
C0266118|T019|PT|750.23|ICD9CM|Atresia, salivary duct|Atresia, salivary duct
C0266118|T019|AB|750.23|ICD9CM|Cong atresia, saliv duct|Cong atresia, saliv duct
C0158669|T019|AB|750.24|ICD9CM|Cong salivary fistula|Cong salivary fistula
C0158669|T019|PT|750.24|ICD9CM|Congenital fistula of salivary gland|Congenital fistula of salivary gland
C0158670|T019|PT|750.25|ICD9CM|Congenital fistula of lip|Congenital fistula of lip
C0158670|T019|AB|750.25|ICD9CM|Congenital lip fistula|Congenital lip fistula
C0158671|T019|AB|750.26|ICD9CM|Mouth anomaly NEC|Mouth anomaly NEC
C0158671|T019|PT|750.26|ICD9CM|Other specified anomalies of mouth|Other specified anomalies of mouth
C0392485|T019|AB|750.27|ICD9CM|Diverticulum of pharynx|Diverticulum of pharynx
C0392485|T019|PT|750.27|ICD9CM|Diverticulum of pharynx|Diverticulum of pharynx
C0158673|T019|PT|750.29|ICD9CM|Other specified anomalies of pharynx|Other specified anomalies of pharynx
C0158673|T019|AB|750.29|ICD9CM|Pharyngeal anomaly NEC|Pharyngeal anomaly NEC
C0009733|T019|AB|750.3|ICD9CM|Cong esoph fistula/atres|Cong esoph fistula/atres
C0009733|T019|PT|750.3|ICD9CM|Tracheoesophageal fistula, esophageal atresia and stenosis|Tracheoesophageal fistula, esophageal atresia and stenosis
C0029758|T019|AB|750.4|ICD9CM|Esophageal anomaly NEC|Esophageal anomaly NEC
C0029758|T019|PT|750.4|ICD9CM|Other specified anomalies of esophagus|Other specified anomalies of esophagus
C0700639|T019|AB|750.5|ICD9CM|Cong pyloric stenosis|Cong pyloric stenosis
C0700639|T019|PT|750.5|ICD9CM|Congenital hypertrophic pyloric stenosis|Congenital hypertrophic pyloric stenosis
C0158674|T019|AB|750.6|ICD9CM|Congenital hiatus hernia|Congenital hiatus hernia
C0158674|T019|PT|750.6|ICD9CM|Congenital hiatus hernia|Congenital hiatus hernia
C2004369|T190|AB|750.7|ICD9CM|Gastric anomaly NEC|Gastric anomaly NEC
C2004369|T190|PT|750.7|ICD9CM|Other specified anomalies of stomach|Other specified anomalies of stomach
C0266021|T019|PT|750.8|ICD9CM|Other specified anomalies of upper alimentary tract|Other specified anomalies of upper alimentary tract
C0266021|T019|AB|750.8|ICD9CM|Upper GI anomaly NEC|Upper GI anomaly NEC
C2004465|T019|PT|750.9|ICD9CM|Unspecified anomaly of upper alimentary tract|Unspecified anomaly of upper alimentary tract
C2004465|T019|AB|750.9|ICD9CM|Upper GI anomaly NOS|Upper GI anomaly NOS
C0158678|T019|HT|751|ICD9CM|Other congenital anomalies of digestive system|Other congenital anomalies of digestive system
C0025037|T019|AB|751.0|ICD9CM|Meckel's diverticulum|Meckel's diverticulum
C0025037|T019|PT|751.0|ICD9CM|Meckel's diverticulum|Meckel's diverticulum
C1261176|T019|PT|751.1|ICD9CM|Atresia and stenosis of small intestine|Atresia and stenosis of small intestine
C1261176|T019|AB|751.1|ICD9CM|Atresia small intestine|Atresia small intestine
C0345205|T019|PT|751.2|ICD9CM|Atresia and stenosis of large intestine, rectum, and anal canal|Atresia and stenosis of large intestine, rectum, and anal canal
C0345205|T019|AB|751.2|ICD9CM|Atresia large intestine|Atresia large intestine
C0019570|T019|AB|751.3|ICD9CM|Hirschsprung's disease|Hirschsprung's disease
C0019570|T047|AB|751.3|ICD9CM|Hirschsprung's disease|Hirschsprung's disease
C0019570|T019|PT|751.3|ICD9CM|Hirschsprung's disease and other congenital functional disorders of colon|Hirschsprung's disease and other congenital functional disorders of colon
C0019570|T047|PT|751.3|ICD9CM|Hirschsprung's disease and other congenital functional disorders of colon|Hirschsprung's disease and other congenital functional disorders of colon
C0158679|T019|PT|751.4|ICD9CM|Anomalies of intestinal fixation|Anomalies of intestinal fixation
C0158679|T019|AB|751.4|ICD9CM|Intestinal fixation anom|Intestinal fixation anom
C0555219|T019|AB|751.5|ICD9CM|Intestinal anomaly NEC|Intestinal anomaly NEC
C0555219|T019|PT|751.5|ICD9CM|Other anomalies of intestine|Other anomalies of intestine
C0158681|T019|HT|751.6|ICD9CM|Anomalies of gallbladder, bile ducts, and liver|Anomalies of gallbladder, bile ducts, and liver
C1456424|T019|AB|751.60|ICD9CM|Biliary & liver anom NOS|Biliary & liver anom NOS
C1456424|T019|PT|751.60|ICD9CM|Unspecified anomaly of gallbladder, bile ducts, and liver|Unspecified anomaly of gallbladder, bile ducts, and liver
C0005411|T019|AB|751.61|ICD9CM|Biliary atresia|Biliary atresia
C0005411|T019|PT|751.61|ICD9CM|Biliary atresia|Biliary atresia
C4551631|T047|AB|751.62|ICD9CM|Cong cystic liver dis|Cong cystic liver dis
C4551631|T047|PT|751.62|ICD9CM|Congenital cystic disease of liver|Congenital cystic disease of liver
C0029554|T019|AB|751.69|ICD9CM|Biliary & liver anom NEC|Biliary & liver anom NEC
C0029554|T019|PT|751.69|ICD9CM|Other anomalies of gallbladder, bile ducts, and liver|Other anomalies of gallbladder, bile ducts, and liver
C0158684|T019|PT|751.7|ICD9CM|Anomalies of pancreas|Anomalies of pancreas
C0158684|T019|AB|751.7|ICD9CM|Pancreas anomalies|Pancreas anomalies
C0478039|T019|AB|751.8|ICD9CM|Anom digestive syst NEC|Anom digestive syst NEC
C0478039|T019|PT|751.8|ICD9CM|Other specified anomalies of digestive system|Other specified anomalies of digestive system
C0266015|T019|AB|751.9|ICD9CM|Anom digestive syst NOS|Anom digestive syst NOS
C0266015|T019|PT|751.9|ICD9CM|Unspecified anomaly of digestive system|Unspecified anomaly of digestive system
C0158687|T019|HT|752|ICD9CM|Congenital anomalies of genital organs|Congenital anomalies of genital organs
C0158688|T019|AB|752.0|ICD9CM|Anomalies of ovaries|Anomalies of ovaries
C0158688|T019|PT|752.0|ICD9CM|Anomalies of ovaries|Anomalies of ovaries
C0158689|T019|HT|752.1|ICD9CM|Anomalies of fallopian tubes and broad ligaments, congenital|Anomalies of fallopian tubes and broad ligaments, congenital
C0158689|T019|AB|752.10|ICD9CM|Tubal/broad lig anom NOS|Tubal/broad lig anom NOS
C0158689|T019|PT|752.10|ICD9CM|Unspecified anomaly of fallopian tubes and broad ligaments|Unspecified anomaly of fallopian tubes and broad ligaments
C0013946|T019|AB|752.11|ICD9CM|Embryonic cyst of adnexa|Embryonic cyst of adnexa
C0013946|T019|PT|752.11|ICD9CM|Embryonic cyst of fallopian tubes and broad ligaments|Embryonic cyst of fallopian tubes and broad ligaments
C0478043|T019|PT|752.19|ICD9CM|Other anomalies of fallopian tubes and broad ligaments|Other anomalies of fallopian tubes and broad ligaments
C0478043|T019|AB|752.19|ICD9CM|Tubal/broad lig anom NEC|Tubal/broad lig anom NEC
C0152240|T019|AB|752.2|ICD9CM|Doubling of uterus|Doubling of uterus
C0152240|T019|PT|752.2|ICD9CM|Doubling of uterus|Doubling of uterus
C0431635|T019|HT|752.3|ICD9CM|Other congenital anomalies of uterus|Other congenital anomalies of uterus
C0266384|T019|AB|752.31|ICD9CM|Agenesis of uterus|Agenesis of uterus
C0266384|T019|PT|752.31|ICD9CM|Agenesis of uterus|Agenesis of uterus
C0266399|T019|PT|752.32|ICD9CM|Hypoplasia of uterus|Hypoplasia of uterus
C0266399|T019|AB|752.32|ICD9CM|Hypoplasia of uterus|Hypoplasia of uterus
C0266389|T019|PT|752.33|ICD9CM|Unicornuate uterus|Unicornuate uterus
C0266389|T019|AB|752.33|ICD9CM|Unicornuate uterus|Unicornuate uterus
C0266387|T019|PT|752.34|ICD9CM|Bicornuate uterus|Bicornuate uterus
C0266387|T019|AB|752.34|ICD9CM|Bicornuate uterus|Bicornuate uterus
C0152240|T019|AB|752.35|ICD9CM|Septate uterus|Septate uterus
C0152240|T019|PT|752.35|ICD9CM|Septate uterus|Septate uterus
C0266385|T019|AB|752.36|ICD9CM|Arcuate uterus|Arcuate uterus
C0266385|T019|PT|752.36|ICD9CM|Arcuate uterus|Arcuate uterus
C0431635|T019|AB|752.39|ICD9CM|Anomalies of uterus NEC|Anomalies of uterus NEC
C0431635|T019|PT|752.39|ICD9CM|Other anomalies of uterus|Other anomalies of uterus
C0158694|T019|HT|752.4|ICD9CM|Anomalies of cervix, vagina, and external female genitalia, congenital|Anomalies of cervix, vagina, and external female genitalia, congenital
C0158694|T019|AB|752.40|ICD9CM|Cervix/fem gen anom NOS|Cervix/fem gen anom NOS
C0158694|T019|PT|752.40|ICD9CM|Unspecified anomaly of cervix, vagina, and external female genitalia|Unspecified anomaly of cervix, vagina, and external female genitalia
C0158695|T019|AB|752.41|ICD9CM|Embryon cyst fem gen NEC|Embryon cyst fem gen NEC
C0158695|T019|PT|752.41|ICD9CM|Embryonic cyst of cervix, vagina, and external female genitalia|Embryonic cyst of cervix, vagina, and external female genitalia
C0152436|T019|AB|752.42|ICD9CM|Imperforate hymen|Imperforate hymen
C0152436|T019|PT|752.42|ICD9CM|Imperforate hymen|Imperforate hymen
C0266404|T019|PT|752.43|ICD9CM|Cervical agenesis|Cervical agenesis
C0266404|T019|AB|752.43|ICD9CM|Cervical agenesis|Cervical agenesis
C2921116|T019|PT|752.44|ICD9CM|Cervical duplication|Cervical duplication
C2921116|T019|AB|752.44|ICD9CM|Cervical duplication|Cervical duplication
C1261251|T019|PT|752.45|ICD9CM|Vaginal agenesis|Vaginal agenesis
C1261251|T019|AB|752.45|ICD9CM|Vaginal agenesis|Vaginal agenesis
C1856006|T033|AB|752.46|ICD9CM|Transv vaginal septum|Transv vaginal septum
C1856006|T033|PT|752.46|ICD9CM|Transverse vaginal septum|Transverse vaginal septum
C1841680|T033|AB|752.47|ICD9CM|Longitud vaginal septum|Longitud vaginal septum
C1841680|T033|PT|752.47|ICD9CM|Longitudinal vaginal septum|Longitudinal vaginal septum
C0029553|T019|AB|752.49|ICD9CM|Cervix/fem gen anom NEC|Cervix/fem gen anom NEC
C0029553|T019|PT|752.49|ICD9CM|Other anomalies of cervix, vagina, and external female genitalia|Other anomalies of cervix, vagina, and external female genitalia
C0520578|T019|HT|752.5|ICD9CM|Undescended and retractile testicle|Undescended and retractile testicle
C0010417|T019|AB|752.51|ICD9CM|Undescended testis|Undescended testis
C0010417|T019|PT|752.51|ICD9CM|Undescended testis|Undescended testis
C0520578|T019|AB|752.52|ICD9CM|Retractile testis|Retractile testis
C0520578|T019|PT|752.52|ICD9CM|Retractile testis|Retractile testis
C0375526|T019|HT|752.6|ICD9CM|Hypospadias and epispadias and other penile anomalies|Hypospadias and epispadias and other penile anomalies
C1691215|T019|AB|752.61|ICD9CM|Hypospadias|Hypospadias
C1691215|T019|PT|752.61|ICD9CM|Hypospadias|Hypospadias
C0563449|T019|AB|752.62|ICD9CM|Epispadias|Epispadias
C0563449|T019|PT|752.62|ICD9CM|Epispadias|Epispadias
C0266436|T019|AB|752.63|ICD9CM|Congenital chordee|Congenital chordee
C0266436|T019|PT|752.63|ICD9CM|Congenital chordee|Congenital chordee
C4551492|T019|AB|752.64|ICD9CM|Micropenis|Micropenis
C4551492|T019|PT|752.64|ICD9CM|Micropenis|Micropenis
C0431668|T019|AB|752.65|ICD9CM|Hidden penis|Hidden penis
C0431668|T019|PT|752.65|ICD9CM|Hidden penis|Hidden penis
C0375528|T019|PT|752.69|ICD9CM|Other penile anomalies|Other penile anomalies
C0375528|T019|AB|752.69|ICD9CM|Penile anomalies NEC|Penile anomalies NEC
C0021193|T019|AB|752.7|ICD9CM|Indeterminate sex|Indeterminate sex
C0021193|T019|PT|752.7|ICD9CM|Indeterminate sex and pseudohermaphroditism|Indeterminate sex and pseudohermaphroditism
C0431614|T019|HT|752.8|ICD9CM|Other specified congenital anomalies of genital organs|Other specified congenital anomalies of genital organs
C1260432|T019|AB|752.81|ICD9CM|Scrotal transposition|Scrotal transposition
C1260432|T019|PT|752.81|ICD9CM|Scrotal transposition|Scrotal transposition
C0431614|T019|AB|752.89|ICD9CM|Genital organ anom NEC|Genital organ anom NEC
C0431614|T019|PT|752.89|ICD9CM|Other specified anomalies of genital organs|Other specified anomalies of genital organs
C0158687|T019|AB|752.9|ICD9CM|Genital organ anom NOS|Genital organ anom NOS
C0158687|T019|PT|752.9|ICD9CM|Unspecified anomaly of genital organs|Unspecified anomaly of genital organs
C0158698|T019|HT|753|ICD9CM|Congenital anomalies of urinary system|Congenital anomalies of urinary system
C0158699|T019|AB|753.0|ICD9CM|Renal agenesis|Renal agenesis
C0158699|T019|PT|753.0|ICD9CM|Renal agenesis and dysgenesis|Renal agenesis and dysgenesis
C0311245|T019|HT|753.1|ICD9CM|Cystic kidney disease|Cystic kidney disease
C0311245|T047|HT|753.1|ICD9CM|Cystic kidney disease|Cystic kidney disease
C0311245|T019|AB|753.10|ICD9CM|Cystic kidney diseas NOS|Cystic kidney diseas NOS
C0311245|T047|AB|753.10|ICD9CM|Cystic kidney diseas NOS|Cystic kidney diseas NOS
C0311245|T019|PT|753.10|ICD9CM|Cystic kidney disease, unspecified|Cystic kidney disease, unspecified
C0311245|T047|PT|753.10|ICD9CM|Cystic kidney disease, unspecified|Cystic kidney disease, unspecified
C3854304|T019|AB|753.11|ICD9CM|Congenital renal cyst|Congenital renal cyst
C3854304|T019|PT|753.11|ICD9CM|Congenital single renal cyst|Congenital single renal cyst
C0022680|T047|AB|753.12|ICD9CM|Polycystic kidney NOS|Polycystic kidney NOS
C0022680|T047|PT|753.12|ICD9CM|Polycystic kidney, unspecified type|Polycystic kidney, unspecified type
C0085413|T047|AB|753.13|ICD9CM|Polycyst kid-autosom dom|Polycyst kid-autosom dom
C0085413|T047|PT|753.13|ICD9CM|Polycystic kidney, autosomal dominant|Polycystic kidney, autosomal dominant
C0085548|T047|AB|753.14|ICD9CM|Polycyst kid-autosom rec|Polycyst kid-autosom rec
C0085548|T047|PT|753.14|ICD9CM|Polycystic kidney, autosomal recessive|Polycystic kidney, autosomal recessive
C3536714|T019|AB|753.15|ICD9CM|Renal dysplasia|Renal dysplasia
C3536714|T019|PT|753.15|ICD9CM|Renal dysplasia|Renal dysplasia
C2939174|T047|AB|753.16|ICD9CM|Medullary cystic kidney|Medullary cystic kidney
C2939174|T047|PT|753.16|ICD9CM|Medullary cystic kidney|Medullary cystic kidney
C0022681|T019|AB|753.17|ICD9CM|Medullary sponge kidney|Medullary sponge kidney
C0022681|T047|AB|753.17|ICD9CM|Medullary sponge kidney|Medullary sponge kidney
C0022681|T019|PT|753.17|ICD9CM|Medullary sponge kidney|Medullary sponge kidney
C0022681|T047|PT|753.17|ICD9CM|Medullary sponge kidney|Medullary sponge kidney
C0431705|T019|AB|753.19|ICD9CM|Cystic kidney diseas NEC|Cystic kidney diseas NEC
C0431705|T047|AB|753.19|ICD9CM|Cystic kidney diseas NEC|Cystic kidney diseas NEC
C0431705|T019|PT|753.19|ICD9CM|Other specified cystic kidney disease|Other specified cystic kidney disease
C0431705|T047|PT|753.19|ICD9CM|Other specified cystic kidney disease|Other specified cystic kidney disease
C0431681|T019|HT|753.2|ICD9CM|Obstructive defects of renal pelvis and ureter, congenital|Obstructive defects of renal pelvis and ureter, congenital
C0431681|T019|AB|753.20|ICD9CM|Obs dfct ren plv&urt NOS|Obs dfct ren plv&urt NOS
C0431681|T019|PT|753.20|ICD9CM|Unspecified obstructive defect of renal pelvis and ureter|Unspecified obstructive defect of renal pelvis and ureter
C0375530|T019|AB|753.21|ICD9CM|Congen obst urtroplv jnc|Congen obst urtroplv jnc
C0375530|T019|PT|753.21|ICD9CM|Congenital obstruction of ureteropelvic junction|Congenital obstruction of ureteropelvic junction
C0266332|T019|AB|753.22|ICD9CM|Cong obst ureteroves jnc|Cong obst ureteroves jnc
C0266332|T019|PT|753.22|ICD9CM|Congenital obstruction of ureterovesical junction|Congenital obstruction of ureterovesical junction
C0474873|T019|AB|753.23|ICD9CM|Congenital ureterocele|Congenital ureterocele
C0474873|T019|PT|753.23|ICD9CM|Congenital ureterocele|Congenital ureterocele
C0478056|T019|AB|753.29|ICD9CM|Obst def ren plv&urt NEC|Obst def ren plv&urt NEC
C0478056|T019|PT|753.29|ICD9CM|Other obstructive defects of renal pelvis and ureter|Other obstructive defects of renal pelvis and ureter
C0478058|T019|AB|753.3|ICD9CM|Kidney anomaly NEC|Kidney anomaly NEC
C0478058|T019|PT|753.3|ICD9CM|Other specified anomalies of kidney|Other specified anomalies of kidney
C0431725|T019|PT|753.4|ICD9CM|Other specified anomalies of ureter|Other specified anomalies of ureter
C0431725|T019|AB|753.4|ICD9CM|Ureteral anomaly NEC|Ureteral anomaly NEC
C0005689|T047|AB|753.5|ICD9CM|Bladder exstrophy|Bladder exstrophy
C0005689|T047|PT|753.5|ICD9CM|Exstrophy of urinary bladder|Exstrophy of urinary bladder
C1305964|T019|PT|753.6|ICD9CM|Atresia and stenosis of urethra and bladder neck|Atresia and stenosis of urethra and bladder neck
C1305964|T019|AB|753.6|ICD9CM|Congen urethral stenosis|Congen urethral stenosis
C0431741|T019|AB|753.7|ICD9CM|Anomalies of urachus|Anomalies of urachus
C0431741|T019|PT|753.7|ICD9CM|Anomalies of urachus|Anomalies of urachus
C0158707|T019|AB|753.8|ICD9CM|Cystourethral anom NEC|Cystourethral anom NEC
C0158707|T019|PT|753.8|ICD9CM|Other specified anomalies of bladder and urethra|Other specified anomalies of bladder and urethra
C0158698|T019|PT|753.9|ICD9CM|Unspecified anomaly of urinary system|Unspecified anomaly of urinary system
C0158698|T019|AB|753.9|ICD9CM|Urinary anomaly NOS|Urinary anomaly NOS
C0158709|T019|HT|754|ICD9CM|Certain congenital musculoskeletal deformities|Certain congenital musculoskeletal deformities
C0432068|T019|AB|754.0|ICD9CM|Cong skull/face/jaw def|Cong skull/face/jaw def
C0432068|T019|PT|754.0|ICD9CM|Congenital musculoskeletal deformities of skull, face, and jaw|Congenital musculoskeletal deformities of skull, face, and jaw
C0345380|T019|PT|754.1|ICD9CM|Congenital musculoskeletal deformities of sternocleidomastoid muscle|Congenital musculoskeletal deformities of sternocleidomastoid muscle
C0345380|T019|AB|754.1|ICD9CM|Congenital torticollis|Congenital torticollis
C0158712|T019|AB|754.2|ICD9CM|Cong postural deformity|Cong postural deformity
C0158712|T019|PT|754.2|ICD9CM|Congenital musculoskeletal deformities of spine|Congenital musculoskeletal deformities of spine
C0019555|T019|HT|754.3|ICD9CM|Congenital dislocation of hip|Congenital dislocation of hip
C0009702|T019|AB|754.30|ICD9CM|Cong hip disloc, unilat|Cong hip disloc, unilat
C0009702|T019|PT|754.30|ICD9CM|Congenital dislocation of hip, unilateral|Congenital dislocation of hip, unilateral
C0158713|T019|AB|754.31|ICD9CM|Congen hip disloc, bilat|Congen hip disloc, bilat
C0158713|T019|PT|754.31|ICD9CM|Congenital dislocation of hip, bilateral|Congenital dislocation of hip, bilateral
C1261276|T019|AB|754.32|ICD9CM|Cong hip sublux, unilat|Cong hip sublux, unilat
C1261276|T019|PT|754.32|ICD9CM|Congenital subluxation of hip, unilateral|Congenital subluxation of hip, unilateral
C0158715|T019|AB|754.33|ICD9CM|Cong hip sublux, bilat|Cong hip sublux, bilat
C0158715|T019|PT|754.33|ICD9CM|Congenital subluxation of hip, bilateral|Congenital subluxation of hip, bilateral
C0158716|T019|AB|754.35|ICD9CM|Cong hip disloc w sublux|Cong hip disloc w sublux
C0158716|T019|PT|754.35|ICD9CM|Congenital dislocation of one hip with subluxation of other hip|Congenital dislocation of one hip with subluxation of other hip
C0431946|T019|HT|754.4|ICD9CM|Congenital genu recurvatum and bowing of long bones of leg|Congenital genu recurvatum and bowing of long bones of leg
C0152235|T019|AB|754.40|ICD9CM|Cong genu recurvatum|Cong genu recurvatum
C0152235|T019|PT|754.40|ICD9CM|Genu recurvatum|Genu recurvatum
C0158718|T019|AB|754.41|ICD9CM|Cong knee dislocation|Cong knee dislocation
C0158718|T019|PT|754.41|ICD9CM|Congenital dislocation of knee (with genu recurvatum)|Congenital dislocation of knee (with genu recurvatum)
C0158719|T019|AB|754.42|ICD9CM|Congen bowing of femur|Congen bowing of femur
C0158719|T019|PT|754.42|ICD9CM|Congenital bowing of femur|Congenital bowing of femur
C0158720|T019|AB|754.43|ICD9CM|Cong bowing tibia/fibula|Cong bowing tibia/fibula
C0158720|T019|PT|754.43|ICD9CM|Congenital bowing of tibia and fibula|Congenital bowing of tibia and fibula
C0152432|T019|AB|754.44|ICD9CM|Cong bowing leg NOS|Cong bowing leg NOS
C0152432|T019|PT|754.44|ICD9CM|Congenital bowing of unspecified long bones of leg|Congenital bowing of unspecified long bones of leg
C0158722|T019|HT|754.5|ICD9CM|Varus deformities of feet, congenital|Varus deformities of feet, congenital
C0158722|T019|AB|754.50|ICD9CM|Talipes varus|Talipes varus
C0158722|T019|PT|754.50|ICD9CM|Talipes varus|Talipes varus
C0009081|T019|AB|754.51|ICD9CM|Talipes equinovarus|Talipes equinovarus
C0009081|T019|PT|754.51|ICD9CM|Talipes equinovarus|Talipes equinovarus
C0265649|T019|AB|754.52|ICD9CM|Metatarsus primus varus|Metatarsus primus varus
C0265649|T019|PT|754.52|ICD9CM|Metatarsus primus varus|Metatarsus primus varus
C0265647|T019|AB|754.53|ICD9CM|Metatarsus varus|Metatarsus varus
C0265647|T019|PT|754.53|ICD9CM|Metatarsus varus|Metatarsus varus
C0158725|T019|AB|754.59|ICD9CM|Cong varus foot def NEC|Cong varus foot def NEC
C0158725|T019|PT|754.59|ICD9CM|Other varus deformities of feet|Other varus deformities of feet
C0158726|T019|HT|754.6|ICD9CM|Valgus deformities of feet, congenital|Valgus deformities of feet, congenital
C0152236|T019|AB|754.60|ICD9CM|Talipes valgus|Talipes valgus
C0152236|T019|PT|754.60|ICD9CM|Talipes valgus|Talipes valgus
C0392477|T019|AB|754.61|ICD9CM|Congenital pes planus|Congenital pes planus
C0392477|T019|PT|754.61|ICD9CM|Congenital pes planus|Congenital pes planus
C4551629|T019|PT|754.62|ICD9CM|Talipes calcaneovalgus|Talipes calcaneovalgus
C4551629|T019|AB|754.62|ICD9CM|Talipes calcaneovalgus|Talipes calcaneovalgus
C0158728|T019|AB|754.69|ICD9CM|Cong valgus foot def NEC|Cong valgus foot def NEC
C0158728|T019|PT|754.69|ICD9CM|Other valgus deformities of feet|Other valgus deformities of feet
C0158729|T019|HT|754.7|ICD9CM|Other congenital deformities of feet|Other congenital deformities of feet
C1301937|T019|AB|754.70|ICD9CM|Talipes NOS|Talipes NOS
C1301937|T019|PT|754.70|ICD9CM|Talipes, unspecified|Talipes, unspecified
C0728829|T019|AB|754.71|ICD9CM|Talipes cavus|Talipes cavus
C0728829|T019|PT|754.71|ICD9CM|Talipes cavus|Talipes cavus
C0158729|T019|AB|754.79|ICD9CM|Cong foot deform NEC|Cong foot deform NEC
C0158729|T019|PT|754.79|ICD9CM|Other deformities of feet|Other deformities of feet
C0158730|T019|HT|754.8|ICD9CM|Other specified nonteratogenic anomalies|Other specified nonteratogenic anomalies
C0016842|T019|AB|754.81|ICD9CM|Pectus excavatum|Pectus excavatum
C0016842|T019|PT|754.81|ICD9CM|Pectus excavatum|Pectus excavatum
C0158731|T019|AB|754.82|ICD9CM|Pectus carinatum|Pectus carinatum
C0158731|T019|PT|754.82|ICD9CM|Pectus carinatum|Pectus carinatum
C0158730|T019|AB|754.89|ICD9CM|Nonteratogenic anom NEC|Nonteratogenic anom NEC
C0158730|T019|PT|754.89|ICD9CM|Other specified nonteratogenic anomalies|Other specified nonteratogenic anomalies
C0158732|T019|HT|755|ICD9CM|Other congenital anomalies of limbs|Other congenital anomalies of limbs
C0152427|T019|HT|755.0|ICD9CM|Polydactyly|Polydactyly
C0152427|T019|AB|755.00|ICD9CM|Polydactyly NOS|Polydactyly NOS
C0152427|T019|PT|755.00|ICD9CM|Polydactyly, unspecified digits|Polydactyly, unspecified digits
C0158733|T019|PT|755.01|ICD9CM|Polydactyly of fingers|Polydactyly of fingers
C0158733|T019|AB|755.01|ICD9CM|Polydactyly, fingers|Polydactyly, fingers
C0158734|T019|PT|755.02|ICD9CM|Polydactyly of toes|Polydactyly of toes
C0158734|T019|AB|755.02|ICD9CM|Polydactyly, toes|Polydactyly, toes
C0039075|T019|HT|755.1|ICD9CM|Syndactyly|Syndactyly
C0265553|T019|PT|755.10|ICD9CM|Syndactyly of multiple and unspecified sites|Syndactyly of multiple and unspecified sites
C0265553|T019|AB|755.10|ICD9CM|Syndactyly, multiple/NOS|Syndactyly, multiple/NOS
C0221352|T019|AB|755.11|ICD9CM|Syndactyl fing-no fusion|Syndactyl fing-no fusion
C0221352|T019|PT|755.11|ICD9CM|Syndactyly of fingers without fusion of bone|Syndactyly of fingers without fusion of bone
C0158736|T019|AB|755.12|ICD9CM|Syndactyl fing w fusion|Syndactyl fing w fusion
C0158736|T019|PT|755.12|ICD9CM|Syndactyly of fingers with fusion of bone|Syndactyly of fingers with fusion of bone
C0345377|T019|AB|755.13|ICD9CM|Syndactyl toe-no fusion|Syndactyl toe-no fusion
C0345377|T019|PT|755.13|ICD9CM|Syndactyly of toes without fusion of bone|Syndactyly of toes without fusion of bone
C0158738|T019|AB|755.14|ICD9CM|Syndactyl toe w fusion|Syndactyl toe w fusion
C0158738|T019|PT|755.14|ICD9CM|Syndactyly of toes with fusion of bone|Syndactyly of toes with fusion of bone
C0265566|T019|HT|755.2|ICD9CM|Reduction deformities of upper limb, congenital|Reduction deformities of upper limb, congenital
C0265566|T019|AB|755.20|ICD9CM|Reduc deform up limb NOS|Reduc deform up limb NOS
C0265566|T019|PT|755.20|ICD9CM|Unspecified reduction deformity of upper limb|Unspecified reduction deformity of upper limb
C0431826|T019|AB|755.21|ICD9CM|Transverse defic arm|Transverse defic arm
C0431826|T019|PT|755.21|ICD9CM|Transverse deficiency of upper limb|Transverse deficiency of upper limb
C0375533|T019|AB|755.22|ICD9CM|Longitud defic arm NEC|Longitud defic arm NEC
C0375533|T019|PT|755.22|ICD9CM|Longitudinal deficiency of upper limb, not elsewhere classified|Longitudinal deficiency of upper limb, not elsewhere classified
C0158743|T019|AB|755.23|ICD9CM|Combin longit defic arm|Combin longit defic arm
C0158743|T019|PT|755.23|ICD9CM|Longitudinal deficiency, combined, involving humerus, radius, and ulna (complete or incomplete)|Longitudinal deficiency, combined, involving humerus, radius, and ulna (complete or incomplete)
C0158744|T019|AB|755.24|ICD9CM|Longitudin defic humerus|Longitudin defic humerus
C0158745|T019|AB|755.25|ICD9CM|Longitud defic radioulna|Longitud defic radioulna
C0158746|T019|AB|755.26|ICD9CM|Longitud defic radius|Longitud defic radius
C0158747|T019|AB|755.27|ICD9CM|Longitudinal defic ulna|Longitudinal defic ulna
C0158748|T019|AB|755.28|ICD9CM|Longitudinal defic hand|Longitudinal defic hand
C0490053|T019|AB|755.29|ICD9CM|Longitud defic phalanges|Longitud defic phalanges
C0490053|T019|PT|755.29|ICD9CM|Longitudinal deficiency, phalanges, complete or partial|Longitudinal deficiency, phalanges, complete or partial
C0265618|T019|HT|755.3|ICD9CM|Reduction deformities of lower limb, congenital|Reduction deformities of lower limb, congenital
C0265618|T019|AB|755.30|ICD9CM|Reduction deform leg NOS|Reduction deform leg NOS
C0265618|T019|PT|755.30|ICD9CM|Unspecified reduction deformity of lower limb|Unspecified reduction deformity of lower limb
C0158752|T019|AB|755.31|ICD9CM|Transverse defic leg|Transverse defic leg
C0158752|T019|PT|755.31|ICD9CM|Transverse deficiency of lower limb|Transverse deficiency of lower limb
C0375534|T190|AB|755.32|ICD9CM|Longitudin defic leg NEC|Longitudin defic leg NEC
C0375534|T190|PT|755.32|ICD9CM|Longitudinal deficiency of lower limb, not elsewhere classified|Longitudinal deficiency of lower limb, not elsewhere classified
C0158754|T019|AB|755.33|ICD9CM|Comb longitudin def leg|Comb longitudin def leg
C0158754|T019|PT|755.33|ICD9CM|Longitudinal deficiency, combined, involving femur, tibia, and fibula (complete or incomplete)|Longitudinal deficiency, combined, involving femur, tibia, and fibula (complete or incomplete)
C0158755|T019|AB|755.34|ICD9CM|Longitudinal defic femur|Longitudinal defic femur
C0158756|T019|AB|755.35|ICD9CM|Tibiofibula longit defic|Tibiofibula longit defic
C0158757|T019|AB|755.36|ICD9CM|Longitudinal defic tibia|Longitudinal defic tibia
C0158758|T019|AB|755.37|ICD9CM|Longitudin defic fibula|Longitudin defic fibula
C0158759|T019|AB|755.38|ICD9CM|Longitudinal defic foot|Longitudinal defic foot
C0490054|T019|AB|755.39|ICD9CM|Longitud defic phalanges|Longitud defic phalanges
C0490054|T019|PT|755.39|ICD9CM|Longitudinal deficiency, phalanges, complete or partial|Longitudinal deficiency, phalanges, complete or partial
C0265547|T019|AB|755.4|ICD9CM|Reduct deform limb NOS|Reduct deform limb NOS
C0265547|T019|PT|755.4|ICD9CM|Reduction deformities, unspecified limb|Reduction deformities, unspecified limb
C0478070|T019|HT|755.5|ICD9CM|Other congenital anomalies of upper limb, including shoulder girdle|Other congenital anomalies of upper limb, including shoulder girdle
C0749794|T019|PT|755.50|ICD9CM|Unspecified anomaly of upper limb|Unspecified anomaly of upper limb
C0749794|T019|AB|755.50|ICD9CM|Upper limb anomaly NOS|Upper limb anomaly NOS
C0158760|T019|AB|755.51|ICD9CM|Cong deformity-clavicle|Cong deformity-clavicle
C0158760|T019|PT|755.51|ICD9CM|Congenital deformity of clavicle|Congenital deformity of clavicle
C0152438|T019|AB|755.52|ICD9CM|Cong elevation-scapula|Cong elevation-scapula
C0152438|T019|PT|755.52|ICD9CM|Congenital elevation of scapula|Congenital elevation of scapula
C0158761|T019|AB|755.53|ICD9CM|Radioulnar synostosis|Radioulnar synostosis
C0158761|T019|PT|755.53|ICD9CM|Radioulnar synostosis|Radioulnar synostosis
C0152441|T019|AB|755.54|ICD9CM|Madelung's deformity|Madelung's deformity
C0152441|T019|PT|755.54|ICD9CM|Madelung's deformity|Madelung's deformity
C1510455|T019|AB|755.55|ICD9CM|Acrocephalosyndactyly|Acrocephalosyndactyly
C1510455|T019|PT|755.55|ICD9CM|Acrocephalosyndactyly|Acrocephalosyndactyly
C0265609|T019|AB|755.56|ICD9CM|Accessory carpal bones|Accessory carpal bones
C0265609|T019|PT|755.56|ICD9CM|Accessory carpal bones|Accessory carpal bones
C0158763|T019|AB|755.57|ICD9CM|Macrodactylia (fingers)|Macrodactylia (fingers)
C0158763|T019|PT|755.57|ICD9CM|Macrodactylia (fingers)|Macrodactylia (fingers)
C0265554|T019|PT|755.58|ICD9CM|Cleft hand, congenital|Cleft hand, congenital
C0265554|T019|AB|755.58|ICD9CM|Congenital cleft hand|Congenital cleft hand
C0478070|T019|PT|755.59|ICD9CM|Other anomalies of upper limb, including shoulder girdle|Other anomalies of upper limb, including shoulder girdle
C0478070|T019|AB|755.59|ICD9CM|Upper limb anomaly NEC|Upper limb anomaly NEC
C0478071|T019|HT|755.6|ICD9CM|Other congenital anomalies of lower limb, including pelvic girdle|Other congenital anomalies of lower limb, including pelvic girdle
C0431943|T019|AB|755.60|ICD9CM|Lower limb anomaly NOS|Lower limb anomaly NOS
C0431943|T019|PT|755.60|ICD9CM|Unspecified anomaly of lower limb|Unspecified anomaly of lower limb
C0152430|T019|AB|755.61|ICD9CM|Congenital coxa valga|Congenital coxa valga
C0152430|T019|PT|755.61|ICD9CM|Coxa valga, congenital|Coxa valga, congenital
C0152431|T019|AB|755.62|ICD9CM|Congenital coxa vara|Congenital coxa vara
C0152431|T019|PT|755.62|ICD9CM|Coxa vara, congenital|Coxa vara, congenital
C0029557|T019|AB|755.63|ICD9CM|Cong hip deformity NEC|Cong hip deformity NEC
C0029557|T019|PT|755.63|ICD9CM|Other congenital deformity of hip (joint)|Other congenital deformity of hip (joint)
C0158767|T019|AB|755.64|ICD9CM|Cong knee deformity|Cong knee deformity
C0158767|T019|PT|755.64|ICD9CM|Congenital deformity of knee (joint)|Congenital deformity of knee (joint)
C0158768|T019|AB|755.65|ICD9CM|Macrodactylia of toes|Macrodactylia of toes
C0158768|T019|PT|755.65|ICD9CM|Macrodactylia of toes|Macrodactylia of toes
C0432018|T019|AB|755.66|ICD9CM|Anomalies of toes NEC|Anomalies of toes NEC
C0432018|T019|PT|755.66|ICD9CM|Other anomalies of toes|Other anomalies of toes
C0868868|T019|AB|755.67|ICD9CM|Anomalies of foot NEC|Anomalies of foot NEC
C0868868|T019|PT|755.67|ICD9CM|Anomalies of foot, not elsewhere classified|Anomalies of foot, not elsewhere classified
C0478071|T019|AB|755.69|ICD9CM|Lower limb anomaly NEC|Lower limb anomaly NEC
C0478071|T019|PT|755.69|ICD9CM|Other anomalies of lower limb, including pelvic girdle|Other anomalies of lower limb, including pelvic girdle
C2733636|T019|AB|755.8|ICD9CM|Congen limb anomaly NEC|Congen limb anomaly NEC
C2733636|T019|PT|755.8|ICD9CM|Other specified anomalies of unspecified limb|Other specified anomalies of unspecified limb
C0206762|T019|AB|755.9|ICD9CM|Congen limb anomaly NOS|Congen limb anomaly NOS
C0206762|T019|PT|755.9|ICD9CM|Unspecified anomaly of unspecified limb|Unspecified anomaly of unspecified limb
C0158773|T019|HT|756|ICD9CM|Other congenital musculoskeletal anomalies|Other congenital musculoskeletal anomalies
C0495615|T019|AB|756.0|ICD9CM|Anomal skull/face bones|Anomal skull/face bones
C0495615|T019|PT|756.0|ICD9CM|Anomalies of skull and face bones|Anomalies of skull and face bones
C0158775|T019|HT|756.1|ICD9CM|Anomalies of spine, congenital|Anomalies of spine, congenital
C0158775|T019|AB|756.10|ICD9CM|Anomaly of spine NOS|Anomaly of spine NOS
C0158775|T019|PT|756.10|ICD9CM|Anomaly of spine, unspecified|Anomaly of spine, unspecified
C0432162|T019|AB|756.11|ICD9CM|Lumbosacr spondylolysis|Lumbosacr spondylolysis
C0432162|T019|PT|756.11|ICD9CM|Spondylolysis, lumbosacral region|Spondylolysis, lumbosacral region
C0038017|T019|AB|756.12|ICD9CM|Spondylolisthesis|Spondylolisthesis
C0038017|T019|PT|756.12|ICD9CM|Spondylolisthesis|Spondylolisthesis
C0158776|T019|PT|756.13|ICD9CM|Absence of vertebra, congenital|Absence of vertebra, congenital
C0158776|T019|AB|756.13|ICD9CM|Cong absence of vertebra|Cong absence of vertebra
C0265677|T019|AB|756.14|ICD9CM|Hemivertebra|Hemivertebra
C0265677|T019|PT|756.14|ICD9CM|Hemivertebra|Hemivertebra
C0265678|T019|AB|756.15|ICD9CM|Congen fusion of spine|Congen fusion of spine
C0265678|T019|PT|756.15|ICD9CM|Fusion of spine (vertebra), congenital|Fusion of spine (vertebra), congenital
C0022738|T047|PT|756.16|ICD9CM|Klippel-Feil syndrome|Klippel-Feil syndrome
C0022738|T047|AB|756.16|ICD9CM|Klippel-feil syndrome|Klippel-feil syndrome
C0080174|T019|AB|756.17|ICD9CM|Spina bifida occulta|Spina bifida occulta
C0080174|T019|PT|756.17|ICD9CM|Spina bifida occulta|Spina bifida occulta
C0432138|T019|AB|756.19|ICD9CM|Anomaly of spine NEC|Anomaly of spine NEC
C0432138|T019|PT|756.19|ICD9CM|Other anomalies of spine|Other anomalies of spine
C0158779|T019|AB|756.2|ICD9CM|Cervical rib|Cervical rib
C0158779|T019|PT|756.2|ICD9CM|Cervical rib|Cervical rib
C0432133|T019|PT|756.3|ICD9CM|Other anomalies of ribs and sternum|Other anomalies of ribs and sternum
C0432133|T019|AB|756.3|ICD9CM|Rib & sternum anomal NEC|Rib & sternum anomal NEC
C0008449|T047|AB|756.4|ICD9CM|Chondrodystrophy|Chondrodystrophy
C0008449|T047|PT|756.4|ICD9CM|Chondrodystrophy|Chondrodystrophy
C0375536|T019|HT|756.5|ICD9CM|Congenital osteodystrophies|Congenital osteodystrophies
C0375536|T047|HT|756.5|ICD9CM|Congenital osteodystrophies|Congenital osteodystrophies
C0375536|T019|PT|756.50|ICD9CM|Congenital osteodystrophy, unspecified|Congenital osteodystrophy, unspecified
C0375536|T047|PT|756.50|ICD9CM|Congenital osteodystrophy, unspecified|Congenital osteodystrophy, unspecified
C0375536|T019|AB|756.50|ICD9CM|Osteodystrophy NOS|Osteodystrophy NOS
C0375536|T047|AB|756.50|ICD9CM|Osteodystrophy NOS|Osteodystrophy NOS
C0029434|T047|AB|756.51|ICD9CM|Osteogenesis imperfecta|Osteogenesis imperfecta
C0029434|T047|PT|756.51|ICD9CM|Osteogenesis imperfecta|Osteogenesis imperfecta
C0029454|T047|AB|756.52|ICD9CM|Osteopetrosis|Osteopetrosis
C0029454|T047|PT|756.52|ICD9CM|Osteopetrosis|Osteopetrosis
C0029455|T047|AB|756.53|ICD9CM|Osteopoikilosis|Osteopoikilosis
C0029455|T047|PT|756.53|ICD9CM|Osteopoikilosis|Osteopoikilosis
C0016065|T019|AB|756.54|ICD9CM|Polyostotic fibros dyspl|Polyostotic fibros dyspl
C0016065|T019|PT|756.54|ICD9CM|Polyostotic fibrous dysplasia of bone|Polyostotic fibrous dysplasia of bone
C0013903|T047|AB|756.55|ICD9CM|Chondroectoderm dysplas|Chondroectoderm dysplas
C0013903|T047|PT|756.55|ICD9CM|Chondroectodermal dysplasia|Chondroectodermal dysplasia
C0026760|T019|AB|756.56|ICD9CM|Mult epiphyseal dysplas|Mult epiphyseal dysplas
C0026760|T019|PT|756.56|ICD9CM|Multiple epiphyseal dysplasia|Multiple epiphyseal dysplasia
C0029559|T019|AB|756.59|ICD9CM|Osteodystrophy NEC|Osteodystrophy NEC
C0029559|T019|PT|756.59|ICD9CM|Other osteodystrophies|Other osteodystrophies
C0158782|T019|AB|756.6|ICD9CM|Anomalies of diaphragm|Anomalies of diaphragm
C0158782|T019|PT|756.6|ICD9CM|Anomalies of diaphragm|Anomalies of diaphragm
C0009680|T019|HT|756.7|ICD9CM|Anomalies of abdominal wall, congenital|Anomalies of abdominal wall, congenital
C0009680|T019|PT|756.70|ICD9CM|Anomaly of abdominal wall, unspecified|Anomaly of abdominal wall, unspecified
C0009680|T019|AB|756.70|ICD9CM|Congn anoml abd wall NOS|Congn anoml abd wall NOS
C0033770|T047|AB|756.71|ICD9CM|Prune belly syndrome|Prune belly syndrome
C0033770|T047|PT|756.71|ICD9CM|Prune belly syndrome|Prune belly syndrome
C0795690|T019|PT|756.72|ICD9CM|Omphalocele|Omphalocele
C0795690|T019|AB|756.72|ICD9CM|Omphalocele|Omphalocele
C0265706|T047|AB|756.73|ICD9CM|Gastroschisis|Gastroschisis
C0265706|T047|PT|756.73|ICD9CM|Gastroschisis|Gastroschisis
C0490010|T019|AB|756.79|ICD9CM|Congn anoml abd wall NEC|Congn anoml abd wall NEC
C0490010|T019|PT|756.79|ICD9CM|Other congenital anomalies of abdominal wall|Other congenital anomalies of abdominal wall
C0029759|T019|HT|756.8|ICD9CM|Other specified congenital anomalies of muscle, tendon, fascia, and connective tissue|Other specified congenital anomalies of muscle, tendon, fascia, and connective tissue
C0439002|T019|PT|756.81|ICD9CM|Absence of muscle and tendon|Absence of muscle and tendon
C0439002|T019|AB|756.81|ICD9CM|Absence of muscle/tendon|Absence of muscle/tendon
C0158784|T019|AB|756.82|ICD9CM|Accessory muscle|Accessory muscle
C0158784|T019|PT|756.82|ICD9CM|Accessory muscle|Accessory muscle
C0013720|T047|PT|756.83|ICD9CM|Ehlers-Danlos syndrome|Ehlers-Danlos syndrome
C0013720|T047|AB|756.83|ICD9CM|Ehlers-danlos syndrome|Ehlers-danlos syndrome
C0029759|T019|PT|756.89|ICD9CM|Other specified anomalies of muscle, tendon, fascia, and connective tissue|Other specified anomalies of muscle, tendon, fascia, and connective tissue
C0029759|T019|AB|756.89|ICD9CM|Soft tissue anomaly NEC|Soft tissue anomaly NEC
C0478080|T019|AB|756.9|ICD9CM|Musculoskel anom NEC/NOS|Musculoskel anom NEC/NOS
C0478080|T019|PT|756.9|ICD9CM|Other and unspecified anomalies of musculoskeletal system|Other and unspecified anomalies of musculoskeletal system
C3536895|T019|HT|757|ICD9CM|Congenital anomalies of the integument|Congenital anomalies of the integument
C1313885|T047|AB|757.0|ICD9CM|Hereditary edema of legs|Hereditary edema of legs
C1313885|T047|PT|757.0|ICD9CM|Hereditary edema of legs|Hereditary edema of legs
C0020758|T047|AB|757.1|ICD9CM|Ichthyosis congenita|Ichthyosis congenita
C0020758|T047|PT|757.1|ICD9CM|Ichthyosis congenita|Ichthyosis congenita
C0432333|T019|AB|757.2|ICD9CM|Dermatoglyphic anomalies|Dermatoglyphic anomalies
C0432333|T019|PT|757.2|ICD9CM|Dermatoglyphic anomalies|Dermatoglyphic anomalies
C2363246|T019|HT|757.3|ICD9CM|Other specified congenital anomalies of skin|Other specified congenital anomalies of skin
C0013575|T047|AB|757.31|ICD9CM|Cong ectodermal dysplas|Cong ectodermal dysplas
C0013575|T047|PT|757.31|ICD9CM|Congenital ectodermal dysplasia|Congenital ectodermal dysplasia
C0265973|T019|AB|757.32|ICD9CM|Vascular hamartomas|Vascular hamartomas
C0265973|T019|PT|757.32|ICD9CM|Vascular hamartomas|Vascular hamartomas
C0009726|T019|AB|757.33|ICD9CM|Cong skin pigment anomal|Cong skin pigment anomal
C0009726|T019|PT|757.33|ICD9CM|Congenital pigmentary anomalies of skin|Congenital pigmentary anomalies of skin
C2363246|T019|PT|757.39|ICD9CM|Other specified anomalies of skin|Other specified anomalies of skin
C2363246|T019|AB|757.39|ICD9CM|Skin anomaly NEC|Skin anomaly NEC
C0432340|T019|AB|757.4|ICD9CM|Hair anomalies NEC|Hair anomalies NEC
C0432340|T019|PT|757.4|ICD9CM|Specified anomalies of hair|Specified anomalies of hair
C0432351|T019|AB|757.5|ICD9CM|Nail anomalies NEC|Nail anomalies NEC
C0432351|T019|PT|757.5|ICD9CM|Specified anomalies of nails|Specified anomalies of nails
C0432354|T019|AB|757.6|ICD9CM|Cong breast anomaly NEC|Cong breast anomaly NEC
C0432354|T019|PT|757.6|ICD9CM|Specified congenital anomalies of breast|Specified congenital anomalies of breast
C0478090|T019|AB|757.8|ICD9CM|Oth integument anomalies|Oth integument anomalies
C0478090|T019|PT|757.8|ICD9CM|Other specified anomalies of the integument|Other specified anomalies of the integument
C3536895|T019|AB|757.9|ICD9CM|Integument anomaly NOS|Integument anomaly NOS
C3536895|T019|PT|757.9|ICD9CM|Unspecified congenital anomaly of the integument|Unspecified congenital anomaly of the integument
C0008626|T019|HT|758|ICD9CM|Chromosomal anomalies|Chromosomal anomalies
C0013080|T047|AB|758.0|ICD9CM|Down's syndrome|Down's syndrome
C0013080|T047|PT|758.0|ICD9CM|Down's syndrome|Down's syndrome
C0152095|T047|AB|758.1|ICD9CM|Patau's syndrome|Patau's syndrome
C0152095|T047|PT|758.1|ICD9CM|Patau's syndrome|Patau's syndrome
C0152096|T047|AB|758.2|ICD9CM|Edwards' syndrome|Edwards' syndrome
C0152096|T047|PT|758.2|ICD9CM|Edwards' syndrome|Edwards' syndrome
C0004402|T047|HT|758.3|ICD9CM|Autosomal deletion syndromes|Autosomal deletion syndromes
C0010314|T047|AB|758.31|ICD9CM|Cri-du-chat syndrome|Cri-du-chat syndrome
C0010314|T047|PT|758.31|ICD9CM|Cri-du-chat syndrome|Cri-du-chat syndrome
C0220704|T047|AB|758.32|ICD9CM|Velo-cardio-facial synd|Velo-cardio-facial synd
C0220704|T047|PT|758.32|ICD9CM|Velo-cardio-facial syndrome|Velo-cardio-facial syndrome
C2910371|T047|AB|758.33|ICD9CM|Microdeletions NEC|Microdeletions NEC
C2910371|T047|PT|758.33|ICD9CM|Other microdeletions|Other microdeletions
C0478100|T046|AB|758.39|ICD9CM|Autosomal deletions NEC|Autosomal deletions NEC
C0478100|T046|PT|758.39|ICD9CM|Other autosomal deletions|Other autosomal deletions
C0029549|T047|AB|758.5|ICD9CM|Autosomal anomalies NEC|Autosomal anomalies NEC
C0029549|T047|PT|758.5|ICD9CM|Other conditions due to autosomal anomalies|Other conditions due to autosomal anomalies
C0018051|T019|AB|758.6|ICD9CM|Gonadal dysgenesis|Gonadal dysgenesis
C0018051|T019|PT|758.6|ICD9CM|Gonadal dysgenesis|Gonadal dysgenesis
C0022735|T047|AB|758.7|ICD9CM|Klinefelter's syndrome|Klinefelter's syndrome
C0022735|T047|PT|758.7|ICD9CM|Klinefelter's syndrome|Klinefelter's syndrome
C1305927|T047|HT|758.8|ICD9CM|Other conditions due to chromosome anomalies|Other conditions due to chromosome anomalies
C0029550|T019|AB|758.81|ICD9CM|Oth cond due to sex chrm|Oth cond due to sex chrm
C0029550|T019|PT|758.81|ICD9CM|Other conditions due to sex chromosome anomalies|Other conditions due to sex chromosome anomalies
C1305927|T047|AB|758.89|ICD9CM|Oth con d/t chrm anm NEC|Oth con d/t chrm anm NEC
C1305927|T047|PT|758.89|ICD9CM|Other conditions due to chromosome anomalies|Other conditions due to chromosome anomalies
C0008626|T019|AB|758.9|ICD9CM|Chromosome anomaly NOS|Chromosome anomaly NOS
C0008626|T019|PT|758.9|ICD9CM|Conditions due to anomaly of unspecified chromosome|Conditions due to anomaly of unspecified chromosome
C0158795|T019|HT|759|ICD9CM|Other and unspecified congenital anomalies|Other and unspecified congenital anomalies
C0700587|T019|AB|759.0|ICD9CM|Anomalies of spleen|Anomalies of spleen
C0700587|T019|PT|759.0|ICD9CM|Anomalies of spleen|Anomalies of spleen
C0158797|T019|AB|759.1|ICD9CM|Adrenal gland anomaly|Adrenal gland anomaly
C0158797|T019|PT|759.1|ICD9CM|Anomalies of adrenal gland|Anomalies of adrenal gland
C0432378|T019|PT|759.2|ICD9CM|Anomalies of other endocrine glands|Anomalies of other endocrine glands
C0432378|T019|AB|759.2|ICD9CM|Endocrine anomaly NEC|Endocrine anomaly NEC
C0037221|T019|AB|759.3|ICD9CM|Situs inversus|Situs inversus
C0037221|T019|PT|759.3|ICD9CM|Situs inversus|Situs inversus
C0041428|T019|AB|759.4|ICD9CM|Conjoined twins|Conjoined twins
C0041428|T019|PT|759.4|ICD9CM|Conjoined twins|Conjoined twins
C0041341|T191|AB|759.5|ICD9CM|Tuberous sclerosis|Tuberous sclerosis
C0041341|T191|PT|759.5|ICD9CM|Tuberous sclerosis|Tuberous sclerosis
C0302397|T019|AB|759.6|ICD9CM|Hamartoses NEC|Hamartoses NEC
C0302397|T019|PT|759.6|ICD9CM|Other hamartoses, not elsewhere classified|Other hamartoses, not elsewhere classified
C0026758|T019|AB|759.7|ICD9CM|Mult congen anomal NEC|Mult congen anomal NEC
C0026758|T019|PT|759.7|ICD9CM|Multiple congenital anomalies, so described|Multiple congenital anomalies, so described
C0478095|T019|HT|759.8|ICD9CM|Other specified anomalies|Other specified anomalies
C0032897|T047|PT|759.81|ICD9CM|Prader-Willi syndrome|Prader-Willi syndrome
C0032897|T047|AB|759.81|ICD9CM|Prader-willi syndrome|Prader-willi syndrome
C0024796|T047|AB|759.82|ICD9CM|Marfan syndrome|Marfan syndrome
C0024796|T047|PT|759.82|ICD9CM|Marfan syndrome|Marfan syndrome
C0016667|T047|PT|759.83|ICD9CM|Fragile X syndrome|Fragile X syndrome
C0016667|T047|AB|759.83|ICD9CM|Fragile x syndrome|Fragile x syndrome
C0478095|T019|PT|759.89|ICD9CM|Other specified congenital anomalies|Other specified congenital anomalies
C0478095|T019|AB|759.89|ICD9CM|Specfied cong anomal NEC|Specfied cong anomal NEC
C0000768|T019|AB|759.9|ICD9CM|Congenital anomaly NOS|Congenital anomaly NOS
C0000768|T019|PT|759.9|ICD9CM|Congenital anomaly, unspecified|Congenital anomaly, unspecified
C0158799|T047|HT|760|ICD9CM|Fetus or newborn affected by maternal conditions which may be unrelated to present pregnancy|Fetus or newborn affected by maternal conditions which may be unrelated to present pregnancy
C0178307|T047|HT|760-779.99|ICD9CM|CERTAIN CONDITIONS ORIGINATING IN THE PERINATAL PERIOD|CERTAIN CONDITIONS ORIGINATING IN THE PERINATAL PERIOD
C0411176|T047|AB|760.0|ICD9CM|Matern hyperten aff NB|Matern hyperten aff NB
C0411176|T047|PT|760.0|ICD9CM|Maternal hypertensive disorders affecting fetus or newborn|Maternal hypertensive disorders affecting fetus or newborn
C0158801|T047|AB|760.1|ICD9CM|Matern urine dis aff NB|Matern urine dis aff NB
C0158801|T047|PT|760.1|ICD9CM|Maternal renal and urinary tract diseases affecting fetus or newborn|Maternal renal and urinary tract diseases affecting fetus or newborn
C0411178|T046|AB|760.2|ICD9CM|Maternal infec aff NB|Maternal infec aff NB
C0411178|T046|PT|760.2|ICD9CM|Maternal infections affecting fetus or newborn|Maternal infections affecting fetus or newborn
C0158803|T047|AB|760.3|ICD9CM|Matern cardioresp aff NB|Matern cardioresp aff NB
C0158803|T047|PT|760.3|ICD9CM|Other chronic maternal circulatory and respiratory diseases affecting fetus or newborn|Other chronic maternal circulatory and respiratory diseases affecting fetus or newborn
C0158804|T047|AB|760.4|ICD9CM|Matern nutrit dis aff NB|Matern nutrit dis aff NB
C0158804|T047|PT|760.4|ICD9CM|Maternal nutritional disorders affecting fetus or newborn|Maternal nutritional disorders affecting fetus or newborn
C0158805|T037|AB|760.5|ICD9CM|Maternal injury aff NB|Maternal injury aff NB
C0158805|T037|PT|760.5|ICD9CM|Maternal injury affecting fetus or newborn|Maternal injury affecting fetus or newborn
C2349661|T033|HT|760.6|ICD9CM|Surgical operation on mother and fetus|Surgical operation on mother and fetus
C2349657|T033|AB|760.61|ICD9CM|Amniocentesis affect NB|Amniocentesis affect NB
C2349657|T033|PT|760.61|ICD9CM|Newborn affected by amniocentesis|Newborn affected by amniocentesis
C2349658|T047|AB|760.62|ICD9CM|In utero proc NEC aff NB|In utero proc NEC aff NB
C2349658|T047|PT|760.62|ICD9CM|Newborn affected by other in utero procedure|Newborn affected by other in utero procedure
C2349659|T047|AB|760.63|ICD9CM|Mat surg dur preg aff NB|Mat surg dur preg aff NB
C2349659|T047|PT|760.63|ICD9CM|Newborn affected by other surgical operations on mother during pregnancy|Newborn affected by other surgical operations on mother during pregnancy
C2349660|T033|PT|760.64|ICD9CM|Newborn affected by previous surgical procedure on mother not associated with pregnancy|Newborn affected by previous surgical procedure on mother not associated with pregnancy
C2349660|T033|AB|760.64|ICD9CM|Prev matern surg aff NB|Prev matern surg aff NB
C0859825|T047|HT|760.7|ICD9CM|Noxious influences affecting fetus or newborn via placenta or breast milk|Noxious influences affecting fetus or newborn via placenta or breast milk
C0158808|T047|AB|760.70|ICD9CM|Nox sub NOS aff NB/fetus|Nox sub NOS aff NB/fetus
C0158808|T047|PT|760.70|ICD9CM|Unspecified noxious substance affecting fetus or newborn via placenta or breast milk|Unspecified noxious substance affecting fetus or newborn via placenta or breast milk
C1542327|T033|PT|760.71|ICD9CM|Alcohol affecting fetus or newborn via placenta or breast milk|Alcohol affecting fetus or newborn via placenta or breast milk
C1542327|T033|AB|760.71|ICD9CM|Maternl alc aff NB/fetus|Maternl alc aff NB/fetus
C0158809|T047|AB|760.72|ICD9CM|Matern narc aff NB/fetus|Matern narc aff NB/fetus
C0158809|T047|PT|760.72|ICD9CM|Narcotics affecting fetus or newborn via placenta or breast milk|Narcotics affecting fetus or newborn via placenta or breast milk
C0158810|T033|PT|760.73|ICD9CM|Hallucinogenic agents affecting fetus or newborn via placenta or breast milk|Hallucinogenic agents affecting fetus or newborn via placenta or breast milk
C0158810|T033|AB|760.73|ICD9CM|Matern halluc af NB/fet|Matern halluc af NB/fet
C0158811|T047|PT|760.74|ICD9CM|Anti-infectives affecting fetus or newborn via placenta or breast milk|Anti-infectives affecting fetus or newborn via placenta or breast milk
C0158811|T047|AB|760.74|ICD9CM|Mat anti-inf aff NB/fet|Mat anti-inf aff NB/fet
C0158812|T047|PT|760.75|ICD9CM|Cocaine affecting fetus or newborn via placenta or breast milk|Cocaine affecting fetus or newborn via placenta or breast milk
C0158812|T047|AB|760.75|ICD9CM|Mat cocaine aff NB/fet|Mat cocaine aff NB/fet
C0375539|T047|PT|760.76|ICD9CM|Diethylstilbestrol [DES] affecting fetus or newborn via placenta or breast milk|Diethylstilbestrol [DES] affecting fetus or newborn via placenta or breast milk
C0375539|T047|AB|760.76|ICD9CM|Maternal DES af NB/fetus|Maternal DES af NB/fetus
C1561781|T046|PT|760.77|ICD9CM|Anticonvulsants affecting fetus or newborn via placenta or breast milk|Anticonvulsants affecting fetus or newborn via placenta or breast milk
C1561781|T046|AB|760.77|ICD9CM|Mat anticonv aff NB/fet|Mat anticonv aff NB/fet
C1561786|T046|PT|760.78|ICD9CM|Antimetabolic agents affecting fetus or newborn via placenta or breast milk|Antimetabolic agents affecting fetus or newborn via placenta or breast milk
C1561786|T046|AB|760.78|ICD9CM|Mat antimetabol aff NB|Mat antimetabol aff NB
C0158813|T047|AB|760.79|ICD9CM|Nox sub NEC aff NB/fetus|Nox sub NEC aff NB/fetus
C0158813|T047|PT|760.79|ICD9CM|Other noxious influences affecting fetus or newborn via placenta or breast milk|Other noxious influences affecting fetus or newborn via placenta or breast milk
C0158814|T047|AB|760.8|ICD9CM|Maternal cond NEC aff NB|Maternal cond NEC aff NB
C0158814|T047|PT|760.8|ICD9CM|Other specified maternal conditions affecting fetus or newborn|Other specified maternal conditions affecting fetus or newborn
C0411175|T047|AB|760.9|ICD9CM|Maternal cond NOS aff NB|Maternal cond NOS aff NB
C0411175|T047|PT|760.9|ICD9CM|Unspecified maternal condition affecting fetus or newborn|Unspecified maternal condition affecting fetus or newborn
C0158816|T046|HT|761|ICD9CM|Fetus or newborn affected by maternal complications of pregnancy|Fetus or newborn affected by maternal complications of pregnancy
C0158817|T046|PT|761.0|ICD9CM|Incompetent cervix affecting fetus or newborn|Incompetent cervix affecting fetus or newborn
C0158817|T046|AB|761.0|ICD9CM|Incompetnt cervix aff NB|Incompetnt cervix aff NB
C0411160|T046|AB|761.1|ICD9CM|Premat rupt memb aff NB|Premat rupt memb aff NB
C0411160|T046|PT|761.1|ICD9CM|Premature rupture of membranes affecting fetus or newborn|Premature rupture of membranes affecting fetus or newborn
C0158819|T046|AB|761.2|ICD9CM|Oligohydramnios aff NB|Oligohydramnios aff NB
C0158819|T046|PT|761.2|ICD9CM|Oligohydramnios affecting fetus or newborn|Oligohydramnios affecting fetus or newborn
C0158820|T046|AB|761.3|ICD9CM|Polyhydramnios aff NB|Polyhydramnios aff NB
C0158820|T046|PT|761.3|ICD9CM|Polyhydramnios affecting fetus or newborn|Polyhydramnios affecting fetus or newborn
C0411164|T046|AB|761.4|ICD9CM|Ectopic pregnancy aff NB|Ectopic pregnancy aff NB
C0411164|T046|PT|761.4|ICD9CM|Ectopic pregnancy affecting fetus or newborn|Ectopic pregnancy affecting fetus or newborn
C0411169|T046|AB|761.5|ICD9CM|Mult pregnancy aff NB|Mult pregnancy aff NB
C0411169|T046|PT|761.5|ICD9CM|Multiple pregnancy affecting fetus or newborn|Multiple pregnancy affecting fetus or newborn
C0158823|T046|AB|761.6|ICD9CM|Maternal death aff NB|Maternal death aff NB
C0158823|T046|PT|761.6|ICD9CM|Maternal death affecting fetus or newborn|Maternal death affecting fetus or newborn
C0473867|T046|AB|761.7|ICD9CM|Antepart malpres aff NB|Antepart malpres aff NB
C0473867|T046|PT|761.7|ICD9CM|Malpresentation before labor affecting fetus or newborn|Malpresentation before labor affecting fetus or newborn
C0158825|T047|AB|761.8|ICD9CM|Matern compl NEC aff NB|Matern compl NEC aff NB
C0158825|T047|PT|761.8|ICD9CM|Other specified maternal complications of pregnancy affecting fetus or newborn|Other specified maternal complications of pregnancy affecting fetus or newborn
C0158816|T046|AB|761.9|ICD9CM|Matern compl NOS aff NB|Matern compl NOS aff NB
C0158816|T046|PT|761.9|ICD9CM|Unspecified maternal complication of pregnancy affecting fetus or newborn|Unspecified maternal complication of pregnancy affecting fetus or newborn
C0270025|T046|HT|762|ICD9CM|Fetus or newborn affected by complications of placenta, cord, and membranes|Fetus or newborn affected by complications of placenta, cord, and membranes
C3662231|T033|AB|762.0|ICD9CM|Placenta previa aff NB|Placenta previa aff NB
C3662231|T033|PT|762.0|ICD9CM|Placenta previa affecting fetus or newborn|Placenta previa affecting fetus or newborn
C0158829|T033|PT|762.1|ICD9CM|Other forms of placental separation and hemorrhage affecting fetus or newborn|Other forms of placental separation and hemorrhage affecting fetus or newborn
C0158829|T033|AB|762.1|ICD9CM|Placenta hem NEC aff NB|Placenta hem NEC aff NB
C0477887|T046|AB|762.2|ICD9CM|Abn plac NEC/NOS aff NB|Abn plac NEC/NOS aff NB
C0158831|T046|AB|762.3|ICD9CM|Placent transfusion syn|Placent transfusion syn
C0158831|T046|PT|762.3|ICD9CM|Placental transfusion syndromes affecting fetus or newborn|Placental transfusion syndromes affecting fetus or newborn
C0158832|T046|AB|762.4|ICD9CM|Prolapsed cord aff NB|Prolapsed cord aff NB
C0158832|T046|PT|762.4|ICD9CM|Prolapsed umbilical cord affecting fetus or newborn|Prolapsed umbilical cord affecting fetus or newborn
C0477888|T047|AB|762.5|ICD9CM|Oth umbil cord compress|Oth umbil cord compress
C0477888|T047|PT|762.5|ICD9CM|Other compression of umbilical cord affecting fetus or newborn|Other compression of umbilical cord affecting fetus or newborn
C0477889|T047|PT|762.6|ICD9CM|Other and unspecified conditions of umbilical cord affecting fetus or newborn|Other and unspecified conditions of umbilical cord affecting fetus or newborn
C0477889|T047|AB|762.6|ICD9CM|Umbil cond NEC aff NB|Umbil cond NEC aff NB
C0158835|T046|AB|762.7|ICD9CM|Chorioamnionitis aff NB|Chorioamnionitis aff NB
C0158835|T046|PT|762.7|ICD9CM|Chorioamnionitis affecting fetus or newborn|Chorioamnionitis affecting fetus or newborn
C0158836|T047|AB|762.8|ICD9CM|Abn amnion NEC aff NB|Abn amnion NEC aff NB
C0158836|T047|PT|762.8|ICD9CM|Other specified abnormalities of chorion and amnion affecting fetus or newborn|Other specified abnormalities of chorion and amnion affecting fetus or newborn
C0158837|T047|AB|762.9|ICD9CM|Abn amnion NOS aff NB|Abn amnion NOS aff NB
C0158837|T047|PT|762.9|ICD9CM|Unspecified abnormality of chorion and amnion affecting fetus or newborn|Unspecified abnormality of chorion and amnion affecting fetus or newborn
C0473833|T046|HT|763|ICD9CM|Fetus or newborn affected by other complications of labor and delivery|Fetus or newborn affected by other complications of labor and delivery
C0158839|T047|AB|763.0|ICD9CM|Breech del/extrac aff NB|Breech del/extrac aff NB
C0158839|T047|PT|763.0|ICD9CM|Breech delivery and extraction affecting fetus or newborn|Breech delivery and extraction affecting fetus or newborn
C0477891|T047|AB|763.1|ICD9CM|Malpos/dispro NEC aff NB|Malpos/dispro NEC aff NB
C0158841|T046|AB|763.2|ICD9CM|Forceps delivery aff NB|Forceps delivery aff NB
C0158841|T046|PT|763.2|ICD9CM|Forceps delivery affecting fetus or newborn|Forceps delivery affecting fetus or newborn
C0158842|T033|PT|763.3|ICD9CM|Delivery by vacuum extractor affecting fetus or newborn|Delivery by vacuum extractor affecting fetus or newborn
C0158842|T033|AB|763.3|ICD9CM|Vacuum extrac del aff NB|Vacuum extrac del aff NB
C0158843|T033|AB|763.4|ICD9CM|Cesarean delivery aff NB|Cesarean delivery aff NB
C0158843|T033|PT|763.4|ICD9CM|Cesarean delivery affecting fetus or newborn|Cesarean delivery affecting fetus or newborn
C0495351|T046|AB|763.5|ICD9CM|Mat anesth/analg aff NB|Mat anesth/analg aff NB
C0495351|T046|PT|763.5|ICD9CM|Maternal anesthesia and analgesia affecting fetus or newborn|Maternal anesthesia and analgesia affecting fetus or newborn
C0158845|T046|AB|763.6|ICD9CM|Precipitate del aff NB|Precipitate del aff NB
C0158845|T046|PT|763.6|ICD9CM|Precipitate delivery affecting fetus or newborn|Precipitate delivery affecting fetus or newborn
C0158846|T033|AB|763.7|ICD9CM|Abn uterine contr aff NB|Abn uterine contr aff NB
C0158846|T033|PT|763.7|ICD9CM|Abnormal uterine contractions affecting fetus or newborn|Abnormal uterine contractions affecting fetus or newborn
C0270067|T033|HT|763.8|ICD9CM|Other specified complications of labor and delivery affecting fetus or newborn|Other specified complications of labor and delivery affecting fetus or newborn
C0695249|T046|AB|763.81|ICD9CM|Ab ftl hrt rt/rh b/f lab|Ab ftl hrt rt/rh b/f lab
C0695249|T046|PT|763.81|ICD9CM|Abnormality in fetal heart rate or rhythm before the onset of labor|Abnormality in fetal heart rate or rhythm before the onset of labor
C0695250|T046|AB|763.82|ICD9CM|Ab ftl hrt rt/rh dur lab|Ab ftl hrt rt/rh dur lab
C0695250|T046|PT|763.82|ICD9CM|Abnormality in fetal heart rate or rhythm during labor|Abnormality in fetal heart rate or rhythm during labor
C0695251|T046|AB|763.83|ICD9CM|Ab ftl hrt rt/rhy NOS|Ab ftl hrt rt/rhy NOS
C0695251|T046|PT|763.83|ICD9CM|Abnormality in fetal heart rate or rhythm, unspecified as to time of onset|Abnormality in fetal heart rate or rhythm, unspecified as to time of onset
C1561790|T046|AB|763.84|ICD9CM|Meconium dur del aff NB|Meconium dur del aff NB
C1561790|T046|PT|763.84|ICD9CM|Meconium passage during delivery|Meconium passage during delivery
C0270067|T033|AB|763.89|ICD9CM|Compl del NEC aff NB|Compl del NEC aff NB
C0270067|T033|PT|763.89|ICD9CM|Other specified complications of labor and delivery affecting fetus or newborn|Other specified complications of labor and delivery affecting fetus or newborn
C0495350|T033|AB|763.9|ICD9CM|Compl deliv NOS aff NB|Compl deliv NOS aff NB
C0495350|T033|PT|763.9|ICD9CM|Unspecified complication of labor and delivery affecting fetus or newborn|Unspecified complication of labor and delivery affecting fetus or newborn
C0158849|T033|HT|764|ICD9CM|Slow fetal growth and fetal malnutrition|Slow fetal growth and fetal malnutrition
C0178309|T046|HT|764-779.99|ICD9CM|OTHER CONDITIONS ORIGINATING IN THE PERINATAL PERIOD|OTHER CONDITIONS ORIGINATING IN THE PERINATAL PERIOD
C1313876|T033|HT|764.0|ICD9CM|"Light-for-dates" without mention of fetal malnutrition|"Light-for-dates" without mention of fetal malnutrition
C0158851|T047|PT|764.00|ICD9CM|"Light-for-dates" without mention of fetal malnutrition, unspecified [weight]|"Light-for-dates" without mention of fetal malnutrition, unspecified [weight]
C0158851|T047|AB|764.00|ICD9CM|Light-for-dates wtNOS|Light-for-dates wtNOS
C0158852|T047|PT|764.01|ICD9CM|"Light-for-dates" without mention of fetal malnutrition, less than 500 grams|"Light-for-dates" without mention of fetal malnutrition, less than 500 grams
C0158852|T047|AB|764.01|ICD9CM|Light-for-dates <500g|Light-for-dates <500g
C0158853|T047|PT|764.02|ICD9CM|"Light-for-dates" without mention of fetal malnutrition, 500-749 grams|"Light-for-dates" without mention of fetal malnutrition, 500-749 grams
C0158853|T047|AB|764.02|ICD9CM|Lt-for-dates 500-749g|Lt-for-dates 500-749g
C0158854|T047|PT|764.03|ICD9CM|"Light-for-dates" without mention of fetal malnutrition, 750-999 grams|"Light-for-dates" without mention of fetal malnutrition, 750-999 grams
C0158854|T047|AB|764.03|ICD9CM|Lt-for-dates 750-999g|Lt-for-dates 750-999g
C0158855|T047|PT|764.04|ICD9CM|"Light-for-dates" without mention of fetal malnutrition, 1,000- 1,249 grams|"Light-for-dates" without mention of fetal malnutrition, 1,000- 1,249 grams
C0158855|T047|AB|764.04|ICD9CM|Lt-for-dates 1000-1249g|Lt-for-dates 1000-1249g
C0158856|T047|PT|764.05|ICD9CM|"Light-for-dates"without mention of fetal malnutrition, 1,250- 1,499 grams|"Light-for-dates"without mention of fetal malnutrition, 1,250- 1,499 grams
C0158856|T047|AB|764.05|ICD9CM|Lt-for-dates 1250-1499g|Lt-for-dates 1250-1499g
C0158857|T047|PT|764.06|ICD9CM|"Light-for-dates" without mention of fetal malnutrition, 1,500- 1,749 grams|"Light-for-dates" without mention of fetal malnutrition, 1,500- 1,749 grams
C0158857|T047|AB|764.06|ICD9CM|Lt-for-dates 1500-1749g|Lt-for-dates 1500-1749g
C0158858|T047|PT|764.07|ICD9CM|"Light-for-dates" without mention of fetal malnutrition, 1,750- 1,999 grams|"Light-for-dates" without mention of fetal malnutrition, 1,750- 1,999 grams
C0158858|T047|AB|764.07|ICD9CM|Lt-for-dates 1750-1999g|Lt-for-dates 1750-1999g
C0158859|T047|PT|764.08|ICD9CM|"Light-for-dates" without mention of fetal malnutrition, 2,000- 2,499 grams|"Light-for-dates" without mention of fetal malnutrition, 2,000- 2,499 grams
C0158859|T047|AB|764.08|ICD9CM|Lt-for-dates 2000-2499g|Lt-for-dates 2000-2499g
C0158860|T047|PT|764.09|ICD9CM|"Light-for-dates" without mention of fetal malnutrition, 2,500 grams and over|"Light-for-dates" without mention of fetal malnutrition, 2,500 grams and over
C0158860|T047|AB|764.09|ICD9CM|Lt-for-dates 2500+g|Lt-for-dates 2500+g
C0158861|T047|HT|764.1|ICD9CM|"Light-for-dates" with signs of fetal malnutrition|"Light-for-dates" with signs of fetal malnutrition
C0158862|T047|PT|764.10|ICD9CM|"Light-for-dates" with signs of fetal malnutrition, unspecified [weight]|"Light-for-dates" with signs of fetal malnutrition, unspecified [weight]
C0158862|T047|AB|764.10|ICD9CM|Lt-for-date w/mal wtNOS|Lt-for-date w/mal wtNOS
C0158863|T047|PT|764.11|ICD9CM|"Light-for-dates" with signs of fetal malnutrition, less than 500 grams|"Light-for-dates" with signs of fetal malnutrition, less than 500 grams
C0158863|T047|AB|764.11|ICD9CM|Lt-for-date w/mal <500g|Lt-for-date w/mal <500g
C0158864|T047|PT|764.12|ICD9CM|"Light-for-dates"with signs of fetal malnutrition, 500-749 grams|"Light-for-dates"with signs of fetal malnutrition, 500-749 grams
C0158864|T047|AB|764.12|ICD9CM|Lt-date w/mal 500-749g|Lt-date w/mal 500-749g
C0158865|T047|PT|764.13|ICD9CM|"Light-for-dates" with signs of fetal malnutrition, 750-999 grams|"Light-for-dates" with signs of fetal malnutrition, 750-999 grams
C0158865|T047|AB|764.13|ICD9CM|Lt-date w/mal 750-999g|Lt-date w/mal 750-999g
C0158866|T047|PT|764.14|ICD9CM|"Light-for-dates" with signs of fetal malnutrition, 1,000-1,249 grams|"Light-for-dates" with signs of fetal malnutrition, 1,000-1,249 grams
C0158866|T047|AB|764.14|ICD9CM|Lt-date w/mal 1000-1249g|Lt-date w/mal 1000-1249g
C0158867|T047|PT|764.15|ICD9CM|"Light-for-dates" with signs of fetal malnutrition, 1,250-1,499 grams|"Light-for-dates" with signs of fetal malnutrition, 1,250-1,499 grams
C0158867|T047|AB|764.15|ICD9CM|Lt-date w/mal 1250-1499g|Lt-date w/mal 1250-1499g
C0158868|T047|PT|764.16|ICD9CM|"Light-for-dates" with signs of fetal malnutrition, 1,500-1,749 grams|"Light-for-dates" with signs of fetal malnutrition, 1,500-1,749 grams
C0158868|T047|AB|764.16|ICD9CM|Lt-date w/mal 1500-1749g|Lt-date w/mal 1500-1749g
C0158869|T047|PT|764.17|ICD9CM|"Light-for-dates" with signs of fetal malnutrition, 1,750-1,999 grams|"Light-for-dates" with signs of fetal malnutrition, 1,750-1,999 grams
C0158869|T047|AB|764.17|ICD9CM|Lt-date w/mal 1750-1999g|Lt-date w/mal 1750-1999g
C0158870|T047|PT|764.18|ICD9CM|"Light-for-dates"with signs of fetal malnutrition, 2,000-2,499 grams|"Light-for-dates"with signs of fetal malnutrition, 2,000-2,499 grams
C0158870|T047|AB|764.18|ICD9CM|Lt-date w/mal 2000-2499g|Lt-date w/mal 2000-2499g
C0158871|T047|PT|764.19|ICD9CM|"Light-for-dates"with signs of fetal malnutrition, 2,500 grams and over|"Light-for-dates"with signs of fetal malnutrition, 2,500 grams and over
C0158871|T047|AB|764.19|ICD9CM|Lt-for-date w/mal 2500+g|Lt-for-date w/mal 2500+g
C1510504|T047|HT|764.2|ICD9CM|Fetal malnutrition without mention of "light-for-dates"|Fetal malnutrition without mention of "light-for-dates"
C0158872|T047|PT|764.20|ICD9CM|Fetal malnutrition without mention of "light-for-dates", unspecified [weight]|Fetal malnutrition without mention of "light-for-dates", unspecified [weight]
C0158872|T047|AB|764.20|ICD9CM|Fetal malnutrition wtNOS|Fetal malnutrition wtNOS
C0158873|T047|AB|764.21|ICD9CM|Fetal malnutrition <500g|Fetal malnutrition <500g
C0158873|T047|PT|764.21|ICD9CM|Fetal malnutrition without mention of "light-for-dates", less than 500 grams|Fetal malnutrition without mention of "light-for-dates", less than 500 grams
C0158874|T047|AB|764.22|ICD9CM|Fetal malnutr 500-749g|Fetal malnutr 500-749g
C0158874|T047|PT|764.22|ICD9CM|Fetal malnutrition without mention of "light-for-dates", 500-749 grams|Fetal malnutrition without mention of "light-for-dates", 500-749 grams
C0158875|T047|AB|764.23|ICD9CM|Fetal mal 750-999g|Fetal mal 750-999g
C0158875|T047|PT|764.23|ICD9CM|Fetal malnutrition without mention of "light-for-dates", 750-999 grams|Fetal malnutrition without mention of "light-for-dates", 750-999 grams
C0158876|T047|AB|764.24|ICD9CM|Fetal mal 1000-1249g|Fetal mal 1000-1249g
C0158876|T047|PT|764.24|ICD9CM|Fetal malnutrition without mention of "light-for-dates", 1,000-1,249 grams|Fetal malnutrition without mention of "light-for-dates", 1,000-1,249 grams
C0158877|T047|AB|764.25|ICD9CM|Fetal mal 1250-1499g|Fetal mal 1250-1499g
C0158877|T047|PT|764.25|ICD9CM|Fetal malnutrition without mention of "light-for-dates", 1,250-1,499 grams|Fetal malnutrition without mention of "light-for-dates", 1,250-1,499 grams
C0158878|T047|AB|764.26|ICD9CM|Fetal mal 1500-1749g|Fetal mal 1500-1749g
C0158878|T047|PT|764.26|ICD9CM|Fetal malnutrition without mention of "light-for-dates", 1,500-1,749 grams|Fetal malnutrition without mention of "light-for-dates", 1,500-1,749 grams
C0158879|T047|AB|764.27|ICD9CM|Fetal malnutr 1750-1999g|Fetal malnutr 1750-1999g
C0158879|T047|PT|764.27|ICD9CM|Fetal malnutrition without mention of "light-for-dates", 1,750-1,999 grams|Fetal malnutrition without mention of "light-for-dates", 1,750-1,999 grams
C0158880|T047|AB|764.28|ICD9CM|Fetal malnutr 2000-2499g|Fetal malnutr 2000-2499g
C0158880|T047|PT|764.28|ICD9CM|Fetal malnutrition without mention of "light-for-dates", 2,000-2,499 grams|Fetal malnutrition without mention of "light-for-dates", 2,000-2,499 grams
C0158881|T047|AB|764.29|ICD9CM|Fetal malnutr 2500+g|Fetal malnutr 2500+g
C0158881|T047|PT|764.29|ICD9CM|Fetal malnutrition without mention of "light-for-dates", 2,500 grams and over|Fetal malnutrition without mention of "light-for-dates", 2,500 grams and over
C0015934|T047|HT|764.9|ICD9CM|Fetal growth retardation, unspecified|Fetal growth retardation, unspecified
C0015934|T047|AB|764.90|ICD9CM|Fet growth retard wtNOS|Fet growth retard wtNOS
C0015934|T047|PT|764.90|ICD9CM|Fetal growth retardation, unspecified, unspecified [weight]|Fetal growth retardation, unspecified, unspecified [weight]
C0158883|T047|AB|764.91|ICD9CM|Fet growth retard <500g|Fet growth retard <500g
C0158883|T047|PT|764.91|ICD9CM|Fetal growth retardation, unspecified, less than 500 grams|Fetal growth retardation, unspecified, less than 500 grams
C0158884|T047|AB|764.92|ICD9CM|Fet growth ret 500-749g|Fet growth ret 500-749g
C0158884|T047|PT|764.92|ICD9CM|Fetal growth retardation, unspecified, 500-749 grams|Fetal growth retardation, unspecified, 500-749 grams
C0158885|T047|AB|764.93|ICD9CM|Fet growth ret 750-999g|Fet growth ret 750-999g
C0158885|T047|PT|764.93|ICD9CM|Fetal growth retardation, unspecified, 750-999 grams|Fetal growth retardation, unspecified, 750-999 grams
C0158886|T047|AB|764.94|ICD9CM|Fet grwth ret 1000-1249g|Fet grwth ret 1000-1249g
C0158886|T047|PT|764.94|ICD9CM|Fetal growth retardation, unspecified, 1,000-1,249 grams|Fetal growth retardation, unspecified, 1,000-1,249 grams
C0158887|T047|AB|764.95|ICD9CM|Fet grwth ret 1250-1499g|Fet grwth ret 1250-1499g
C0158887|T047|PT|764.95|ICD9CM|Fetal growth retardation, unspecified, 1,250-1,499 grams|Fetal growth retardation, unspecified, 1,250-1,499 grams
C0158888|T047|AB|764.96|ICD9CM|Fet grwth ret 1500-1749g|Fet grwth ret 1500-1749g
C0158888|T047|PT|764.96|ICD9CM|Fetal growth retardation, unspecified, 1,500-1,749 grams|Fetal growth retardation, unspecified, 1,500-1,749 grams
C0158889|T047|AB|764.97|ICD9CM|Fet grwth ret 1750-1999g|Fet grwth ret 1750-1999g
C0158889|T047|PT|764.97|ICD9CM|Fetal growth retardation, unspecified, 1,750-1,999 grams|Fetal growth retardation, unspecified, 1,750-1,999 grams
C0158890|T047|AB|764.98|ICD9CM|Fet grwth ret 2000-2499g|Fet grwth ret 2000-2499g
C0158890|T047|PT|764.98|ICD9CM|Fetal growth retardation, unspecified, 2,000-2,499 grams|Fetal growth retardation, unspecified, 2,000-2,499 grams
C0158891|T047|AB|764.99|ICD9CM|Fet growth ret 2500+g|Fet growth ret 2500+g
C0158891|T047|PT|764.99|ICD9CM|Fetal growth retardation, unspecified, 2,500 grams and over|Fetal growth retardation, unspecified, 2,500 grams and over
C0158892|T047|HT|765|ICD9CM|Disorders relating to short gestation and unspecified low birthweight|Disorders relating to short gestation and unspecified low birthweight
C0270078|T047|HT|765.0|ICD9CM|Extreme immaturity|Extreme immaturity
C0158894|T047|AB|765.00|ICD9CM|Extreme immatur wtNOS|Extreme immatur wtNOS
C0158894|T047|PT|765.00|ICD9CM|Extreme immaturity, unspecified [weight]|Extreme immaturity, unspecified [weight]
C0158895|T047|AB|765.01|ICD9CM|Extreme immatur <500g|Extreme immatur <500g
C0158895|T047|PT|765.01|ICD9CM|Extreme immaturity, less than 500 grams|Extreme immaturity, less than 500 grams
C0158896|T047|AB|765.02|ICD9CM|Extreme immatur 500-749g|Extreme immatur 500-749g
C0158896|T047|PT|765.02|ICD9CM|Extreme immaturity, 500-749 grams|Extreme immaturity, 500-749 grams
C0158897|T047|AB|765.03|ICD9CM|Extreme immatur 750-999g|Extreme immatur 750-999g
C0158897|T047|PT|765.03|ICD9CM|Extreme immaturity, 750-999 grams|Extreme immaturity, 750-999 grams
C0158898|T047|AB|765.04|ICD9CM|Extreme immat 1000-1249g|Extreme immat 1000-1249g
C0158898|T047|PT|765.04|ICD9CM|Extreme immaturity, 1,000-1,249 grams|Extreme immaturity, 1,000-1,249 grams
C0158899|T047|AB|765.05|ICD9CM|Extreme immat 1250-1499g|Extreme immat 1250-1499g
C0158899|T047|PT|765.05|ICD9CM|Extreme immaturity, 1,250-1,499 grams|Extreme immaturity, 1,250-1,499 grams
C0158900|T047|AB|765.06|ICD9CM|Extreme immat 1500-1749g|Extreme immat 1500-1749g
C0158900|T047|PT|765.06|ICD9CM|Extreme immaturity, 1,500-1,749 grams|Extreme immaturity, 1,500-1,749 grams
C0158901|T047|AB|765.07|ICD9CM|Extreme immat 1750-1999g|Extreme immat 1750-1999g
C0158901|T047|PT|765.07|ICD9CM|Extreme immaturity, 1,750-1,999 grams|Extreme immaturity, 1,750-1,999 grams
C0158902|T047|AB|765.08|ICD9CM|Extreme immat 2000-2499g|Extreme immat 2000-2499g
C0158902|T047|PT|765.08|ICD9CM|Extreme immaturity, 2,000-2,499 grams|Extreme immaturity, 2,000-2,499 grams
C0158903|T047|AB|765.09|ICD9CM|Extreme immat 2500+g|Extreme immat 2500+g
C0158903|T047|PT|765.09|ICD9CM|Extreme immaturity, 2,500 grams and over|Extreme immaturity, 2,500 grams and over
C0029713|T047|HT|765.1|ICD9CM|Other preterm infants|Other preterm infants
C0029713|T047|PT|765.10|ICD9CM|Other preterm infants, unspecified [weight]|Other preterm infants, unspecified [weight]
C0029713|T047|AB|765.10|ICD9CM|Preterm infant NEC wtNOS|Preterm infant NEC wtNOS
C1135241|T033|HT|765.2|ICD9CM|Weeks of gestation|Weeks of gestation
C1135241|T033|PT|765.20|ICD9CM|Unspecified weeks of gestation|Unspecified weeks of gestation
C1135241|T033|AB|765.20|ICD9CM|Weeks of gestation NOS|Weeks of gestation NOS
C0730521|T033|AB|765.21|ICD9CM|<24 comp wks gestation|<24 comp wks gestation
C0730521|T033|PT|765.21|ICD9CM|Less than 24 completed weeks of gestation|Less than 24 completed weeks of gestation
C0730522|T033|AB|765.22|ICD9CM|24 comp weeks gestation|24 comp weeks gestation
C0730522|T033|PT|765.22|ICD9CM|24 completed weeks of gestation|24 completed weeks of gestation
C1135242|T033|AB|765.23|ICD9CM|25-26 comp wks gestation|25-26 comp wks gestation
C1135242|T033|PT|765.23|ICD9CM|25-26 completed weeks of gestation|25-26 completed weeks of gestation
C1135243|T033|AB|765.24|ICD9CM|27-28 comp wks gestation|27-28 comp wks gestation
C1135243|T033|PT|765.24|ICD9CM|27-28 completed weeks of gestation|27-28 completed weeks of gestation
C1135244|T033|AB|765.25|ICD9CM|29-30 comp wks gestation|29-30 comp wks gestation
C1135244|T033|PT|765.25|ICD9CM|29-30 completed weeks of gestation|29-30 completed weeks of gestation
C1135245|T037|AB|765.26|ICD9CM|31-32 comp wks gestation|31-32 comp wks gestation
C1135245|T037|PT|765.26|ICD9CM|31-32 completed weeks of gestation|31-32 completed weeks of gestation
C1135246|T033|AB|765.27|ICD9CM|33-34 comp wks gestation|33-34 comp wks gestation
C1135246|T033|PT|765.27|ICD9CM|33-34 completed weeks of gestation|33-34 completed weeks of gestation
C1135247|T033|AB|765.28|ICD9CM|35-36 comp wks gestation|35-36 comp wks gestation
C1135247|T033|PT|765.28|ICD9CM|35-36 completed weeks of gestation|35-36 completed weeks of gestation
C1135248|T047|PT|765.29|ICD9CM|37 or more completed weeks of gestation|37 or more completed weeks of gestation
C1135248|T047|AB|765.29|ICD9CM|37+ comp wks gestation|37+ comp wks gestation
C0158914|T047|HT|766|ICD9CM|Disorders relating to long gestation and high birthweight|Disorders relating to long gestation and high birthweight
C2242834|T033|AB|766.0|ICD9CM|Exceptionally large baby|Exceptionally large baby
C2242834|T033|PT|766.0|ICD9CM|Exceptionally large baby|Exceptionally large baby
C0477897|T047|AB|766.1|ICD9CM|Heavy-for-date infan NEC|Heavy-for-date infan NEC
C0477897|T047|PT|766.1|ICD9CM|Other "heavy-for-dates" infants|Other "heavy-for-dates" infants
C0158917|T047|HT|766.2|ICD9CM|Late infant, not "heavy-for-dates"|Late infant, not "heavy-for-dates"
C2909960|T046|AB|766.22|ICD9CM|Prolong gestation-infant|Prolong gestation-infant
C2909960|T046|PT|766.22|ICD9CM|Prolonged gestation of infant|Prolonged gestation of infant
C0005604|T037|HT|767|ICD9CM|Birth trauma|Birth trauma
C0836917|T046|AB|767.0|ICD9CM|Cerebral hem at birth|Cerebral hem at birth
C0836917|T046|PT|767.0|ICD9CM|Subdural and cerebral hemorrhage|Subdural and cerebral hemorrhage
C0270089|T037|HT|767.1|ICD9CM|Injuries to scalp due to birth trauma|Injuries to scalp due to birth trauma
C0270092|T046|AB|767.11|ICD9CM|Epicranial subapo hemorr|Epicranial subapo hemorr
C0270092|T046|PT|767.11|ICD9CM|Epicranial subaponeurotic hemorrhage (massive)|Epicranial subaponeurotic hemorrhage (massive)
C1260437|T037|AB|767.19|ICD9CM|Injuries to scalp NEC|Injuries to scalp NEC
C1260437|T037|PT|767.19|ICD9CM|Other injuries to scalp|Other injuries to scalp
C0270094|T037|AB|767.2|ICD9CM|Clavicle fx at birth|Clavicle fx at birth
C0270094|T037|PT|767.2|ICD9CM|Fracture of clavicle due to birth trauma|Fracture of clavicle due to birth trauma
C0700643|T037|AB|767.3|ICD9CM|Bone injury NEC at birth|Bone injury NEC at birth
C0700643|T037|PT|767.3|ICD9CM|Other injuries to skeleton due to birth trauma|Other injuries to skeleton due to birth trauma
C0411063|T037|PT|767.4|ICD9CM|Injury to spine and spinal cord due to birth trauma|Injury to spine and spinal cord due to birth trauma
C0411063|T037|AB|767.4|ICD9CM|Spinal cord inj at birth|Spinal cord inj at birth
C0270103|T037|AB|767.5|ICD9CM|Facial nerve inj-birth|Facial nerve inj-birth
C0270103|T037|PT|767.5|ICD9CM|Facial nerve injury due to birth trauma|Facial nerve injury due to birth trauma
C0270105|T037|AB|767.6|ICD9CM|Brach plexus inj-birth|Brach plexus inj-birth
C0270105|T037|PT|767.6|ICD9CM|Injury to brachial plexus due to birth trauma|Injury to brachial plexus due to birth trauma
C0158925|T037|AB|767.7|ICD9CM|Nerve inj NEC at birth|Nerve inj NEC at birth
C0158925|T037|PT|767.7|ICD9CM|Other cranial and peripheral nerve injuries due to birth trauma|Other cranial and peripheral nerve injuries due to birth trauma
C0477903|T037|AB|767.8|ICD9CM|Birth trauma NEC|Birth trauma NEC
C0477903|T037|PT|767.8|ICD9CM|Other specified birth trauma|Other specified birth trauma
C0005604|T037|AB|767.9|ICD9CM|Birth trauma NOS|Birth trauma NOS
C0005604|T037|PT|767.9|ICD9CM|Birth trauma, unspecified|Birth trauma, unspecified
C2003945|T047|HT|768|ICD9CM|Intrauterine hypoxia and birth asphyxia|Intrauterine hypoxia and birth asphyxia
C0270131|T046|PT|768.0|ICD9CM|Fetal death from asphyxia or anoxia before onset of labor or at unspecified time|Fetal death from asphyxia or anoxia before onset of labor or at unspecified time
C0270131|T046|AB|768.0|ICD9CM|Fetal death-anoxia NOS|Fetal death-anoxia NOS
C0158928|T046|AB|768.1|ICD9CM|Fet death-anoxia dur lab|Fet death-anoxia dur lab
C0158928|T046|PT|768.1|ICD9CM|Fetal death from asphyxia or anoxia during labor|Fetal death from asphyxia or anoxia during labor
C0158929|T046|AB|768.2|ICD9CM|Fet distress befor labor|Fet distress befor labor
C0158929|T046|PT|768.2|ICD9CM|Fetal distress before onset of labor, in liveborn infant|Fetal distress before onset of labor, in liveborn infant
C1719625|T046|PT|768.3|ICD9CM|Fetal distress first noted during labor and delivery, in liveborn infant|Fetal distress first noted during labor and delivery, in liveborn infant
C1719625|T046|AB|768.3|ICD9CM|Fetal distrs dur lab/del|Fetal distrs dur lab/del
C0270124|T047|AB|768.4|ICD9CM|Fetal distress NOS|Fetal distress NOS
C0270124|T047|PT|768.4|ICD9CM|Fetal distress, unspecified as to time of onset, in liveborn infant|Fetal distress, unspecified as to time of onset, in liveborn infant
C0158931|T046|AB|768.5|ICD9CM|Severe birth asphyxia|Severe birth asphyxia
C0158931|T046|PT|768.5|ICD9CM|Severe birth asphyxia|Severe birth asphyxia
C0456089|T046|PT|768.6|ICD9CM|Mild or moderate birth asphyxia|Mild or moderate birth asphyxia
C0456089|T046|AB|768.6|ICD9CM|Mild/mod birth asphyxia|Mild/mod birth asphyxia
C0752304|T047|HT|768.7|ICD9CM|Hypoxic-ischemic encephalopathy (HIE)|Hypoxic-ischemic encephalopathy (HIE)
C0752304|T047|AB|768.70|ICD9CM|Hypoxc-ischem enceph NOS|Hypoxc-ischem enceph NOS
C0752304|T047|PT|768.70|ICD9CM|Hypoxic-ischemic encephalopathy, unspecified|Hypoxic-ischemic encephalopathy, unspecified
C2712358|T047|AB|768.71|ICD9CM|Mild hypox-ischem enceph|Mild hypox-ischem enceph
C2712358|T047|PT|768.71|ICD9CM|Mild hypoxic-ischemic encephalopathy|Mild hypoxic-ischemic encephalopathy
C2712359|T047|AB|768.72|ICD9CM|Mod hypox-ischem enceph|Mod hypox-ischem enceph
C2712359|T047|PT|768.72|ICD9CM|Moderate hypoxic-ischemic encephalopathy|Moderate hypoxic-ischemic encephalopathy
C2712360|T047|AB|768.73|ICD9CM|Sev hypox-ischem enceph|Sev hypox-ischem enceph
C2712360|T047|PT|768.73|ICD9CM|Severe hypoxic-ischemic encephalopathy|Severe hypoxic-ischemic encephalopathy
C0004045|T047|AB|768.9|ICD9CM|Birth asphyxia NOS|Birth asphyxia NOS
C0004045|T047|PT|768.9|ICD9CM|Unspecified severity of birth asphyxia in liveborn infant|Unspecified severity of birth asphyxia in liveborn infant
C0035220|T047|AB|769|ICD9CM|Respiratory distress syn|Respiratory distress syn
C0035220|T047|PT|769|ICD9CM|Respiratory distress syndrome in newborn|Respiratory distress syndrome in newborn
C0158934|T047|HT|770|ICD9CM|Other respiratory conditions of fetus and newborn|Other respiratory conditions of fetus and newborn
C0158935|T047|AB|770.0|ICD9CM|Congenital pneumonia|Congenital pneumonia
C0158935|T047|PT|770.0|ICD9CM|Congenital pneumonia|Congenital pneumonia
C1561805|T046|HT|770.1|ICD9CM|Fetal and newborn aspiration|Fetal and newborn aspiration
C1561791|T046|AB|770.10|ICD9CM|Fetal & newborn asp NOS|Fetal & newborn asp NOS
C1561791|T046|PT|770.10|ICD9CM|Fetal and newborn aspiration, unspecified|Fetal and newborn aspiration, unspecified
C1561792|T046|AB|770.11|ICD9CM|Meconium asp wo resp sym|Meconium asp wo resp sym
C1561792|T046|PT|770.11|ICD9CM|Meconium aspiration without respiratory symptoms|Meconium aspiration without respiratory symptoms
C1561793|T046|AB|770.12|ICD9CM|Meconium asp w resp symp|Meconium asp w resp symp
C1561793|T046|PT|770.12|ICD9CM|Meconium aspiration with respiratory symptoms|Meconium aspiration with respiratory symptoms
C1561794|T046|AB|770.13|ICD9CM|Amniotc asp w/o resp sym|Amniotc asp w/o resp sym
C1561794|T046|PT|770.13|ICD9CM|Aspiration of clear amniotic fluid without respiratory symptoms|Aspiration of clear amniotic fluid without respiratory symptoms
C1561796|T046|AB|770.14|ICD9CM|Amniotic asp w resp sym|Amniotic asp w resp sym
C1561796|T046|PT|770.14|ICD9CM|Aspiration of clear amniotic fluid with respiratory symptoms|Aspiration of clear amniotic fluid with respiratory symptoms
C1561799|T046|PT|770.15|ICD9CM|Aspiration of blood without respiratory symptoms|Aspiration of blood without respiratory symptoms
C1561799|T046|AB|770.15|ICD9CM|Blood asp w/o resp sympt|Blood asp w/o resp sympt
C1561800|T046|PT|770.16|ICD9CM|Aspiration of blood with respiratory symptoms|Aspiration of blood with respiratory symptoms
C1561800|T046|AB|770.16|ICD9CM|Blood asp w resp sympt|Blood asp w resp sympt
C1561801|T046|AB|770.17|ICD9CM|NB asp w/o resp symp NEC|NB asp w/o resp symp NEC
C1561801|T046|PT|770.17|ICD9CM|Other fetal and newborn aspiration without respiratory symptoms|Other fetal and newborn aspiration without respiratory symptoms
C1561802|T046|AB|770.18|ICD9CM|NB asp w resp symp NEC|NB asp w resp symp NEC
C1561802|T046|PT|770.18|ICD9CM|Other fetal and newborn aspiration with respiratory symptoms|Other fetal and newborn aspiration with respiratory symptoms
C0158936|T047|PT|770.2|ICD9CM|Interstitial emphysema and related conditions|Interstitial emphysema and related conditions
C0158936|T047|AB|770.2|ICD9CM|NB interstit emphysema|NB interstit emphysema
C0475713|T046|AB|770.3|ICD9CM|NB pulmonary hemorrhage|NB pulmonary hemorrhage
C0475713|T046|PT|770.3|ICD9CM|Pulmonary hemorrhage|Pulmonary hemorrhage
C0270163|T046|AB|770.4|ICD9CM|Primary atelectasis|Primary atelectasis
C0270163|T046|PT|770.4|ICD9CM|Primary atelectasis|Primary atelectasis
C0158939|T047|AB|770.5|ICD9CM|NB atelectasis NEC/NOS|NB atelectasis NEC/NOS
C0158939|T047|PT|770.5|ICD9CM|Other and unspecified atelectasis|Other and unspecified atelectasis
C0158940|T047|AB|770.6|ICD9CM|NB transitory tachypnea|NB transitory tachypnea
C0158940|T047|PT|770.6|ICD9CM|Transitory tachypnea of newborn|Transitory tachypnea of newborn
C0456017|T047|PT|770.7|ICD9CM|Chronic respiratory disease arising in the perinatal period|Chronic respiratory disease arising in the perinatal period
C0456017|T047|AB|770.7|ICD9CM|Perinatal chr resp dis|Perinatal chr resp dis
C0158942|T047|HT|770.8|ICD9CM|Other newborn respiratory problems|Other newborn respiratory problems
C2316590|T047|AB|770.81|ICD9CM|Primary apnea of newborn|Primary apnea of newborn
C2316590|T047|PT|770.81|ICD9CM|Primary apnea of newborn|Primary apnea of newborn
C0477914|T046|AB|770.82|ICD9CM|Other apnea of newborn|Other apnea of newborn
C0477914|T046|PT|770.82|ICD9CM|Other apnea of newborn|Other apnea of newborn
C0270148|T047|AB|770.83|ICD9CM|Cyanotic attack, newborn|Cyanotic attack, newborn
C0270148|T047|PT|770.83|ICD9CM|Cyanotic attacks of newborn|Cyanotic attacks of newborn
C0521648|T047|AB|770.84|ICD9CM|Resp failure of newborn|Resp failure of newborn
C0521648|T047|PT|770.84|ICD9CM|Respiratory failure of newborn|Respiratory failure of newborn
C1561806|T046|PT|770.85|ICD9CM|Aspiration of postnatal stomach contents without respiratory symptoms|Aspiration of postnatal stomach contents without respiratory symptoms
C1561806|T046|AB|770.85|ICD9CM|Stomch cont asp w/o resp|Stomch cont asp w/o resp
C1561808|T046|PT|770.86|ICD9CM|Aspiration of postnatal stomach contents with respiratory symptoms|Aspiration of postnatal stomach contents with respiratory symptoms
C1561808|T046|AB|770.86|ICD9CM|Stomach cont asp w resp|Stomach cont asp w resp
C0235065|T046|AB|770.87|ICD9CM|NB respiratory arrest|NB respiratory arrest
C0235065|T046|PT|770.87|ICD9CM|Respiratory arrest of newborn|Respiratory arrest of newborn
C2316692|T047|PT|770.88|ICD9CM|Hypoxemia of newborn|Hypoxemia of newborn
C2316692|T047|AB|770.88|ICD9CM|NB hypoxia|NB hypoxia
C1135250|T047|PT|770.89|ICD9CM|Other respiratory problems after birth|Other respiratory problems after birth
C1135250|T047|AB|770.89|ICD9CM|Resp prob after brth NEC|Resp prob after brth NEC
C0270146|T047|AB|770.9|ICD9CM|NB respiratory cond NOS|NB respiratory cond NOS
C0270146|T047|PT|770.9|ICD9CM|Unspecified respiratory condition of fetus and newborn|Unspecified respiratory condition of fetus and newborn
C0158944|T047|HT|771|ICD9CM|Infections specific to the perinatal period|Infections specific to the perinatal period
C0035921|T047|AB|771.0|ICD9CM|Congenital rubella|Congenital rubella
C0035921|T047|PT|771.0|ICD9CM|Congenital rubella|Congenital rubella
C0158945|T047|AB|771.1|ICD9CM|Cong cytomegalovirus inf|Cong cytomegalovirus inf
C0158945|T047|PT|771.1|ICD9CM|Congenital cytomegalovirus infection|Congenital cytomegalovirus infection
C0158946|T047|AB|771.2|ICD9CM|Congenital infec NEC|Congenital infec NEC
C0158946|T047|PT|771.2|ICD9CM|Other congenital infections specific to the perinatal period|Other congenital infections specific to the perinatal period
C0343312|T047|AB|771.3|ICD9CM|Tetanus neonatorum|Tetanus neonatorum
C0343312|T047|PT|771.3|ICD9CM|Tetanus neonatorum|Tetanus neonatorum
C0158947|T047|AB|771.4|ICD9CM|Omphalitis of newborn|Omphalitis of newborn
C0158947|T047|PT|771.4|ICD9CM|Omphalitis of the newborn|Omphalitis of the newborn
C0158948|T047|AB|771.5|ICD9CM|Neonatal infec mastitis|Neonatal infec mastitis
C0158948|T047|PT|771.5|ICD9CM|Neonatal infective mastitis|Neonatal infective mastitis
C0027611|T047|AB|771.6|ICD9CM|Neonatal conjunctivitis|Neonatal conjunctivitis
C0027611|T047|PT|771.6|ICD9CM|Neonatal conjunctivitis and dacryocystitis|Neonatal conjunctivitis and dacryocystitis
C0276682|T047|AB|771.7|ICD9CM|Neonatal candida infect|Neonatal candida infect
C0276682|T047|PT|771.7|ICD9CM|Neonatal Candida infection|Neonatal Candida infection
C0158950|T046|HT|771.8|ICD9CM|Other infection specific to the perinatal period|Other infection specific to the perinatal period
C1135251|T047|AB|771.81|ICD9CM|NB septicemia [sepsis]|NB septicemia [sepsis]
C1135251|T047|PT|771.81|ICD9CM|Septicemia [sepsis] of newborn|Septicemia [sepsis] of newborn
C0235815|T047|AB|771.82|ICD9CM|NB urinary tract infectn|NB urinary tract infectn
C0235815|T047|PT|771.82|ICD9CM|Urinary tract infection of newborn|Urinary tract infection of newborn
C1135253|T047|AB|771.83|ICD9CM|Bacteremia of newborn|Bacteremia of newborn
C1135253|T047|PT|771.83|ICD9CM|Bacteremia of newborn|Bacteremia of newborn
C0158950|T046|PT|771.89|ICD9CM|Other infections specific to the perinatal period|Other infections specific to the perinatal period
C0158950|T046|AB|771.89|ICD9CM|Perinatal infection NEC|Perinatal infection NEC
C0473800|T046|HT|772|ICD9CM|Fetal and neonatal hemorrhage|Fetal and neonatal hemorrhage
C0158951|T046|PT|772.0|ICD9CM|Fetal blood loss|Fetal blood loss
C0158951|T046|AB|772.0|ICD9CM|NB fetal blood loss NEC|NB fetal blood loss NEC
C0270191|T046|HT|772.1|ICD9CM|Intraventricular hemorrhage of fetus or newborn|Intraventricular hemorrhage of fetus or newborn
C0949141|T047|PT|772.10|ICD9CM|Intraventricular hemorrhage unspecified grade|Intraventricular hemorrhage unspecified grade
C0949141|T047|AB|772.10|ICD9CM|NB intraven hem NOS|NB intraven hem NOS
C0949142|T047|PT|772.11|ICD9CM|Intraventricular hemorrhage, grade I|Intraventricular hemorrhage, grade I
C0949142|T047|AB|772.11|ICD9CM|NB intraven hem,grade i|NB intraven hem,grade i
C0949143|T047|PT|772.12|ICD9CM|Intraventricular hemorrhage, grade II|Intraventricular hemorrhage, grade II
C0949143|T047|AB|772.12|ICD9CM|NB intraven hem,grade ii|NB intraven hem,grade ii
C0949144|T047|PT|772.13|ICD9CM|Intraventricular hemorrhage, grade III|Intraventricular hemorrhage, grade III
C0949144|T047|AB|772.13|ICD9CM|NB intravn hem,grade iii|NB intravn hem,grade iii
C0949145|T047|PT|772.14|ICD9CM|Intraventricular hemorrhage, grade IV|Intraventricular hemorrhage, grade IV
C0949145|T047|AB|772.14|ICD9CM|NB intraven hem,grade iv|NB intraven hem,grade iv
C0854172|T046|AB|772.2|ICD9CM|NB subarachnoid hemorr|NB subarachnoid hemorr
C0854172|T046|PT|772.2|ICD9CM|Subarachnoid hemorrhage of fetus or newborn|Subarachnoid hemorrhage of fetus or newborn
C0473789|T046|AB|772.3|ICD9CM|Post-birth umbil hemorr|Post-birth umbil hemorr
C0473789|T046|PT|772.3|ICD9CM|Umbilical hemorrhage after birth|Umbilical hemorrhage after birth
C0158956|T047|PT|772.4|ICD9CM|Gastrointestinal hemorrhage of fetus or newborn|Gastrointestinal hemorrhage of fetus or newborn
C0158956|T047|AB|772.4|ICD9CM|NB GI hemorrhage|NB GI hemorrhage
C0158957|T046|PT|772.5|ICD9CM|Adrenal hemorrhage of fetus or newborn|Adrenal hemorrhage of fetus or newborn
C0158957|T046|AB|772.5|ICD9CM|NB adrenal hemorrhage|NB adrenal hemorrhage
C1390180|T046|PT|772.6|ICD9CM|Cutaneous hemorrhage of fetus or newborn|Cutaneous hemorrhage of fetus or newborn
C1390180|T046|AB|772.6|ICD9CM|NB cutaneous hemorrhage|NB cutaneous hemorrhage
C0158959|T046|AB|772.8|ICD9CM|Neonatal hemorrhage NEC|Neonatal hemorrhage NEC
C0158959|T046|PT|772.8|ICD9CM|Other specified hemorrhage of fetus or newborn|Other specified hemorrhage of fetus or newborn
C0270183|T046|AB|772.9|ICD9CM|Neonatal hemorrhage NOS|Neonatal hemorrhage NOS
C0270183|T046|PT|772.9|ICD9CM|Unspecified hemorrhage of newborn|Unspecified hemorrhage of newborn
C0014761|T047|HT|773|ICD9CM|Hemolytic disease of fetus or newborn, due to isoimmunization|Hemolytic disease of fetus or newborn, due to isoimmunization
C0158962|T047|PT|773.0|ICD9CM|Hemolytic disease of fetus or newborn due to Rh isoimmunization|Hemolytic disease of fetus or newborn due to Rh isoimmunization
C0158962|T047|AB|773.0|ICD9CM|NB hemolyt dis:rh isoimm|NB hemolyt dis:rh isoimm
C0270202|T047|PT|773.1|ICD9CM|Hemolytic disease of fetus or newborn due to ABO isoimmunization|Hemolytic disease of fetus or newborn due to ABO isoimmunization
C0270202|T047|AB|773.1|ICD9CM|NB hemolyt dis-abo isoim|NB hemolyt dis-abo isoim
C0014761|T047|PT|773.2|ICD9CM|Hemolytic disease of fetus or newborn due to other and unspecified isoimmunization|Hemolytic disease of fetus or newborn due to other and unspecified isoimmunization
C0014761|T047|AB|773.2|ICD9CM|NB hemolyt dis-isoim NEC|NB hemolyt dis-isoim NEC
C0455990|T047|PT|773.3|ICD9CM|Hydrops fetalis due to isoimmunization|Hydrops fetalis due to isoimmunization
C0455990|T047|AB|773.3|ICD9CM|Hydrops fetalis:isoimm|Hydrops fetalis:isoimm
C0270204|T047|PT|773.4|ICD9CM|Kernicterus of fetus or newborn due to isoimmunization|Kernicterus of fetus or newborn due to isoimmunization
C0270204|T047|AB|773.4|ICD9CM|NB kernicterus:isoimmun|NB kernicterus:isoimmun
C0158967|T047|PT|773.5|ICD9CM|Late anemia of fetus or newborn due to isoimmunization|Late anemia of fetus or newborn due to isoimmunization
C0158967|T047|AB|773.5|ICD9CM|NB late anemia:isoimmun|NB late anemia:isoimmun
C0158968|T046|HT|774|ICD9CM|Other perinatal jaundice|Other perinatal jaundice
C0158969|T047|AB|774.0|ICD9CM|Perinat jaund-hered anem|Perinat jaund-hered anem
C0158969|T047|PT|774.0|ICD9CM|Perinatal jaundice from hereditary hemolytic anemias|Perinatal jaundice from hereditary hemolytic anemias
C0701144|T047|AB|774.1|ICD9CM|Perinat jaund:hemolysis|Perinat jaund:hemolysis
C0701144|T047|PT|774.1|ICD9CM|Perinatal jaundice from other excessive hemolysis|Perinatal jaundice from other excessive hemolysis
C0158971|T046|AB|774.2|ICD9CM|Neonat jaund preterm del|Neonat jaund preterm del
C0158971|T046|PT|774.2|ICD9CM|Neonatal jaundice associated with preterm delivery|Neonatal jaundice associated with preterm delivery
C0158972|T047|HT|774.3|ICD9CM|Neonatal jaundice due to delayed conjugation from other causes|Neonatal jaundice due to delayed conjugation from other causes
C0375543|T046|AB|774.30|ICD9CM|Delay conjugat jaund NOS|Delay conjugat jaund NOS
C0375543|T046|PT|774.30|ICD9CM|Neonatal jaundice due to delayed conjugation, cause unspecified|Neonatal jaundice due to delayed conjugation, cause unspecified
C0158974|T047|AB|774.31|ICD9CM|Neonat jaund in oth dis|Neonat jaund in oth dis
C0158974|T047|PT|774.31|ICD9CM|Neonatal jaundice due to delayed conjugation in diseases classified elsewhere|Neonatal jaundice due to delayed conjugation in diseases classified elsewhere
C0158975|T046|AB|774.39|ICD9CM|Delay conjugat jaund NEC|Delay conjugat jaund NEC
C0158975|T046|PT|774.39|ICD9CM|Other neonatal jaundice due to delayed conjugation from other causes|Other neonatal jaundice due to delayed conjugation from other causes
C0158976|T047|AB|774.4|ICD9CM|Fetal/neonatal hepatitis|Fetal/neonatal hepatitis
C0158976|T047|PT|774.4|ICD9CM|Perinatal jaundice due to hepatocellular damage|Perinatal jaundice due to hepatocellular damage
C0158977|T047|PT|774.5|ICD9CM|Perinatal jaundice from other causes|Perinatal jaundice from other causes
C0158977|T047|AB|774.5|ICD9CM|Perinatal jaundice NEC|Perinatal jaundice NEC
C0270206|T047|AB|774.6|ICD9CM|Fetal/neonatal jaund NOS|Fetal/neonatal jaund NOS
C0270206|T047|PT|774.6|ICD9CM|Unspecified fetal and neonatal jaundice|Unspecified fetal and neonatal jaundice
C0158978|T047|PT|774.7|ICD9CM|Kernicterus of fetus or newborn not due to isoimmunization|Kernicterus of fetus or newborn not due to isoimmunization
C0158978|T047|AB|774.7|ICD9CM|NB kernicterus|NB kernicterus
C0158979|T047|HT|775|ICD9CM|Endocrine and metabolic disturbances specific to the fetus and newborn|Endocrine and metabolic disturbances specific to the fetus and newborn
C0270221|T047|AB|775.0|ICD9CM|Infant diabet mother syn|Infant diabet mother syn
C0270221|T047|PT|775.0|ICD9CM|Syndrome of "infant of a diabetic mother"|Syndrome of "infant of a diabetic mother"
C0158981|T047|AB|775.1|ICD9CM|Neonat diabetes mellitus|Neonat diabetes mellitus
C0158981|T047|PT|775.1|ICD9CM|Neonatal diabetes mellitus|Neonatal diabetes mellitus
C0158982|T047|AB|775.2|ICD9CM|Neonat myasthenia gravis|Neonat myasthenia gravis
C0158982|T047|PT|775.2|ICD9CM|Neonatal myasthenia gravis|Neonatal myasthenia gravis
C0158983|T047|AB|775.3|ICD9CM|Neonatal thyrotoxicosis|Neonatal thyrotoxicosis
C0158983|T047|PT|775.3|ICD9CM|Neonatal thyrotoxicosis|Neonatal thyrotoxicosis
C0158984|T047|AB|775.4|ICD9CM|Hypocalcem/hypomagnes NB|Hypocalcem/hypomagnes NB
C0158984|T047|PT|775.4|ICD9CM|Hypocalcemia and hypomagnesemia of newborn|Hypocalcemia and hypomagnesemia of newborn
C0495447|T047|AB|775.5|ICD9CM|Neonatal dehydration|Neonatal dehydration
C0495447|T047|PT|775.5|ICD9CM|Other transitory neonatal electrolyte disturbances|Other transitory neonatal electrolyte disturbances
C0158986|T047|AB|775.6|ICD9CM|Neonatal hypoglycemia|Neonatal hypoglycemia
C0158986|T047|PT|775.6|ICD9CM|Neonatal hypoglycemia|Neonatal hypoglycemia
C0158987|T033|AB|775.7|ICD9CM|Late metab acidosis NB|Late metab acidosis NB
C0158987|T033|PT|775.7|ICD9CM|Late metabolic acidosis of newborn|Late metabolic acidosis of newborn
C1719633|T047|HT|775.8|ICD9CM|Other neonatal endocrine and metabolic disturbances|Other neonatal endocrine and metabolic disturbances
C1719629|T047|AB|775.81|ICD9CM|NB acidosis NEC|NB acidosis NEC
C1719629|T047|PT|775.81|ICD9CM|Other acidosis of newborn|Other acidosis of newborn
C1719633|T047|AB|775.89|ICD9CM|Neonat endo/met dis NEC|Neonat endo/met dis NEC
C1719633|T047|PT|775.89|ICD9CM|Other neonatal endocrine and metabolic disturbances|Other neonatal endocrine and metabolic disturbances
C0158989|T047|AB|775.9|ICD9CM|Transient met dis NB NOS|Transient met dis NB NOS
C0158989|T047|PT|775.9|ICD9CM|Unspecified endocrine and metabolic disturbances specific to the fetus and newborn|Unspecified endocrine and metabolic disturbances specific to the fetus and newborn
C1285368|T047|HT|776|ICD9CM|Hematological disorders of newborn|Hematological disorders of newborn
C0019088|T047|PT|776.0|ICD9CM|Hemorrhagic disease of newborn|Hemorrhagic disease of newborn
C0019088|T047|AB|776.0|ICD9CM|NB hemorrhagic disease|NB hemorrhagic disease
C0158991|T047|AB|776.1|ICD9CM|Neonatal thrombocytopen|Neonatal thrombocytopen
C0158991|T047|PT|776.1|ICD9CM|Transient neonatal thrombocytopenia|Transient neonatal thrombocytopenia
C0158992|T047|AB|776.2|ICD9CM|Dissem intravasc coag NB|Dissem intravasc coag NB
C0158992|T047|PT|776.2|ICD9CM|Disseminated intravascular coagulation in newborn|Disseminated intravascular coagulation in newborn
C0158993|T047|AB|776.3|ICD9CM|Oth neonatal coag dis|Oth neonatal coag dis
C0158993|T047|PT|776.3|ICD9CM|Other transient neonatal disorders of coagulation|Other transient neonatal disorders of coagulation
C0272153|T047|AB|776.4|ICD9CM|Polycythemia neonatorum|Polycythemia neonatorum
C0272153|T047|PT|776.4|ICD9CM|Polycythemia neonatorum|Polycythemia neonatorum
C0158995|T047|AB|776.5|ICD9CM|Congenital anemia|Congenital anemia
C0158995|T047|PT|776.5|ICD9CM|Congenital anemia|Congenital anemia
C0158996|T047|AB|776.6|ICD9CM|Anemia of prematurity|Anemia of prematurity
C0158996|T047|PT|776.6|ICD9CM|Anemia of prematurity|Anemia of prematurity
C0158997|T047|AB|776.7|ICD9CM|Neonatal neutropenia|Neonatal neutropenia
C0158997|T047|PT|776.7|ICD9CM|Transient neonatal neutropenia|Transient neonatal neutropenia
C0158998|T047|PT|776.8|ICD9CM|Other specified transient hematological disorders of fetus or newborn|Other specified transient hematological disorders of fetus or newborn
C0158998|T047|AB|776.8|ICD9CM|Transient hemat dis NEC|Transient hemat dis NEC
C0158999|T047|AB|776.9|ICD9CM|NB hematological dis NOS|NB hematological dis NOS
C0158999|T047|PT|776.9|ICD9CM|Unspecified hematological disorder specific to newborn|Unspecified hematological disorder specific to newborn
C0159000|T047|HT|777|ICD9CM|Perinatal disorders of digestive system|Perinatal disorders of digestive system
C0270246|T047|AB|777.1|ICD9CM|Meconium obstruction|Meconium obstruction
C0270246|T047|PT|777.1|ICD9CM|Meconium obstruction in fetus or newborn|Meconium obstruction in fetus or newborn
C0400853|T047|AB|777.2|ICD9CM|Intest obst-inspiss milk|Intest obst-inspiss milk
C0400853|T047|PT|777.2|ICD9CM|Intestinal obstruction in newborn due to inspissated milk|Intestinal obstruction in newborn due to inspissated milk
C0270249|T046|PT|777.3|ICD9CM|Hematemesis and melena of newborn due to swallowed maternal blood|Hematemesis and melena of newborn due to swallowed maternal blood
C0270249|T046|AB|777.3|ICD9CM|Swallowed blood syndrome|Swallowed blood syndrome
C0159004|T020|AB|777.4|ICD9CM|Transitory ileus of NB|Transitory ileus of NB
C0159004|T020|PT|777.4|ICD9CM|Transitory ileus of newborn|Transitory ileus of newborn
C2349669|T047|HT|777.5|ICD9CM|Necrotizing enterocolitis in newborn|Necrotizing enterocolitis in newborn
C2349662|T047|AB|777.50|ICD9CM|Nec enterocoltis NB NOS|Nec enterocoltis NB NOS
C2349662|T047|PT|777.50|ICD9CM|Necrotizing enterocolitis in newborn, unspecified|Necrotizing enterocolitis in newborn, unspecified
C2910076|T047|PT|777.51|ICD9CM|Stage I necrotizing enterocolitis in newborn|Stage I necrotizing enterocolitis in newborn
C2910076|T047|AB|777.51|ICD9CM|Stg I nec enterocol NB|Stg I nec enterocol NB
C2910077|T047|PT|777.52|ICD9CM|Stage II necrotizing enterocolitis in newborn|Stage II necrotizing enterocolitis in newborn
C2910077|T047|AB|777.52|ICD9CM|Stg II nec enterocol NB|Stg II nec enterocol NB
C2910078|T047|PT|777.53|ICD9CM|Stage III necrotizing enterocolitis in newborn|Stage III necrotizing enterocolitis in newborn
C2910078|T047|AB|777.53|ICD9CM|Stg III nec enterocol NB|Stg III nec enterocol NB
C0159006|T047|AB|777.6|ICD9CM|Perinatal intest perfor|Perinatal intest perfor
C0159006|T047|PT|777.6|ICD9CM|Perinatal intestinal perforation|Perinatal intestinal perforation
C0159007|T047|PT|777.8|ICD9CM|Other specified perinatal disorders of digestive system|Other specified perinatal disorders of digestive system
C0159007|T047|AB|777.8|ICD9CM|Perinat GI sys dis NEC|Perinat GI sys dis NEC
C0159000|T047|AB|777.9|ICD9CM|Perinat GI sys dis NOS|Perinat GI sys dis NOS
C0159000|T047|PT|777.9|ICD9CM|Unspecified perinatal disorder of digestive system|Unspecified perinatal disorder of digestive system
C0159009|T046|HT|778|ICD9CM|Conditions involving the integument and temperature regulation of fetus and newborn|Conditions involving the integument and temperature regulation of fetus and newborn
C0455988|T047|AB|778.0|ICD9CM|Hydrops fetalis no isoim|Hydrops fetalis no isoim
C0455988|T047|PT|778.0|ICD9CM|Hydrops fetalis not due to isoimmunization|Hydrops fetalis not due to isoimmunization
C0036415|T019|AB|778.1|ICD9CM|Sclerema neonatorum|Sclerema neonatorum
C0036415|T019|PT|778.1|ICD9CM|Sclerema neonatorum|Sclerema neonatorum
C0159011|T047|PT|778.2|ICD9CM|Cold injury syndrome of newborn|Cold injury syndrome of newborn
C0159011|T047|AB|778.2|ICD9CM|NB cold injury syndrome|NB cold injury syndrome
C0159012|T046|AB|778.3|ICD9CM|NB hypothermia NEC|NB hypothermia NEC
C0159012|T046|PT|778.3|ICD9CM|Other hypothermia of newborn|Other hypothermia of newborn
C0159013|T047|AB|778.4|ICD9CM|NB temp regulat dis NEC|NB temp regulat dis NEC
C0159013|T047|PT|778.4|ICD9CM|Other disturbances of temperature regulation of newborn|Other disturbances of temperature regulation of newborn
C0159014|T046|AB|778.5|ICD9CM|Edema of newborn NEC/NOS|Edema of newborn NEC/NOS
C0159014|T046|PT|778.5|ICD9CM|Other and unspecified edema of newborn|Other and unspecified edema of newborn
C0159015|T019|AB|778.6|ICD9CM|Congenital hydrocele|Congenital hydrocele
C0159015|T019|PT|778.6|ICD9CM|Congenital hydrocele|Congenital hydrocele
C1449721|T047|PT|778.7|ICD9CM|Breast engorgement in newborn|Breast engorgement in newborn
C1449721|T047|AB|778.7|ICD9CM|NB breast engorgement|NB breast engorgement
C0477961|T047|AB|778.8|ICD9CM|NB integument cond NEC|NB integument cond NEC
C0477961|T047|PT|778.8|ICD9CM|Other specified conditions involving the integument of fetus and newborn|Other specified conditions involving the integument of fetus and newborn
C0159018|T047|AB|778.9|ICD9CM|NB integument cond NOS|NB integument cond NOS
C0159018|T047|PT|778.9|ICD9CM|Unspecified condition involving the integument and temperature regulation of fetus and newborn|Unspecified condition involving the integument and temperature regulation of fetus and newborn
C0159019|T047|HT|779|ICD9CM|Other and ill-defined conditions originating in the perinatal period|Other and ill-defined conditions originating in the perinatal period
C0159020|T047|AB|779.0|ICD9CM|Convulsions in newborn|Convulsions in newborn
C0159020|T047|PT|779.0|ICD9CM|Convulsions in newborn|Convulsions in newborn
C0159021|T047|AB|779.1|ICD9CM|NB cereb irrit NEC/NOS|NB cereb irrit NEC/NOS
C0159021|T047|PT|779.1|ICD9CM|Other and unspecified cerebral irritability in newborn|Other and unspecified cerebral irritability in newborn
C0159022|T047|PT|779.2|ICD9CM|Cerebral depression, coma, and other abnormal cerebral signs in fetus or newborn|Cerebral depression, coma, and other abnormal cerebral signs in fetus or newborn
C0159022|T047|AB|779.2|ICD9CM|Cns dysfunction syn NB|Cns dysfunction syn NB
C2712941|T047|HT|779.3|ICD9CM|Disorder of stomach function and feeding problems in newborn|Disorder of stomach function and feeding problems in newborn
C0159023|T033|PT|779.31|ICD9CM|Feeding problems in newborn|Feeding problems in newborn
C0159023|T033|AB|779.31|ICD9CM|NB feeding problems|NB feeding problems
C2712362|T184|PT|779.32|ICD9CM|Bilious vomiting in newborn|Bilious vomiting in newborn
C2712362|T184|AB|779.32|ICD9CM|NB bilious vomiting|NB bilious vomiting
C2712363|T047|AB|779.33|ICD9CM|NB other vomiting|NB other vomiting
C2712363|T047|PT|779.33|ICD9CM|Other vomiting in newborn|Other vomiting in newborn
C2712364|T047|PT|779.34|ICD9CM|Failure to thrive in newborn|Failure to thrive in newborn
C2712364|T047|AB|779.34|ICD9CM|NB failure to thrive|NB failure to thrive
C0270275|T037|PT|779.4|ICD9CM|Drug reactions and intoxications specific to newborn|Drug reactions and intoxications specific to newborn
C0270275|T037|AB|779.4|ICD9CM|NB drug reaction/intoxic|NB drug reaction/intoxic
C0027609|T047|PT|779.5|ICD9CM|Drug withdrawal syndrome in newborn|Drug withdrawal syndrome in newborn
C0027609|T047|AB|779.5|ICD9CM|NB drug withdrawal syndr|NB drug withdrawal syndr
C1704300|T033|AB|779.6|ICD9CM|Termination of pregnancy|Termination of pregnancy
C1704300|T033|PT|779.6|ICD9CM|Termination of pregnancy (fetus)|Termination of pregnancy (fetus)
C0023529|T047|AB|779.7|ICD9CM|Perivent leukomalacia|Perivent leukomalacia
C0023529|T047|PT|779.7|ICD9CM|Periventricular leukomalacia|Periventricular leukomalacia
C0159027|T047|HT|779.8|ICD9CM|Other specified conditions originating in the perinatal period|Other specified conditions originating in the perinatal period
C1112488|T046|AB|779.81|ICD9CM|Neonatal bradycardia|Neonatal bradycardia
C1112488|T046|PT|779.81|ICD9CM|Neonatal bradycardia|Neonatal bradycardia
C0877308|T046|AB|779.82|ICD9CM|Neonatal tachycardia|Neonatal tachycardia
C0877308|T046|PT|779.82|ICD9CM|Neonatal tachycardia|Neonatal tachycardia
C1260438|T046|AB|779.83|ICD9CM|Delay separate umbl cord|Delay separate umbl cord
C1260438|T046|PT|779.83|ICD9CM|Delayed separation of umbilical cord|Delayed separation of umbilical cord
C1112318|T046|AB|779.84|ICD9CM|Meconium staining|Meconium staining
C1112318|T046|PT|779.84|ICD9CM|Meconium staining|Meconium staining
C1410098|T046|PT|779.85|ICD9CM|Cardiac arrest of newborn|Cardiac arrest of newborn
C1410098|T046|AB|779.85|ICD9CM|NB cardiac arrest|NB cardiac arrest
C0159027|T047|PT|779.89|ICD9CM|Other specified conditions originating in the perinatal period|Other specified conditions originating in the perinatal period
C0159027|T047|AB|779.89|ICD9CM|Perinatal condition NEC|Perinatal condition NEC
C0270075|T047|AB|779.9|ICD9CM|Perinatal condition NOS|Perinatal condition NOS
C0270075|T047|PT|779.9|ICD9CM|Unspecified condition originating in the perinatal period|Unspecified condition originating in the perinatal period
C0159028|T184|HT|780|ICD9CM|General symptoms|General symptoms
C1457887|T184|HT|780-789.99|ICD9CM|SYMPTOMS|SYMPTOMS
C0178310|T184|HT|780-799.99|ICD9CM|SYMPTOMS, SIGNS, AND ILL-DEFINED CONDITIONS|SYMPTOMS, SIGNS, AND ILL-DEFINED CONDITIONS
C0234428|T033|HT|780.0|ICD9CM|Alteration of consciousness|Alteration of consciousness
C0009421|T047|AB|780.01|ICD9CM|Coma|Coma
C0009421|T047|PT|780.01|ICD9CM|Coma|Coma
C0221539|T184|AB|780.02|ICD9CM|Trans alter awareness|Trans alter awareness
C0221539|T184|PT|780.02|ICD9CM|Transient alteration of awareness|Transient alteration of awareness
C0242670|T047|PT|780.03|ICD9CM|Persistent vegetative state|Persistent vegetative state
C0242670|T047|AB|780.03|ICD9CM|Persistent vegtv state|Persistent vegtv state
C0221540|T184|AB|780.09|ICD9CM|Other alter consciousnes|Other alter consciousnes
C0221540|T184|PT|780.09|ICD9CM|Other alteration of consciousness|Other alteration of consciousness
C0018524|T048|AB|780.1|ICD9CM|Hallucinations|Hallucinations
C0018524|T048|PT|780.1|ICD9CM|Hallucinations|Hallucinations
C0039070|T184|AB|780.2|ICD9CM|Syncope and collapse|Syncope and collapse
C0039070|T184|PT|780.2|ICD9CM|Syncope and collapse|Syncope and collapse
C4048158|T184|HT|780.3|ICD9CM|Convulsions|Convulsions
C0009952|T047|PT|780.31|ICD9CM|Febrile convulsions (simple), unspecified|Febrile convulsions (simple), unspecified
C0009952|T047|AB|780.31|ICD9CM|Febrile convulsions NOS|Febrile convulsions NOS
C0751057|T047|PT|780.32|ICD9CM|Complex febrile convulsions|Complex febrile convulsions
C0751057|T047|AB|780.32|ICD9CM|Complx febrile convulsns|Complx febrile convulsns
C2921125|T047|PT|780.33|ICD9CM|Post traumatic seizures|Post traumatic seizures
C2921125|T047|AB|780.33|ICD9CM|Post traumatic seizures|Post traumatic seizures
C0490011|T184|AB|780.39|ICD9CM|Convulsions NEC|Convulsions NEC
C0490011|T184|PT|780.39|ICD9CM|Other convulsions|Other convulsions
C0476206|T184|AB|780.4|ICD9CM|Dizziness and giddiness|Dizziness and giddiness
C0476206|T184|PT|780.4|ICD9CM|Dizziness and giddiness|Dizziness and giddiness
C0037317|T184|HT|780.5|ICD9CM|Sleep disturbances|Sleep disturbances
C0037317|T184|AB|780.50|ICD9CM|Sleep disturbance NOS|Sleep disturbance NOS
C0037317|T184|PT|780.50|ICD9CM|Sleep disturbance, unspecified|Sleep disturbance, unspecified
C1561813|T184|AB|780.51|ICD9CM|Insomn w sleep apnea NOS|Insomn w sleep apnea NOS
C1561813|T184|PT|780.51|ICD9CM|Insomnia with sleep apnea, unspecified|Insomnia with sleep apnea, unspecified
C0917801|T184|AB|780.52|ICD9CM|Insomnia NOS|Insomnia NOS
C0917801|T184|PT|780.52|ICD9CM|Insomnia, unspecified|Insomnia, unspecified
C1561815|T184|AB|780.53|ICD9CM|Hypersom w slp apnea NOS|Hypersom w slp apnea NOS
C1561815|T184|PT|780.53|ICD9CM|Hypersomnia with sleep apnea, unspecified|Hypersomnia with sleep apnea, unspecified
C0917799|T047|AB|780.54|ICD9CM|Hypersomnia NOS|Hypersomnia NOS
C0917799|T047|PT|780.54|ICD9CM|Hypersomnia, unspecified|Hypersomnia, unspecified
C1561817|T184|PT|780.55|ICD9CM|Disruption of 24 hour sleep wake cycle, unspecified|Disruption of 24 hour sleep wake cycle, unspecified
C1561817|T184|AB|780.55|ICD9CM|Irreg sleep-wake rhy NOS|Irreg sleep-wake rhy NOS
C0013373|T048|PT|780.56|ICD9CM|Dysfunctions associated with sleep stages or arousal from sleep|Dysfunctions associated with sleep stages or arousal from sleep
C0013373|T048|AB|780.56|ICD9CM|Sleep stage dysfunctions|Sleep stage dysfunctions
C0037315|T047|AB|780.57|ICD9CM|Sleep apnea NOS|Sleep apnea NOS
C0037315|T047|PT|780.57|ICD9CM|Unspecified sleep apnea|Unspecified sleep apnea
C1561818|T047|AB|780.58|ICD9CM|Sleep rel move disor NOS|Sleep rel move disor NOS
C1561818|T047|PT|780.58|ICD9CM|Sleep related movement disorder, unspecified|Sleep related movement disorder, unspecified
C1962929|T047|PT|780.59|ICD9CM|Other sleep disturbances|Other sleep disturbances
C1962929|T047|AB|780.59|ICD9CM|Sleep disturbances NEC|Sleep disturbances NEC
C2349675|T184|HT|780.6|ICD9CM|Fever and other physiologic disturbances of temperature regulation|Fever and other physiologic disturbances of temperature regulation
C0015967|T184|AB|780.60|ICD9CM|Fever NOS|Fever NOS
C0015967|T184|PT|780.60|ICD9CM|Fever, unspecified|Fever, unspecified
C2349670|T047|AB|780.61|ICD9CM|Fever in other diseases|Fever in other diseases
C2349670|T047|PT|780.61|ICD9CM|Fever presenting with conditions classified elsewhere|Fever presenting with conditions classified elsewhere
C2349671|T046|PT|780.62|ICD9CM|Postprocedural fever|Postprocedural fever
C2349671|T046|AB|780.62|ICD9CM|Postprocedural fever|Postprocedural fever
C2349672|T046|PT|780.63|ICD9CM|Postvaccination fever|Postvaccination fever
C2349672|T046|AB|780.63|ICD9CM|Postvaccination fever|Postvaccination fever
C2349674|T184|PT|780.64|ICD9CM|Chills (without fever)|Chills (without fever)
C2349674|T184|AB|780.64|ICD9CM|Chills (without fever)|Chills (without fever)
C3542020|T033|PT|780.65|ICD9CM|Hypothermia not associated with low environmental temperature|Hypothermia not associated with low environmental temperature
C3542020|T033|AB|780.65|ICD9CM|Hypothrm-wo low env tmp|Hypothrm-wo low env tmp
C1739123|T046|AB|780.66|ICD9CM|Feb nonhemo transf react|Feb nonhemo transf react
C1739123|T046|PT|780.66|ICD9CM|Febrile nonhemolytic transfusion reaction|Febrile nonhemolytic transfusion reaction
C0024528|T184|HT|780.7|ICD9CM|Malaise and fatigue|Malaise and fatigue
C0015674|T047|AB|780.71|ICD9CM|Chronic fatigue syndrome|Chronic fatigue syndrome
C0015674|T047|PT|780.71|ICD9CM|Chronic fatigue syndrome|Chronic fatigue syndrome
C3543852|T047|PT|780.72|ICD9CM|Functional quadriplegia|Functional quadriplegia
C3543852|T047|AB|780.72|ICD9CM|Functional quadriplegia|Functional quadriplegia
C0695252|T184|AB|780.79|ICD9CM|Malaise and fatigue NEC|Malaise and fatigue NEC
C0695252|T184|PT|780.79|ICD9CM|Other malaise and fatigue|Other malaise and fatigue
C0476476|T033|AB|780.8|ICD9CM|Generalizd hyperhidrosis|Generalizd hyperhidrosis
C0476476|T033|PT|780.8|ICD9CM|Generalized hyperhidrosis|Generalized hyperhidrosis
C0029625|T184|HT|780.9|ICD9CM|Other general symptoms|Other general symptoms
C1135254|T047|PT|780.91|ICD9CM|Fussy infant (baby)|Fussy infant (baby)
C1135254|T047|AB|780.91|ICD9CM|Fussy infant/baby|Fussy infant/baby
C0497134|T033|AB|780.92|ICD9CM|Excess cry infant/baby|Excess cry infant/baby
C0497134|T033|PT|780.92|ICD9CM|Excessive crying of infant (baby)|Excessive crying of infant (baby)
C0751295|T184|AB|780.93|ICD9CM|Memory loss|Memory loss
C0751295|T184|PT|780.93|ICD9CM|Memory loss|Memory loss
C0239233|T184|AB|780.94|ICD9CM|Early satiety|Early satiety
C0239233|T184|PT|780.94|ICD9CM|Early satiety|Early satiety
C1719639|T033|PT|780.95|ICD9CM|Excessive crying of child, adolescent, or adult|Excessive crying of child, adolescent, or adult
C1719639|T033|AB|780.95|ICD9CM|Excs cry chld,adol,adult|Excs cry chld,adol,adult
C0281856|T184|PT|780.96|ICD9CM|Generalized pain|Generalized pain
C0281856|T184|AB|780.96|ICD9CM|Generalized pain|Generalized pain
C0278061|T048|PT|780.97|ICD9CM|Altered mental status|Altered mental status
C0278061|T048|AB|780.97|ICD9CM|Altered mental status|Altered mental status
C0029625|T184|AB|780.99|ICD9CM|Other general symptoms|Other general symptoms
C0029625|T184|PT|780.99|ICD9CM|Other general symptoms|Other general symptoms
C0159033|T184|HT|781|ICD9CM|Symptoms involving nervous and musculoskeletal systems|Symptoms involving nervous and musculoskeletal systems
C0392702|T047|AB|781.0|ICD9CM|Abn involun movement NEC|Abn involun movement NEC
C0392702|T047|PT|781.0|ICD9CM|Abnormal involuntary movements|Abnormal involuntary movements
C0495689|T033|PT|781.1|ICD9CM|Disturbances of sensation of smell and taste|Disturbances of sensation of smell and taste
C0495689|T033|AB|781.1|ICD9CM|Smell & taste disturb|Smell & taste disturb
C0575081|T033|AB|781.2|ICD9CM|Abnormality of gait|Abnormality of gait
C0575081|T033|PT|781.2|ICD9CM|Abnormality of gait|Abnormality of gait
C0520966|T033|AB|781.3|ICD9CM|Lack of coordination|Lack of coordination
C0520966|T033|PT|781.3|ICD9CM|Lack of coordination|Lack of coordination
C0159034|T184|AB|781.4|ICD9CM|Transient limb paralysis|Transient limb paralysis
C0159034|T184|PT|781.4|ICD9CM|Transient paralysis of limb|Transient paralysis of limb
C0009080|T190|AB|781.5|ICD9CM|Clubbing of fingers|Clubbing of fingers
C0009080|T190|PT|781.5|ICD9CM|Clubbing of fingers|Clubbing of fingers
C0025287|T184|AB|781.6|ICD9CM|Meningismus|Meningismus
C0025287|T184|PT|781.6|ICD9CM|Meningismus|Meningismus
C0039621|T033|AB|781.7|ICD9CM|Tetany|Tetany
C0039621|T033|PT|781.7|ICD9CM|Tetany|Tetany
C0840927|T047|AB|781.8|ICD9CM|Neurologic neglect syndr|Neurologic neglect syndr
C0840927|T047|PT|781.8|ICD9CM|Neurologic neglect syndrome|Neurologic neglect syndrome
C0159036|T184|HT|781.9|ICD9CM|Other symptoms involving nervous and musculoskeletal systems|Other symptoms involving nervous and musculoskeletal systems
C0424641|T033|AB|781.91|ICD9CM|Loss of height|Loss of height
C0424641|T033|PT|781.91|ICD9CM|Loss of height|Loss of height
C0231471|T033|AB|781.92|ICD9CM|Abnormal posture|Abnormal posture
C0231471|T033|PT|781.92|ICD9CM|Abnormal posture|Abnormal posture
C0028856|T047|AB|781.93|ICD9CM|Ocular torticollis|Ocular torticollis
C0028856|T047|PT|781.93|ICD9CM|Ocular torticollis|Ocular torticollis
C0427055|T047|AB|781.94|ICD9CM|Facial weakness|Facial weakness
C0427055|T047|PT|781.94|ICD9CM|Facial weakness|Facial weakness
C0159036|T184|AB|781.99|ICD9CM|Nerve/musculskel sym NEC|Nerve/musculskel sym NEC
C0159036|T184|PT|781.99|ICD9CM|Other symptoms involving nervous and musculoskeletal systems|Other symptoms involving nervous and musculoskeletal systems
C0159037|T184|HT|782|ICD9CM|Symptoms involving skin and other integumentary tissue|Symptoms involving skin and other integumentary tissue
C0012766|T184|PT|782.0|ICD9CM|Disturbance of skin sensation|Disturbance of skin sensation
C0012766|T184|AB|782.0|ICD9CM|Skin sensation disturb|Skin sensation disturb
C0015230|T184|AB|782.1|ICD9CM|Nonspecif skin erupt NEC|Nonspecif skin erupt NEC
C0015230|T184|PT|782.1|ICD9CM|Rash and other nonspecific skin eruption|Rash and other nonspecific skin eruption
C0476228|T184|AB|782.2|ICD9CM|Local suprficial swellng|Local suprficial swellng
C0476228|T184|PT|782.2|ICD9CM|Localized superficial swelling, mass, or lump|Localized superficial swelling, mass, or lump
C0013604|T046|AB|782.3|ICD9CM|Edema|Edema
C0013604|T046|PT|782.3|ICD9CM|Edema|Edema
C0476232|T184|AB|782.4|ICD9CM|Jaundice NOS|Jaundice NOS
C0476232|T184|PT|782.4|ICD9CM|Jaundice, unspecified, not of newborn|Jaundice, unspecified, not of newborn
C0010520|T184|AB|782.5|ICD9CM|Cyanosis|Cyanosis
C0010520|T184|PT|782.5|ICD9CM|Cyanosis|Cyanosis
C0159038|T184|HT|782.6|ICD9CM|Pallor and flushing|Pallor and flushing
C0030232|T033|AB|782.61|ICD9CM|Pallor|Pallor
C0030232|T033|PT|782.61|ICD9CM|Pallor|Pallor
C0016382|T184|AB|782.62|ICD9CM|Flushing|Flushing
C0016382|T184|PT|782.62|ICD9CM|Flushing|Flushing
C0159039|T046|AB|782.7|ICD9CM|Spontaneous ecchymoses|Spontaneous ecchymoses
C0159039|T046|PT|782.7|ICD9CM|Spontaneous ecchymoses|Spontaneous ecchymoses
C0159040|T184|AB|782.8|ICD9CM|Changes in skin texture|Changes in skin texture
C0159040|T184|PT|782.8|ICD9CM|Changes in skin texture|Changes in skin texture
C0159037|T184|AB|782.9|ICD9CM|Integument tiss symp NEC|Integument tiss symp NEC
C0159037|T184|PT|782.9|ICD9CM|Other symptoms involving skin and integumentary tissues|Other symptoms involving skin and integumentary tissues
C0476235|T184|HT|783|ICD9CM|Symptoms concerning nutrition, metabolism, and development|Symptoms concerning nutrition, metabolism, and development
C0003123|T047|AB|783.0|ICD9CM|Anorexia|Anorexia
C0003123|T047|PT|783.0|ICD9CM|Anorexia|Anorexia
C0332544|T184|AB|783.1|ICD9CM|Abnormal weight gain|Abnormal weight gain
C0332544|T184|PT|783.1|ICD9CM|Abnormal weight gain|Abnormal weight gain
C0878752|T184|HT|783.2|ICD9CM|Abnormal loss of weight and underweight|Abnormal loss of weight and underweight
C1262477|T033|AB|783.21|ICD9CM|Abnormal loss of weight|Abnormal loss of weight
C1262477|T033|PT|783.21|ICD9CM|Loss of weight|Loss of weight
C0041667|T033|AB|783.22|ICD9CM|Underweight|Underweight
C0041667|T033|PT|783.22|ICD9CM|Underweight|Underweight
C0699815|T033|PT|783.3|ICD9CM|Feeding difficulties and mismanagement|Feeding difficulties and mismanagement
C0699815|T033|AB|783.3|ICD9CM|Feeding problem|Feeding problem
C0878753|T184|HT|783.4|ICD9CM|Lack of expected normal physiological development in childhood|Lack of expected normal physiological development in childhood
C0878706|T184|AB|783.40|ICD9CM|Lack norm physio dev NOS|Lack norm physio dev NOS
C0878706|T184|PT|783.40|ICD9CM|Lack of normal physiological development, unspecified|Lack of normal physiological development, unspecified
C0015544|T047|PT|783.41|ICD9CM|Failure to thrive|Failure to thrive
C0015544|T047|AB|783.41|ICD9CM|Failure to thrive-child|Failure to thrive-child
C0476241|T033|AB|783.42|ICD9CM|Delayed milestones|Delayed milestones
C0476241|T033|PT|783.42|ICD9CM|Delayed milestones|Delayed milestones
C0349588|T033|AB|783.43|ICD9CM|Short stature|Short stature
C0349588|T033|PT|783.43|ICD9CM|Short stature|Short stature
C0085602|T184|AB|783.5|ICD9CM|Polydipsia|Polydipsia
C0085602|T184|PT|783.5|ICD9CM|Polydipsia|Polydipsia
C0020505|T033|AB|783.6|ICD9CM|Polyphagia|Polyphagia
C0020505|T033|PT|783.6|ICD9CM|Polyphagia|Polyphagia
C1998978|T047|PT|783.7|ICD9CM|Adult failure to thrive|Adult failure to thrive
C1998978|T047|AB|783.7|ICD9CM|Failure to thrive-adult|Failure to thrive-adult
C0159043|T184|AB|783.9|ICD9CM|Nutr/metab/devel sym NEC|Nutr/metab/devel sym NEC
C0159043|T184|PT|783.9|ICD9CM|Other symptoms concerning nutrition, metabolism, and development|Other symptoms concerning nutrition, metabolism, and development
C0476247|T184|HT|784|ICD9CM|Symptoms involving head and neck|Symptoms involving head and neck
C0018681|T184|AB|784.0|ICD9CM|Headache|Headache
C0018681|T184|PT|784.0|ICD9CM|Headache|Headache
C0242429|T184|AB|784.1|ICD9CM|Throat pain|Throat pain
C0242429|T184|PT|784.1|ICD9CM|Throat pain|Throat pain
C0159045|T184|AB|784.2|ICD9CM|Swelling in head & neck|Swelling in head & neck
C0159045|T184|PT|784.2|ICD9CM|Swelling, mass, or lump in head and neck|Swelling, mass, or lump in head and neck
C0003537|T048|AB|784.3|ICD9CM|Aphasia|Aphasia
C0003537|T048|PT|784.3|ICD9CM|Aphasia|Aphasia
C2712707|T046|HT|784.4|ICD9CM|Voice and resonance disorders|Voice and resonance disorders
C2712365|T046|PT|784.40|ICD9CM|Voice and resonance disorder, unspecified|Voice and resonance disorder, unspecified
C2712365|T046|AB|784.40|ICD9CM|Voice/resonance dis NOS|Voice/resonance dis NOS
C0003564|T184|AB|784.41|ICD9CM|Aphonia|Aphonia
C0003564|T184|PT|784.41|ICD9CM|Aphonia|Aphonia
C1527344|T048|AB|784.42|ICD9CM|Dysphonia|Dysphonia
C1527344|T048|PT|784.42|ICD9CM|Dysphonia|Dysphonia
C0264614|T047|PT|784.43|ICD9CM|Hypernasality|Hypernasality
C0264614|T047|AB|784.43|ICD9CM|Hypernasality|Hypernasality
C0264618|T047|AB|784.44|ICD9CM|Hyponasality|Hyponasality
C0264618|T047|PT|784.44|ICD9CM|Hyponasality|Hyponasality
C2712366|T184|PT|784.49|ICD9CM|Other voice and resonance disorders|Other voice and resonance disorders
C2712366|T184|AB|784.49|ICD9CM|Voice/resonance dis NEC|Voice/resonance dis NEC
C0478144|T184|HT|784.5|ICD9CM|Other speech disturbance|Other speech disturbance
C0013362|T048|PT|784.51|ICD9CM|Dysarthria|Dysarthria
C0013362|T048|AB|784.51|ICD9CM|Dysarthria|Dysarthria
C2921127|T047|AB|784.52|ICD9CM|Flncy dsord cond elsewhr|Flncy dsord cond elsewhr
C2921127|T047|PT|784.52|ICD9CM|Fluency disorder in conditions classified elsewhere|Fluency disorder in conditions classified elsewhere
C2712367|T184|PT|784.59|ICD9CM|Other speech disturbance|Other speech disturbance
C2712367|T184|AB|784.59|ICD9CM|Speech disturbance NEC|Speech disturbance NEC
C0478145|T184|HT|784.6|ICD9CM|Other symbolic dysfunction|Other symbolic dysfunction
C0159047|T048|AB|784.60|ICD9CM|Symbolic dysfunction NOS|Symbolic dysfunction NOS
C0159047|T048|PT|784.60|ICD9CM|Symbolic dysfunction, unspecified|Symbolic dysfunction, unspecified
C0002019|T048|AB|784.61|ICD9CM|Alexia and dyslexia|Alexia and dyslexia
C0002019|T048|PT|784.61|ICD9CM|Alexia and dyslexia|Alexia and dyslexia
C0478145|T184|PT|784.69|ICD9CM|Other symbolic dysfunction|Other symbolic dysfunction
C0478145|T184|AB|784.69|ICD9CM|Symbolic dysfunction NEC|Symbolic dysfunction NEC
C0014591|T046|AB|784.7|ICD9CM|Epistaxis|Epistaxis
C0014591|T046|PT|784.7|ICD9CM|Epistaxis|Epistaxis
C0576995|T046|AB|784.8|ICD9CM|Hemorrhage from throat|Hemorrhage from throat
C0576995|T046|PT|784.8|ICD9CM|Hemorrhage from throat|Hemorrhage from throat
C0029855|T184|HT|784.9|ICD9CM|Other symptoms involving head and neck|Other symptoms involving head and neck
C0032781|T184|PT|784.91|ICD9CM|Postnasal drip|Postnasal drip
C0032781|T184|AB|784.91|ICD9CM|Postnasal drip|Postnasal drip
C0236000|T184|PT|784.92|ICD9CM|Jaw pain|Jaw pain
C0236000|T184|AB|784.92|ICD9CM|Jaw pain|Jaw pain
C0029855|T184|AB|784.99|ICD9CM|Head & neck symptoms NEC|Head & neck symptoms NEC
C0029855|T184|PT|784.99|ICD9CM|Other symptoms involving head and neck|Other symptoms involving head and neck
C0159049|T184|HT|785|ICD9CM|Symptoms involving cardiovascular system|Symptoms involving cardiovascular system
C0039231|T033|AB|785.0|ICD9CM|Tachycardia NOS|Tachycardia NOS
C0039231|T033|PT|785.0|ICD9CM|Tachycardia, unspecified|Tachycardia, unspecified
C0030252|T033|AB|785.1|ICD9CM|Palpitations|Palpitations
C0030252|T033|PT|785.1|ICD9CM|Palpitations|Palpitations
C0375546|T184|AB|785.2|ICD9CM|Cardiac murmurs NEC|Cardiac murmurs NEC
C0375546|T184|PT|785.2|ICD9CM|Undiagnosed cardiac murmurs|Undiagnosed cardiac murmurs
C0159050|T033|AB|785.3|ICD9CM|Abnorm heart sounds NEC|Abnorm heart sounds NEC
C0159050|T033|PT|785.3|ICD9CM|Other abnormal heart sounds|Other abnormal heart sounds
C0017086|T047|AB|785.4|ICD9CM|Gangrene|Gangrene
C0017086|T047|PT|785.4|ICD9CM|Gangrene|Gangrene
C0159051|T184|HT|785.5|ICD9CM|Shock without mention of trauma|Shock without mention of trauma
C0036974|T046|AB|785.50|ICD9CM|Shock NOS|Shock NOS
C0036974|T046|PT|785.50|ICD9CM|Shock, unspecified|Shock, unspecified
C0036980|T046|AB|785.51|ICD9CM|Cardiogenic shock|Cardiogenic shock
C0036980|T046|PT|785.51|ICD9CM|Cardiogenic shock|Cardiogenic shock
C0036983|T046|AB|785.52|ICD9CM|Septic shock|Septic shock
C0036983|T046|PT|785.52|ICD9CM|Septic shock|Septic shock
C0029737|T046|PT|785.59|ICD9CM|Other shock without mention of trauma|Other shock without mention of trauma
C0029737|T046|AB|785.59|ICD9CM|Shock w/o trauma NEC|Shock w/o trauma NEC
C4282165|T033|AB|785.6|ICD9CM|Enlargement lymph nodes|Enlargement lymph nodes
C4282165|T033|PT|785.6|ICD9CM|Enlargement of lymph nodes|Enlargement of lymph nodes
C0029854|T184|AB|785.9|ICD9CM|Cardiovas sys symp NEC|Cardiovas sys symp NEC
C0029854|T184|PT|785.9|ICD9CM|Other symptoms involving cardiovascular system|Other symptoms involving cardiovascular system
C0476271|T184|HT|786|ICD9CM|Symptoms involving respiratory system and other chest symptoms|Symptoms involving respiratory system and other chest symptoms
C0159053|T033|HT|786.0|ICD9CM|Dyspnea and respiratory abnormalities|Dyspnea and respiratory abnormalities
C1260922|T033|AB|786.00|ICD9CM|Respiratory abnorm NOS|Respiratory abnorm NOS
C1260922|T033|PT|786.00|ICD9CM|Respiratory abnormality, unspecified|Respiratory abnormality, unspecified
C0020578|T033|AB|786.01|ICD9CM|Hyperventilation|Hyperventilation
C0020578|T033|PT|786.01|ICD9CM|Hyperventilation|Hyperventilation
C0085619|T033|AB|786.02|ICD9CM|Orthopnea|Orthopnea
C0085619|T033|PT|786.02|ICD9CM|Orthopnea|Orthopnea
C0003578|T184|AB|786.03|ICD9CM|Apnea|Apnea
C0003578|T184|PT|786.03|ICD9CM|Apnea|Apnea
C0008039|T184|PT|786.04|ICD9CM|Cheyne-Stokes respiration|Cheyne-Stokes respiration
C0008039|T184|AB|786.04|ICD9CM|Cheyne-stokes respiratn|Cheyne-stokes respiratn
C0013404|T184|AB|786.05|ICD9CM|Shortness of breath|Shortness of breath
C0013404|T184|PT|786.05|ICD9CM|Shortness of breath|Shortness of breath
C0231835|T033|AB|786.06|ICD9CM|Tachypnea|Tachypnea
C0231835|T033|PT|786.06|ICD9CM|Tachypnea|Tachypnea
C0043144|T184|AB|786.07|ICD9CM|Wheezing|Wheezing
C0043144|T184|PT|786.07|ICD9CM|Wheezing|Wheezing
C0029601|T046|PT|786.09|ICD9CM|Other respiratory abnormalities|Other respiratory abnormalities
C0029601|T046|AB|786.09|ICD9CM|Respiratory abnorm NEC|Respiratory abnorm NEC
C0038450|T184|AB|786.1|ICD9CM|Stridor|Stridor
C0038450|T184|PT|786.1|ICD9CM|Stridor|Stridor
C0010200|T184|AB|786.2|ICD9CM|Cough|Cough
C0010200|T184|PT|786.2|ICD9CM|Cough|Cough
C0019079|T184|HT|786.3|ICD9CM|Hemoptysis|Hemoptysis
C0019079|T184|AB|786.30|ICD9CM|Hemoptysis NOS|Hemoptysis NOS
C0019079|T184|PT|786.30|ICD9CM|Hemoptysis, unspecified|Hemoptysis, unspecified
C2921130|T046|AB|786.31|ICD9CM|Ac idio pul hemrg infant|Ac idio pul hemrg infant
C2921130|T046|PT|786.31|ICD9CM|Acute idiopathic pulmonary hemorrhage in infants [AIPHI]|Acute idiopathic pulmonary hemorrhage in infants [AIPHI]
C2921131|T184|AB|786.39|ICD9CM|Hemoptysis NEC|Hemoptysis NEC
C2921131|T184|PT|786.39|ICD9CM|Other hemoptysis|Other hemoptysis
C0159054|T033|AB|786.4|ICD9CM|Abnormal sputum|Abnormal sputum
C0159054|T033|PT|786.4|ICD9CM|Abnormal sputum|Abnormal sputum
C0008031|T184|HT|786.5|ICD9CM|Chest pain|Chest pain
C0008031|T184|AB|786.50|ICD9CM|Chest pain NOS|Chest pain NOS
C0008031|T184|PT|786.50|ICD9CM|Chest pain, unspecified|Chest pain, unspecified
C0232286|T184|AB|786.51|ICD9CM|Precordial pain|Precordial pain
C0232286|T184|PT|786.51|ICD9CM|Precordial pain|Precordial pain
C0423729|T184|AB|786.52|ICD9CM|Painful respiration|Painful respiration
C0423729|T184|PT|786.52|ICD9CM|Painful respiration|Painful respiration
C0029537|T184|AB|786.59|ICD9CM|Chest pain NEC|Chest pain NEC
C0029537|T184|PT|786.59|ICD9CM|Other chest pain|Other chest pain
C0159055|T184|AB|786.6|ICD9CM|Chest swelling/mass/lump|Chest swelling/mass/lump
C0159055|T184|PT|786.6|ICD9CM|Swelling, mass, or lump in chest|Swelling, mass, or lump in chest
C0159056|T184|AB|786.7|ICD9CM|Abnormal chest sounds|Abnormal chest sounds
C0159056|T184|PT|786.7|ICD9CM|Abnormal chest sounds|Abnormal chest sounds
C0019521|T033|AB|786.8|ICD9CM|Hiccough|Hiccough
C0019521|T033|PT|786.8|ICD9CM|Hiccough|Hiccough
C0159057|T184|PT|786.9|ICD9CM|Other symptoms involving respiratory system and chest|Other symptoms involving respiratory system and chest
C0159057|T184|AB|786.9|ICD9CM|Resp sys/chest symp NEC|Resp sys/chest symp NEC
C0159058|T184|HT|787|ICD9CM|Symptoms involving digestive system|Symptoms involving digestive system
C0027498|T184|HT|787.0|ICD9CM|Nausea and vomiting|Nausea and vomiting
C0027498|T184|AB|787.01|ICD9CM|Nausea with vomiting|Nausea with vomiting
C0027498|T184|PT|787.01|ICD9CM|Nausea with vomiting|Nausea with vomiting
C0375548|T033|AB|787.02|ICD9CM|Nausea alone|Nausea alone
C0375548|T033|PT|787.02|ICD9CM|Nausea alone|Nausea alone
C0728950|T184|AB|787.03|ICD9CM|Vomiting alone|Vomiting alone
C0728950|T184|PT|787.03|ICD9CM|Vomiting alone|Vomiting alone
C0232599|T033|AB|787.04|ICD9CM|Bilious emesis|Bilious emesis
C0232599|T033|PT|787.04|ICD9CM|Bilious emesis|Bilious emesis
C0018834|T184|AB|787.1|ICD9CM|Heartburn|Heartburn
C0018834|T184|PT|787.1|ICD9CM|Heartburn|Heartburn
C0011168|T047|HT|787.2|ICD9CM|Dysphagia|Dysphagia
C0011168|T047|AB|787.20|ICD9CM|Dysphagia NOS|Dysphagia NOS
C0011168|T047|PT|787.20|ICD9CM|Dysphagia, unspecified|Dysphagia, unspecified
C2315800|T047|PT|787.21|ICD9CM|Dysphagia, oral phase|Dysphagia, oral phase
C2315800|T047|AB|787.21|ICD9CM|Dysphagia, oral phase|Dysphagia, oral phase
C0267071|T047|AB|787.22|ICD9CM|Dysphagia, oropharyngeal|Dysphagia, oropharyngeal
C0267071|T047|PT|787.22|ICD9CM|Dysphagia, oropharyngeal phase|Dysphagia, oropharyngeal phase
C1955516|T184|AB|787.23|ICD9CM|Dysphagia, pharyngeal|Dysphagia, pharyngeal
C1955516|T184|PT|787.23|ICD9CM|Dysphagia, pharyngeal phase|Dysphagia, pharyngeal phase
C1955517|T184|PT|787.24|ICD9CM|Dysphagia, pharyngoesophageal phase|Dysphagia, pharyngoesophageal phase
C1955517|T184|AB|787.24|ICD9CM|Dysphagia,pharyngoesoph|Dysphagia,pharyngoesoph
C1955518|T047|AB|787.29|ICD9CM|Dysphagia NEC|Dysphagia NEC
C1955518|T047|PT|787.29|ICD9CM|Other dysphagia|Other dysphagia
C0016205|T184|AB|787.3|ICD9CM|Flatul/eructat/gas pain|Flatul/eructat/gas pain
C0016205|T184|PT|787.3|ICD9CM|Flatulence, eructation, and gas pain|Flatulence, eructation, and gas pain
C0159059|T033|AB|787.4|ICD9CM|Visible peristalsis|Visible peristalsis
C0159059|T033|PT|787.4|ICD9CM|Visible peristalsis|Visible peristalsis
C0159060|T033|AB|787.5|ICD9CM|Abnormal bowel sounds|Abnormal bowel sounds
C0159060|T033|PT|787.5|ICD9CM|Abnormal bowel sounds|Abnormal bowel sounds
C0015732|T047|HT|787.6|ICD9CM|Incontinence of feces|Incontinence of feces
C2921132|T184|PT|787.60|ICD9CM|Full incontinence of feces|Full incontinence of feces
C2921132|T184|AB|787.60|ICD9CM|Full incontinence-feces|Full incontinence-feces
C0239167|T033|AB|787.61|ICD9CM|Incomplete defecation|Incomplete defecation
C0239167|T033|PT|787.61|ICD9CM|Incomplete defecation|Incomplete defecation
C4759678|T184|PT|787.62|ICD9CM|Fecal smearing|Fecal smearing
C4759678|T184|AB|787.62|ICD9CM|Fecal smearing|Fecal smearing
C0426636|T184|PT|787.63|ICD9CM|Fecal urgency|Fecal urgency
C0426636|T184|AB|787.63|ICD9CM|Fecal urgency|Fecal urgency
C0162287|T033|AB|787.7|ICD9CM|Abnormal feces|Abnormal feces
C0162287|T033|PT|787.7|ICD9CM|Abnormal feces|Abnormal feces
C0159061|T184|HT|787.9|ICD9CM|Other symptoms involving digestive system|Other symptoms involving digestive system
C0011991|T184|AB|787.91|ICD9CM|Diarrhea|Diarrhea
C0011991|T184|PT|787.91|ICD9CM|Diarrhea|Diarrhea
C0159061|T184|AB|787.99|ICD9CM|Digestve syst symptm NEC|Digestve syst symptm NEC
C0159061|T184|PT|787.99|ICD9CM|Other symptoms involving digestive system|Other symptoms involving digestive system
C0476293|T184|HT|788|ICD9CM|Symptoms involving urinary system|Symptoms involving urinary system
C0152169|T184|AB|788.0|ICD9CM|Renal colic|Renal colic
C0152169|T184|PT|788.0|ICD9CM|Renal colic|Renal colic
C0013428|T184|AB|788.1|ICD9CM|Dysuria|Dysuria
C0013428|T184|PT|788.1|ICD9CM|Dysuria|Dysuria
C0080274|T033|HT|788.2|ICD9CM|Retention of urine|Retention of urine
C0080274|T033|PT|788.20|ICD9CM|Retention of urine, unspecified|Retention of urine, unspecified
C0080274|T033|AB|788.20|ICD9CM|Retention urine NOS|Retention urine NOS
C0344365|T184|AB|788.21|ICD9CM|Incmplet bldder emptying|Incmplet bldder emptying
C0344365|T184|PT|788.21|ICD9CM|Incomplete bladder emptying|Incomplete bladder emptying
C0375549|T046|AB|788.29|ICD9CM|Oth spcf retention urine|Oth spcf retention urine
C0375549|T046|PT|788.29|ICD9CM|Other specified retention of urine|Other specified retention of urine
C0042024|T046|HT|788.3|ICD9CM|Urinary incontinence|Urinary incontinence
C0042024|T046|AB|788.30|ICD9CM|Urinary incontinence NOS|Urinary incontinence NOS
C0042024|T046|PT|788.30|ICD9CM|Urinary incontinence, unspecified|Urinary incontinence, unspecified
C0150045|T033|AB|788.31|ICD9CM|Urge incontinence|Urge incontinence
C0150045|T033|PT|788.31|ICD9CM|Urge incontinence|Urge incontinence
C0302505|T046|AB|788.32|ICD9CM|Stress incontinence male|Stress incontinence male
C0302505|T046|PT|788.32|ICD9CM|Stress incontinence, male|Stress incontinence, male
C0869256|T184|AB|788.33|ICD9CM|Mixed incontinence|Mixed incontinence
C0869256|T184|PT|788.33|ICD9CM|Mixed incontinence (male) (female)|Mixed incontinence (male) (female)
C0375551|T046|PT|788.34|ICD9CM|Incontinence without sensory awareness|Incontinence without sensory awareness
C0375551|T046|AB|788.34|ICD9CM|Incontnce wo sensr aware|Incontnce wo sensr aware
C0375552|T184|AB|788.35|ICD9CM|Post-void dribbling|Post-void dribbling
C0375552|T184|PT|788.35|ICD9CM|Post-void dribbling|Post-void dribbling
C0270327|T048|AB|788.36|ICD9CM|Nocturnal enuresis|Nocturnal enuresis
C0270327|T048|PT|788.36|ICD9CM|Nocturnal enuresis|Nocturnal enuresis
C0375553|T184|AB|788.37|ICD9CM|Continuous leakage|Continuous leakage
C0375553|T184|PT|788.37|ICD9CM|Continuous leakage|Continuous leakage
C0312413|T033|AB|788.38|ICD9CM|Overflow incontinence|Overflow incontinence
C0312413|T033|PT|788.38|ICD9CM|Overflow incontinence|Overflow incontinence
C0375554|T046|AB|788.39|ICD9CM|Oth urinry incontinence|Oth urinry incontinence
C0375554|T046|PT|788.39|ICD9CM|Other urinary incontinence|Other urinary incontinence
C0016708|T184|HT|788.4|ICD9CM|Frequency of urination and polyuria|Frequency of urination and polyuria
C0042023|T033|AB|788.41|ICD9CM|Urinary frequency|Urinary frequency
C0042023|T033|PT|788.41|ICD9CM|Urinary frequency|Urinary frequency
C0032617|T184|AB|788.42|ICD9CM|Polyuria|Polyuria
C0032617|T184|PT|788.42|ICD9CM|Polyuria|Polyuria
C0028734|T047|AB|788.43|ICD9CM|Nocturia|Nocturia
C0028734|T047|PT|788.43|ICD9CM|Nocturia|Nocturia
C0028962|T184|AB|788.5|ICD9CM|Oliguria & anuria|Oliguria & anuria
C0028962|T184|PT|788.5|ICD9CM|Oliguria and anuria|Oliguria and anuria
C0159063|T184|HT|788.6|ICD9CM|Other abnormality of urination|Other abnormality of urination
C0232855|T184|PT|788.61|ICD9CM|Splitting of urinary stream|Splitting of urinary stream
C0232855|T184|AB|788.61|ICD9CM|Splitting urinary stream|Splitting urinary stream
C0232854|T184|PT|788.62|ICD9CM|Slowing of urinary stream|Slowing of urinary stream
C0232854|T184|AB|788.62|ICD9CM|Slowing urinary stream|Slowing urinary stream
C0085606|T184|AB|788.63|ICD9CM|Urgency of urination|Urgency of urination
C0085606|T184|PT|788.63|ICD9CM|Urgency of urination|Urgency of urination
C0152032|T184|PT|788.64|ICD9CM|Urinary hesitancy|Urinary hesitancy
C0152032|T184|AB|788.64|ICD9CM|Urinary hesitancy|Urinary hesitancy
C0426365|T033|PT|788.65|ICD9CM|Straining on urination|Straining on urination
C0426365|T033|AB|788.65|ICD9CM|Straining on urination|Straining on urination
C0159063|T184|AB|788.69|ICD9CM|Oth abnormalt urination|Oth abnormalt urination
C0159063|T184|PT|788.69|ICD9CM|Other abnormality of urination|Other abnormality of urination
C0152447|T184|AB|788.7|ICD9CM|Urethral discharge|Urethral discharge
C0152447|T184|PT|788.7|ICD9CM|Urethral discharge|Urethral discharge
C0152245|T046|AB|788.8|ICD9CM|Extravasation of urine|Extravasation of urine
C0152245|T046|PT|788.8|ICD9CM|Extravasation of urine|Extravasation of urine
C0159064|T184|HT|788.9|ICD9CM|Other symptoms involving urinary system|Other symptoms involving urinary system
C0150042|T033|AB|788.91|ICD9CM|Fnctnl urinary incontnce|Fnctnl urinary incontnce
C0150042|T033|PT|788.91|ICD9CM|Functional urinary incontinence|Functional urinary incontinence
C0159064|T184|AB|788.99|ICD9CM|Oth symptm urinary systm|Oth symptm urinary systm
C0159064|T184|PT|788.99|ICD9CM|Other symptoms involving urinary system|Other symptoms involving urinary system
C0159065|T184|HT|789|ICD9CM|Other symptoms involving abdomen and pelvis|Other symptoms involving abdomen and pelvis
C0000737|T184|HT|789.0|ICD9CM|Abdominal pain|Abdominal pain
C0000737|T184|AB|789.00|ICD9CM|Abdmnal pain unspcf site|Abdmnal pain unspcf site
C0000737|T184|PT|789.00|ICD9CM|Abdominal pain, unspecified site|Abdominal pain, unspecified site
C0235299|T184|AB|789.01|ICD9CM|Abdmnal pain rt upr quad|Abdmnal pain rt upr quad
C0235299|T184|PT|789.01|ICD9CM|Abdominal pain, right upper quadrant|Abdominal pain, right upper quadrant
C0238552|T184|AB|789.02|ICD9CM|Abdmnal pain lft up quad|Abdmnal pain lft up quad
C0238552|T184|PT|789.02|ICD9CM|Abdominal pain, left upper quadrant|Abdominal pain, left upper quadrant
C0694551|T184|AB|789.03|ICD9CM|Abdmnal pain rt lwr quad|Abdmnal pain rt lwr quad
C0694551|T184|PT|789.03|ICD9CM|Abdominal pain, right lower quadrant|Abdominal pain, right lower quadrant
C0238551|T184|AB|789.04|ICD9CM|Abdmnal pain lt lwr quad|Abdmnal pain lt lwr quad
C0238551|T184|PT|789.04|ICD9CM|Abdominal pain, left lower quadrant|Abdominal pain, left lower quadrant
C1096624|T033|AB|789.05|ICD9CM|Abdmnal pain periumbilic|Abdmnal pain periumbilic
C1096624|T033|PT|789.05|ICD9CM|Abdominal pain, periumbilic|Abdominal pain, periumbilic
C0232493|T184|AB|789.06|ICD9CM|Abdmnal pain epigastric|Abdmnal pain epigastric
C0232493|T184|PT|789.06|ICD9CM|Abdominal pain, epigastric|Abdominal pain, epigastric
C0344304|T184|AB|789.07|ICD9CM|Abdmnal pain generalized|Abdmnal pain generalized
C0344304|T184|PT|789.07|ICD9CM|Abdominal pain, generalized|Abdominal pain, generalized
C0375555|T184|AB|789.09|ICD9CM|Abdmnal pain oth spcf st|Abdmnal pain oth spcf st
C0375555|T184|PT|789.09|ICD9CM|Abdominal pain, other specified site|Abdominal pain, other specified site
C0019209|T033|AB|789.1|ICD9CM|Hepatomegaly|Hepatomegaly
C0019209|T033|PT|789.1|ICD9CM|Hepatomegaly|Hepatomegaly
C0038002|T033|AB|789.2|ICD9CM|Splenomegaly|Splenomegaly
C0038002|T033|PT|789.2|ICD9CM|Splenomegaly|Splenomegaly
C0476310|T184|HT|789.3|ICD9CM|Abdominal or pelvic swelling, mass, or lump|Abdominal or pelvic swelling, mass, or lump
C0375556|T184|AB|789.30|ICD9CM|Abdmnal mass unspcf site|Abdmnal mass unspcf site
C0375556|T184|PT|789.30|ICD9CM|Abdominal or pelvic swelling, mass, or lump, unspecified site|Abdominal or pelvic swelling, mass, or lump, unspecified site
C0375557|T184|AB|789.31|ICD9CM|Abdmnal mass rt upr quad|Abdmnal mass rt upr quad
C0375557|T184|PT|789.31|ICD9CM|Abdominal or pelvic swelling, mass, or lump, right upper quadrant|Abdominal or pelvic swelling, mass, or lump, right upper quadrant
C0375558|T184|AB|789.32|ICD9CM|Abdmnal mass lft up quad|Abdmnal mass lft up quad
C0375558|T184|PT|789.32|ICD9CM|Abdominal or pelvic swelling, mass, or lump, left upper quadrant|Abdominal or pelvic swelling, mass, or lump, left upper quadrant
C0375559|T184|AB|789.33|ICD9CM|Abdmnal mass rt lwr quad|Abdmnal mass rt lwr quad
C0375559|T184|PT|789.33|ICD9CM|Abdominal or pelvic swelling, mass, or lump, right lower quadrant|Abdominal or pelvic swelling, mass, or lump, right lower quadrant
C0375560|T184|AB|789.34|ICD9CM|Abdmnal mass lt lwr quad|Abdmnal mass lt lwr quad
C0375560|T184|PT|789.34|ICD9CM|Abdominal or pelvic swelling, mass, or lump, left lower quadrant|Abdominal or pelvic swelling, mass, or lump, left lower quadrant
C0375561|T184|AB|789.35|ICD9CM|Abdmnal mass periumbilic|Abdmnal mass periumbilic
C0375561|T184|PT|789.35|ICD9CM|Abdominal or pelvic swelling, mass, or lump, periumbilic|Abdominal or pelvic swelling, mass, or lump, periumbilic
C0375562|T184|AB|789.36|ICD9CM|Abdmnal mass epigastric|Abdmnal mass epigastric
C0375562|T184|PT|789.36|ICD9CM|Abdominal or pelvic swelling, mass, or lump, epigastric|Abdominal or pelvic swelling, mass, or lump, epigastric
C0375563|T184|AB|789.37|ICD9CM|Abdmnal mass generalized|Abdmnal mass generalized
C0375563|T184|PT|789.37|ICD9CM|Abdominal or pelvic swelling, mass, or lump, generalized|Abdominal or pelvic swelling, mass, or lump, generalized
C0375564|T184|AB|789.39|ICD9CM|Abdmnal mass oth spcf st|Abdmnal mass oth spcf st
C0375564|T184|PT|789.39|ICD9CM|Abdominal or pelvic swelling, mass, or lump, other specified site|Abdominal or pelvic swelling, mass, or lump, other specified site
C0159066|T184|HT|789.4|ICD9CM|Abdominal rigidity|Abdominal rigidity
C0159066|T184|AB|789.40|ICD9CM|Abdmnal rgdt unspcf site|Abdmnal rgdt unspcf site
C0159066|T184|PT|789.40|ICD9CM|Abdominal rigidity, unspecified site|Abdominal rigidity, unspecified site
C0375565|T184|AB|789.41|ICD9CM|Abdmnal rgdt rt upr quad|Abdmnal rgdt rt upr quad
C0375565|T184|PT|789.41|ICD9CM|Abdominal rigidity, right upper quadrant|Abdominal rigidity, right upper quadrant
C2585165|T184|AB|789.42|ICD9CM|Abdmnal rgdt lft up quad|Abdmnal rgdt lft up quad
C2585165|T184|PT|789.42|ICD9CM|Abdominal rigidity, left upper quadrant|Abdominal rigidity, left upper quadrant
C2585545|T184|AB|789.43|ICD9CM|Abdmnal rgdt rt lwr quad|Abdmnal rgdt rt lwr quad
C2585545|T184|PT|789.43|ICD9CM|Abdominal rigidity, right lower quadrant|Abdominal rigidity, right lower quadrant
C2585546|T184|AB|789.44|ICD9CM|Abdmnal rgdt lt lwr quad|Abdmnal rgdt lt lwr quad
C2585546|T184|PT|789.44|ICD9CM|Abdominal rigidity, left lower quadrant|Abdominal rigidity, left lower quadrant
C2127287|T033|AB|789.45|ICD9CM|Abdmnal rgdt periumbilic|Abdmnal rgdt periumbilic
C2127287|T033|PT|789.45|ICD9CM|Abdominal rigidity, periumbilic|Abdominal rigidity, periumbilic
C0375570|T184|AB|789.46|ICD9CM|Abdmnal rgdt epigastric|Abdmnal rgdt epigastric
C0375570|T184|PT|789.46|ICD9CM|Abdominal rigidity, epigastric|Abdominal rigidity, epigastric
C0375571|T184|AB|789.47|ICD9CM|Abdmnal rgdt generalized|Abdmnal rgdt generalized
C0375571|T184|PT|789.47|ICD9CM|Abdominal rigidity, generalized|Abdominal rigidity, generalized
C0375572|T184|AB|789.49|ICD9CM|Abdmnal rgdt oth spcf st|Abdmnal rgdt oth spcf st
C0375572|T184|PT|789.49|ICD9CM|Abdominal rigidity, other specified site|Abdominal rigidity, other specified site
C0003962|T047|HT|789.5|ICD9CM|Ascites|Ascites
C0220656|T191|PT|789.51|ICD9CM|Malignant ascites|Malignant ascites
C0220656|T191|AB|789.51|ICD9CM|Malignant ascites|Malignant ascites
C1955521|T047|AB|789.59|ICD9CM|Ascites NEC|Ascites NEC
C1955521|T047|PT|789.59|ICD9CM|Other ascites|Other ascites
C0232498|T184|HT|789.6|ICD9CM|Abdominal tenderness|Abdominal tenderness
C0232498|T184|AB|789.60|ICD9CM|Abdmnal tndr unspcf site|Abdmnal tndr unspcf site
C0232498|T184|PT|789.60|ICD9CM|Abdominal tenderness, unspecified site|Abdominal tenderness, unspecified site
C0238571|T184|AB|789.61|ICD9CM|Abdmnal tndr rt upr quad|Abdmnal tndr rt upr quad
C0238571|T184|PT|789.61|ICD9CM|Abdominal tenderness, right upper quadrant|Abdominal tenderness, right upper quadrant
C0238566|T184|AB|789.62|ICD9CM|Abdmnal tndr lft up quad|Abdmnal tndr lft up quad
C0238566|T184|PT|789.62|ICD9CM|Abdominal tenderness, left upper quadrant|Abdominal tenderness, left upper quadrant
C0238570|T184|AB|789.63|ICD9CM|Abdmnal tndr rt lwr quad|Abdmnal tndr rt lwr quad
C0238570|T184|PT|789.63|ICD9CM|Abdominal tenderness, right lower quadrant|Abdominal tenderness, right lower quadrant
C2585306|T184|AB|789.64|ICD9CM|Abdmnal tndr lt lwr quad|Abdmnal tndr lt lwr quad
C2585306|T184|PT|789.64|ICD9CM|Abdominal tenderness, left lower quadrant|Abdominal tenderness, left lower quadrant
C0375573|T184|AB|789.65|ICD9CM|Abdmnal tndr periumbilic|Abdmnal tndr periumbilic
C0375573|T184|PT|789.65|ICD9CM|Abdominal tenderness, periumbilic|Abdominal tenderness, periumbilic
C0239280|T184|AB|789.66|ICD9CM|Abdmnal tndr epigastric|Abdmnal tndr epigastric
C0239280|T184|PT|789.66|ICD9CM|Abdominal tenderness, epigastric|Abdominal tenderness, epigastric
C0302540|T184|AB|789.67|ICD9CM|Abdmnal tndr generalized|Abdmnal tndr generalized
C0302540|T184|PT|789.67|ICD9CM|Abdominal tenderness, generalized|Abdominal tenderness, generalized
C0375574|T184|AB|789.69|ICD9CM|Abdmnal tndr oth spcf st|Abdmnal tndr oth spcf st
C0375574|T184|PT|789.69|ICD9CM|Abdominal tenderness, other specified site|Abdominal tenderness, other specified site
C0232488|T033|PT|789.7|ICD9CM|Colic|Colic
C0232488|T033|AB|789.7|ICD9CM|Colic|Colic
C0159065|T184|AB|789.9|ICD9CM|Abdomen/pelvis symp NEC|Abdomen/pelvis symp NEC
C0159065|T184|PT|789.9|ICD9CM|Other symptoms involving abdomen and pelvis|Other symptoms involving abdomen and pelvis
C0476319|T033|HT|790|ICD9CM|Nonspecific findings on examination of blood|Nonspecific findings on examination of blood
C2004518|T033|HT|790-796.99|ICD9CM|NONSPECIFIC ABNORMAL FINDINGS|NONSPECIFIC ABNORMAL FINDINGS
C0391870|T033|HT|790.0|ICD9CM|Abnormality of red blood cells|Abnormality of red blood cells
C0878707|T184|AB|790.01|ICD9CM|Drop, hematocrit, precip|Drop, hematocrit, precip
C0878707|T184|PT|790.01|ICD9CM|Precipitous drop in hematocrit|Precipitous drop in hematocrit
C0878708|T033|AB|790.09|ICD9CM|Abnormal RBC NEC|Abnormal RBC NEC
C0878708|T033|PT|790.09|ICD9CM|Other abnormality of red blood cells|Other abnormality of red blood cells
C0151632|T033|AB|790.1|ICD9CM|Elevated sediment rate|Elevated sediment rate
C0151632|T033|PT|790.1|ICD9CM|Elevated sedimentation rate|Elevated sedimentation rate
C0580546|T033|HT|790.2|ICD9CM|Abnormal glucose|Abnormal glucose
C1272092|T033|AB|790.21|ICD9CM|Impaired fasting glucose|Impaired fasting glucose
C1272092|T033|PT|790.21|ICD9CM|Impaired fasting glucose|Impaired fasting glucose
C2830475|T033|PT|790.22|ICD9CM|Impaired glucose tolerance test (oral)|Impaired glucose tolerance test (oral)
C2830475|T033|AB|790.22|ICD9CM|Impaired oral glucse tol|Impaired oral glucse tol
C1260443|T033|AB|790.29|ICD9CM|Abnormal glucose NEC|Abnormal glucose NEC
C1260443|T033|PT|790.29|ICD9CM|Other abnormal glucose|Other abnormal glucose
C0159070|T033|AB|790.3|ICD9CM|Excess blood-alcohol lev|Excess blood-alcohol lev
C0159070|T033|PT|790.3|ICD9CM|Excessive blood level of alcohol|Excessive blood level of alcohol
C0159071|T033|AB|790.4|ICD9CM|Elev transaminase/ldh|Elev transaminase/ldh
C0159071|T033|PT|790.4|ICD9CM|Nonspecific elevation of levels of transaminase or lactic acid dehydrogenase [LDH]|Nonspecific elevation of levels of transaminase or lactic acid dehydrogenase [LDH]
C0159072|T046|AB|790.5|ICD9CM|Abn serum enzy level NEC|Abn serum enzy level NEC
C0159072|T046|PT|790.5|ICD9CM|Other nonspecific abnormal serum enzyme levels|Other nonspecific abnormal serum enzyme levels
C0029481|T046|AB|790.6|ICD9CM|Abn blood chemistry NEC|Abn blood chemistry NEC
C0029481|T046|PT|790.6|ICD9CM|Other abnormal blood chemistry|Other abnormal blood chemistry
C0004610|T047|AB|790.7|ICD9CM|Bacteremia|Bacteremia
C0004610|T047|PT|790.7|ICD9CM|Bacteremia|Bacteremia
C0042749|T047|AB|790.8|ICD9CM|Viremia NOS|Viremia NOS
C0042749|T047|PT|790.8|ICD9CM|Viremia, unspecified|Viremia, unspecified
C0159073|T033|HT|790.9|ICD9CM|Other nonspecific findings on examination of blood|Other nonspecific findings on examination of blood
C0375575|T033|PT|790.91|ICD9CM|Abnormal arterial blood gases|Abnormal arterial blood gases
C0375575|T033|AB|790.91|ICD9CM|Abnrml art blood gases|Abnrml art blood gases
C0375576|T033|PT|790.92|ICD9CM|Abnormal coagulation profile|Abnormal coagulation profile
C0375576|T033|AB|790.92|ICD9CM|Abnrml coagultion prfile|Abnrml coagultion prfile
C0178415|T033|PT|790.93|ICD9CM|Elevated prostate specific antigen [PSA]|Elevated prostate specific antigen [PSA]
C0178415|T033|AB|790.93|ICD9CM|Elvtd prstate spcf antgn|Elvtd prstate spcf antgn
C0015190|T047|AB|790.94|ICD9CM|Euthyroid sick syndrome|Euthyroid sick syndrome
C0015190|T047|PT|790.94|ICD9CM|Euthyroid sick syndrome|Euthyroid sick syndrome
C1455884|T033|AB|790.95|ICD9CM|Elev C-reactive protein|Elev C-reactive protein
C1455884|T033|PT|790.95|ICD9CM|Elevated C-reactive protein (CRP)|Elevated C-reactive protein (CRP)
C0159073|T033|AB|790.99|ICD9CM|Oth nspcf finding blood|Oth nspcf finding blood
C0159073|T033|PT|790.99|ICD9CM|Other nonspecific findings on examination of blood|Other nonspecific findings on examination of blood
C0476338|T033|HT|791|ICD9CM|Nonspecific findings on examination of urine|Nonspecific findings on examination of urine
C0033687|T033|AB|791.0|ICD9CM|Proteinuria|Proteinuria
C0033687|T033|PT|791.0|ICD9CM|Proteinuria|Proteinuria
C0159075|T184|AB|791.1|ICD9CM|Chyluria|Chyluria
C0159075|T184|PT|791.1|ICD9CM|Chyluria|Chyluria
C0019048|T033|AB|791.2|ICD9CM|Hemoglobinuria|Hemoglobinuria
C0019048|T033|PT|791.2|ICD9CM|Hemoglobinuria|Hemoglobinuria
C0027080|T033|AB|791.3|ICD9CM|Myoglobinuria|Myoglobinuria
C0027080|T033|PT|791.3|ICD9CM|Myoglobinuria|Myoglobinuria
C0159076|T033|AB|791.4|ICD9CM|Biliuria|Biliuria
C0159076|T033|PT|791.4|ICD9CM|Biliuria|Biliuria
C0017979|T033|AB|791.5|ICD9CM|Glycosuria|Glycosuria
C0017979|T033|PT|791.5|ICD9CM|Glycosuria|Glycosuria
C0162275|T047|AB|791.6|ICD9CM|Acetonuria|Acetonuria
C0162275|T047|PT|791.6|ICD9CM|Acetonuria|Acetonuria
C0159077|T033|AB|791.7|ICD9CM|Oth cells/casts in urine|Oth cells/casts in urine
C0159077|T033|PT|791.7|ICD9CM|Other cells and casts in urine|Other cells and casts in urine
C0159078|T033|AB|791.9|ICD9CM|Abn urine findings NEC|Abn urine findings NEC
C0159078|T033|PT|791.9|ICD9CM|Other nonspecific findings on examination of urine|Other nonspecific findings on examination of urine
C0159079|T033|HT|792|ICD9CM|Nonspecific abnormal findings in other body substances|Nonspecific abnormal findings in other body substances
C0151583|T033|AB|792.0|ICD9CM|Abn fnd-cerebrospinal fl|Abn fnd-cerebrospinal fl
C0151583|T033|PT|792.0|ICD9CM|Nonspecific abnormal findings in cerebrospinal fluid|Nonspecific abnormal findings in cerebrospinal fluid
C0476346|T033|AB|792.1|ICD9CM|Abn find-stool contents|Abn find-stool contents
C0476346|T033|PT|792.1|ICD9CM|Nonspecific abnormal findings in stool contents|Nonspecific abnormal findings in stool contents
C0235756|T033|AB|792.2|ICD9CM|Abn findings-semen|Abn findings-semen
C0235756|T033|PT|792.2|ICD9CM|Nonspecific abnormal findings in semen|Nonspecific abnormal findings in semen
C0266781|T033|AB|792.3|ICD9CM|Abn find-amniotic fluid|Abn find-amniotic fluid
C0266781|T033|PT|792.3|ICD9CM|Nonspecific abnormal findings in amniotic fluid|Nonspecific abnormal findings in amniotic fluid
C0159084|T033|AB|792.4|ICD9CM|Abn findings-saliva|Abn findings-saliva
C0159084|T033|PT|792.4|ICD9CM|Nonspecific abnormal findings in saliva|Nonspecific abnormal findings in saliva
C0878709|T184|PT|792.5|ICD9CM|Cloudy (hemodialysis) (peritoneal) dialysis effluent|Cloudy (hemodialysis) (peritoneal) dialysis effluent
C0878709|T184|AB|792.5|ICD9CM|Cloudy dialysis effluent|Cloudy dialysis effluent
C0159079|T033|AB|792.9|ICD9CM|Abn find-body subst NEC|Abn find-body subst NEC
C0159079|T033|PT|792.9|ICD9CM|Other nonspecific abnormal findings in body substances|Other nonspecific abnormal findings in body substances
C0159085|T033|HT|793|ICD9CM|Nonspecific (abnormal) findings on radiological and other examination of body structure|Nonspecific (abnormal) findings on radiological and other examination of body structure
C0476359|T033|AB|793.0|ICD9CM|Nonsp abn fd-skull/head|Nonsp abn fd-skull/head
C0476359|T033|PT|793.0|ICD9CM|Nonspecific (abnormal) findings on radiological and other examination of skull and head|Nonspecific (abnormal) findings on radiological and other examination of skull and head
C0476365|T033|HT|793.1|ICD9CM|Nonspecific abnormal findings on radiological and other examination of lung field|Nonspecific abnormal findings on radiological and other examination of lung field
C2350019|T191|PT|793.11|ICD9CM|Solitary pulmonary nodule|Solitary pulmonary nodule
C2350019|T191|AB|793.11|ICD9CM|Solitary pulmonry nodule|Solitary pulmonry nodule
C3161126|T033|AB|793.19|ICD9CM|Ot nonsp ab fnd lung fld|Ot nonsp ab fnd lung fld
C3161126|T033|PT|793.19|ICD9CM|Other nonspecific abnormal finding of lung field|Other nonspecific abnormal finding of lung field
C0159088|T033|AB|793.2|ICD9CM|Nonsp abn intrathor NEC|Nonsp abn intrathor NEC
C0159088|T033|PT|793.2|ICD9CM|Nonspecific (abnormal) findings on radiological and other examination of other intrathoracic organs|Nonspecific (abnormal) findings on radiological and other examination of other intrathoracic organs
C0159089|T033|AB|793.3|ICD9CM|Nonsp abn fd-bilry tract|Nonsp abn fd-bilry tract
C0159089|T033|PT|793.3|ICD9CM|Nonspecific (abnormal) findings on radiological and other examination of biliary tract|Nonspecific (abnormal) findings on radiological and other examination of biliary tract
C0159090|T033|AB|793.4|ICD9CM|Nonsp abn find-gi tract|Nonsp abn find-gi tract
C0159090|T033|PT|793.4|ICD9CM|Nonspecific (abnormal) findings on radiological and other examination of gastrointestinal tract|Nonspecific (abnormal) findings on radiological and other examination of gastrointestinal tract
C0476376|T033|AB|793.5|ICD9CM|Nonsp abn find-gu organs|Nonsp abn find-gu organs
C0476376|T033|PT|793.5|ICD9CM|Nonspecific (abnormal) findings on radiological and other examination of genitourinary organs|Nonspecific (abnormal) findings on radiological and other examination of genitourinary organs
C0159092|T033|AB|793.6|ICD9CM|Nonsp abn fnd-abdom area|Nonsp abn fnd-abdom area
C0159093|T033|AB|793.7|ICD9CM|Nonsp abn find-ms system|Nonsp abn find-ms system
C0159093|T033|PT|793.7|ICD9CM|Nonspecific (abnormal) findings on radiological and other examination of musculoskeletal system|Nonspecific (abnormal) findings on radiological and other examination of musculoskeletal system
C0159094|T033|HT|793.8|ICD9CM|Nonspecific abnormal findings on radiological and other examination of breast|Nonspecific abnormal findings on radiological and other examination of breast
C0949146|T047|AB|793.80|ICD9CM|Ab mammogram NOS|Ab mammogram NOS
C0949146|T047|PT|793.80|ICD9CM|Abnormal mammogram, unspecified|Abnormal mammogram, unspecified
C2830589|T033|AB|793.81|ICD9CM|Mammographic microcalcif|Mammographic microcalcif
C2830589|T033|PT|793.81|ICD9CM|Mammographic microcalcification|Mammographic microcalcification
C2712369|T033|PT|793.82|ICD9CM|Inconclusive mammogram|Inconclusive mammogram
C2712369|T033|AB|793.82|ICD9CM|Inconclusive mammogram|Inconclusive mammogram
C0949148|T047|AB|793.89|ICD9CM|Abn finding-breast NEC|Abn finding-breast NEC
C0949148|T047|PT|793.89|ICD9CM|Other (abnormal) findings on radiological examination of breast|Other (abnormal) findings on radiological examination of breast
C0028315|T033|HT|793.9|ICD9CM|Nonspecific abnormal findings on radiological and other examination of other sites of body|Nonspecific abnormal findings on radiological and other examination of other sites of body
C1719644|T033|AB|793.91|ICD9CM|Image test incon d/t fat|Image test incon d/t fat
C1719644|T033|PT|793.91|ICD9CM|Image test inconclusive due to excess body fat|Image test inconclusive due to excess body fat
C1719645|T033|AB|793.99|ICD9CM|Nonsp abn find-body NEC|Nonsp abn find-body NEC
C1719645|T033|PT|793.99|ICD9CM|Other nonspecific (abnormal) findings on radiological and other examinations of body structure|Other nonspecific (abnormal) findings on radiological and other examinations of body structure
C0476388|T033|HT|794|ICD9CM|Nonspecific abnormal results of function studies|Nonspecific abnormal results of function studies
C0476389|T033|HT|794.0|ICD9CM|Nonspecific abnormal results of function study of brain and central nervous system|Nonspecific abnormal results of function study of brain and central nervous system
C0476389|T033|AB|794.00|ICD9CM|Abn cns funct study NOS|Abn cns funct study NOS
C0476389|T033|PT|794.00|ICD9CM|Abnormal function study of brain and central nervous system, unspecified|Abnormal function study of brain and central nervous system, unspecified
C0476391|T033|AB|794.01|ICD9CM|Abnorm echoencephalogram|Abnorm echoencephalogram
C0476391|T033|PT|794.01|ICD9CM|Nonspecific abnormal echoencephalogram|Nonspecific abnormal echoencephalogram
C0159099|T033|AB|794.02|ICD9CM|Abn electroencephalogram|Abn electroencephalogram
C0159099|T033|PT|794.02|ICD9CM|Nonspecific abnormal electroencephalogram [EEG]|Nonspecific abnormal electroencephalogram [EEG]
C0159100|T033|AB|794.09|ICD9CM|Abn cns funct study NEC|Abn cns funct study NEC
C0159100|T033|PT|794.09|ICD9CM|Other nonspecific abnormal results of function study of brain and central nervous system|Other nonspecific abnormal results of function study of brain and central nervous system
C0495795|T033|HT|794.1|ICD9CM|Nonspecific abnormal results of function study of peripheral nervous system and special senses|Nonspecific abnormal results of function study of peripheral nervous system and special senses
C0159102|T033|AB|794.10|ICD9CM|Abn stimul response NOS|Abn stimul response NOS
C0159102|T033|PT|794.10|ICD9CM|Nonspecific abnormal response to nerve stimulation, unspecified|Nonspecific abnormal response to nerve stimulation, unspecified
C0476396|T033|AB|794.11|ICD9CM|Abn retinal funct study|Abn retinal funct study
C0476396|T033|PT|794.11|ICD9CM|Nonspecific abnormal retinal function studies|Nonspecific abnormal retinal function studies
C0159104|T033|AB|794.12|ICD9CM|Abnorm electro-oculogram|Abnorm electro-oculogram
C0159104|T033|PT|794.12|ICD9CM|Nonspecific abnormal electro-oculogram [EOG]|Nonspecific abnormal electro-oculogram [EOG]
C0522214|T033|AB|794.13|ICD9CM|Abnormal vep|Abnormal vep
C0522214|T033|PT|794.13|ICD9CM|Nonspecific abnormal visually evoked potential|Nonspecific abnormal visually evoked potential
C0159106|T033|AB|794.14|ICD9CM|Abn oculomotor studies|Abn oculomotor studies
C0159106|T033|PT|794.14|ICD9CM|Nonspecific abnormal oculomotor studies|Nonspecific abnormal oculomotor studies
C0159107|T033|AB|794.15|ICD9CM|Abn auditory funct study|Abn auditory funct study
C0159107|T033|PT|794.15|ICD9CM|Nonspecific abnormal auditory function studies|Nonspecific abnormal auditory function studies
C0476402|T033|AB|794.16|ICD9CM|Abn vestibular func stud|Abn vestibular func stud
C0476402|T033|PT|794.16|ICD9CM|Nonspecific abnormal vestibular function studies|Nonspecific abnormal vestibular function studies
C0476403|T033|AB|794.17|ICD9CM|Abnorm electromyogram|Abnorm electromyogram
C0476403|T033|PT|794.17|ICD9CM|Nonspecific abnormal electromyogram [EMG]|Nonspecific abnormal electromyogram [EMG]
C0159110|T033|AB|794.19|ICD9CM|Abn periph nerv stud NEC|Abn periph nerv stud NEC
C0159110|T033|PT|794.19|ICD9CM|Other nonspecific abnormal results of function study of peripheral nervous system and special senses|Other nonspecific abnormal results of function study of peripheral nervous system and special senses
C0476405|T033|AB|794.2|ICD9CM|Abn pulmonary func study|Abn pulmonary func study
C0476405|T033|PT|794.2|ICD9CM|Nonspecific abnormal results of pulmonary function study|Nonspecific abnormal results of pulmonary function study
C0476409|T033|HT|794.3|ICD9CM|Nonspecific abnormal results of function study, cardiovascular|Nonspecific abnormal results of function study, cardiovascular
C0476409|T033|AB|794.30|ICD9CM|Abn cardiovasc study NOS|Abn cardiovasc study NOS
C0476409|T033|PT|794.30|ICD9CM|Abnormal cardiovascular function study, unspecified|Abnormal cardiovascular function study, unspecified
C0236140|T033|AB|794.31|ICD9CM|Abnorm electrocardiogram|Abnorm electrocardiogram
C0236140|T033|PT|794.31|ICD9CM|Nonspecific abnormal electrocardiogram [ECG] [EKG]|Nonspecific abnormal electrocardiogram [ECG] [EKG]
C2711989|T033|AB|794.39|ICD9CM|Abn cardiovasc study NEC|Abn cardiovasc study NEC
C2711989|T033|PT|794.39|ICD9CM|Other nonspecific abnormal results of function study of cardiovascular system|Other nonspecific abnormal results of function study of cardiovascular system
C0236151|T033|AB|794.4|ICD9CM|Abn kidney funct study|Abn kidney funct study
C0236151|T033|PT|794.4|ICD9CM|Nonspecific abnormal results of function study of kidney|Nonspecific abnormal results of function study of kidney
C0476414|T033|AB|794.5|ICD9CM|Abn thyroid funct study|Abn thyroid funct study
C0476414|T033|PT|794.5|ICD9CM|Nonspecific abnormal results of function study of thyroid|Nonspecific abnormal results of function study of thyroid
C0159117|T033|AB|794.6|ICD9CM|Abn endocrine study NEC|Abn endocrine study NEC
C0159117|T033|PT|794.6|ICD9CM|Nonspecific abnormal results of other endocrine function study|Nonspecific abnormal results of other endocrine function study
C0159118|T033|AB|794.7|ICD9CM|Abn basal metabol study|Abn basal metabol study
C0159118|T033|PT|794.7|ICD9CM|Nonspecific abnormal results of function study of basal metabolism|Nonspecific abnormal results of function study of basal metabolism
C0151766|T033|AB|794.8|ICD9CM|Abn liver function study|Abn liver function study
C0151766|T033|PT|794.8|ICD9CM|Nonspecific abnormal results of function study of liver|Nonspecific abnormal results of function study of liver
C0159120|T033|AB|794.9|ICD9CM|Abn function study NEC|Abn function study NEC
C0159120|T033|PT|794.9|ICD9CM|Nonspecific abnormal results of other specified function study|Nonspecific abnormal results of other specified function study
C1455902|T033|HT|795|ICD9CM|Other and nonspecific abnormal cytological, histological, immunological and DNA test findings|Other and nonspecific abnormal cytological, histological, immunological and DNA test findings
C1455899|T033|HT|795.0|ICD9CM|Abnormal Papanicolaou smear of cervix and cervical HPV|Abnormal Papanicolaou smear of cervix and cervical HPV
C1455885|T033|AB|795.00|ICD9CM|Abn glandular pap smear|Abn glandular pap smear
C1455885|T033|PT|795.00|ICD9CM|Abnormal glandular Papanicolaou smear of cervix|Abnormal glandular Papanicolaou smear of cervix
C1455889|T033|AB|795.01|ICD9CM|Pap smear (ASC-US)|Pap smear (ASC-US)
C1455889|T033|PT|795.01|ICD9CM|Papanicolaou smear of cervix with atypical squamous cells of undetermined significance (ASC-US)|Papanicolaou smear of cervix with atypical squamous cells of undetermined significance (ASC-US)
C1455890|T033|AB|795.02|ICD9CM|Pap smear (ASC-H)|Pap smear (ASC-H)
C1455891|T033|AB|795.03|ICD9CM|Pap smear cervix w LGSIL|Pap smear cervix w LGSIL
C1455891|T033|PT|795.03|ICD9CM|Papanicolaou smear of cervix with low grade squamous intraepithelial lesion (LGSIL)|Papanicolaou smear of cervix with low grade squamous intraepithelial lesion (LGSIL)
C1455892|T033|AB|795.04|ICD9CM|Pap smear cervix w HGSIL|Pap smear cervix w HGSIL
C1455892|T033|PT|795.04|ICD9CM|Papanicolaou smear of cervix with high grade squamous intraepithelial lesion (HGSIL)|Papanicolaou smear of cervix with high grade squamous intraepithelial lesion (HGSIL)
C1455894|T033|AB|795.05|ICD9CM|Cervical (HPV) DNA pos|Cervical (HPV) DNA pos
C1455894|T033|PT|795.05|ICD9CM|Cervical high risk human papillomavirus (HPV) DNA test positive|Cervical high risk human papillomavirus (HPV) DNA test positive
C1719648|T033|AB|795.06|ICD9CM|Pap smr cytol evid malig|Pap smr cytol evid malig
C1719648|T033|PT|795.06|ICD9CM|Papanicolaou smear of cervix with cytologic evidence of malignancy|Papanicolaou smear of cervix with cytologic evidence of malignancy
C2349680|T033|AB|795.07|ICD9CM|Sat cerv smr-no trnsfrm|Sat cerv smr-no trnsfrm
C2349680|T033|PT|795.07|ICD9CM|Satisfactory cervical smear but lacking transformation zone|Satisfactory cervical smear but lacking transformation zone
C2349681|T033|AB|795.08|ICD9CM|Unsat cerv cytlogy smear|Unsat cerv cytlogy smear
C2349681|T033|PT|795.08|ICD9CM|Unsatisfactory cervical cytology smear|Unsatisfactory cervical cytology smear
C1455897|T047|AB|795.09|ICD9CM|Abn pap cervix HPV NEC|Abn pap cervix HPV NEC
C1455897|T047|PT|795.09|ICD9CM|Other abnormal Papanicolaou smear of cervix and cervical HPV|Other abnormal Papanicolaou smear of cervix and cervical HPV
C2349696|T033|HT|795.1|ICD9CM|Abnormal Papanicolaou smear of vagina and vaginal HPV|Abnormal Papanicolaou smear of vagina and vaginal HPV
C2349683|T033|AB|795.10|ICD9CM|Abn gland pap smr vagina|Abn gland pap smr vagina
C2349683|T033|PT|795.10|ICD9CM|Abnormal glandular Papanicolaou smear of vagina|Abnormal glandular Papanicolaou smear of vagina
C2349685|T033|AB|795.11|ICD9CM|Pap smear vag w ASC-US|Pap smear vag w ASC-US
C2349685|T033|PT|795.11|ICD9CM|Papanicolaou smear of vagina with atypical squamous cells of undetermined significance (ASC-US)|Papanicolaou smear of vagina with atypical squamous cells of undetermined significance (ASC-US)
C2349686|T033|AB|795.12|ICD9CM|Pap smear vagina w ASC-H|Pap smear vagina w ASC-H
C2349687|T033|AB|795.13|ICD9CM|Pap smear vagina w LGSIL|Pap smear vagina w LGSIL
C2349687|T033|PT|795.13|ICD9CM|Papanicolaou smear of vagina with low grade squamous intraepithelial lesion (LGSIL)|Papanicolaou smear of vagina with low grade squamous intraepithelial lesion (LGSIL)
C2349688|T033|AB|795.14|ICD9CM|Pap smear vagina w HGSIL|Pap smear vagina w HGSIL
C2349688|T033|PT|795.14|ICD9CM|Papanicolaou smear of vagina with high grade squamous intraepithelial lesion (HGSIL)|Papanicolaou smear of vagina with high grade squamous intraepithelial lesion (HGSIL)
C2349689|T033|AB|795.15|ICD9CM|Vag hi risk HPV-DNA pos|Vag hi risk HPV-DNA pos
C2349689|T033|PT|795.15|ICD9CM|Vaginal high risk human papillomavirus (HPV) DNA test positive|Vaginal high risk human papillomavirus (HPV) DNA test positive
C2349690|T033|AB|795.16|ICD9CM|Pap smr vag-cytol malig|Pap smr vag-cytol malig
C2349690|T033|PT|795.16|ICD9CM|Papanicolaou smear of vagina with cytologic evidence of malignancy|Papanicolaou smear of vagina with cytologic evidence of malignancy
C2830555|T033|PT|795.18|ICD9CM|Unsatisfactory vaginal cytology smear|Unsatisfactory vaginal cytology smear
C2830555|T033|AB|795.18|ICD9CM|Vaginl cytol smr unsatis|Vaginl cytol smr unsatis
C2349693|T033|AB|795.19|ICD9CM|Oth abn Pap smr vag/HPV|Oth abn Pap smr vag/HPV
C2349693|T033|PT|795.19|ICD9CM|Other abnormal Papanicolaou smear of vagina and vaginal HPV|Other abnormal Papanicolaou smear of vagina and vaginal HPV
C0476431|T033|AB|795.2|ICD9CM|Abn chromosomal analysis|Abn chromosomal analysis
C0476431|T033|PT|795.2|ICD9CM|Nonspecific abnormal findings on chromosomal analysis|Nonspecific abnormal findings on chromosomal analysis
C0159125|T033|HT|795.3|ICD9CM|Nonspecific positive culture findings|Nonspecific positive culture findings
C1135260|T047|AB|795.31|ICD9CM|Nonsp postv find-anthrax|Nonsp postv find-anthrax
C1135260|T047|PT|795.31|ICD9CM|Nonspecific positive findings for anthrax|Nonspecific positive findings for anthrax
C1135261|T047|AB|795.39|ICD9CM|Nonsp positive cult NEC|Nonsp positive cult NEC
C1135261|T047|PT|795.39|ICD9CM|Other nonspecific positive culture findings|Other nonspecific positive culture findings
C0159126|T033|AB|795.4|ICD9CM|Abn histologic find NEC|Abn histologic find NEC
C0159126|T033|PT|795.4|ICD9CM|Other nonspecific abnormal histological findings|Other nonspecific abnormal histological findings
C3161127|T033|HT|795.5|ICD9CM|Nonspecific reaction to tuberculin skin test without active tuberculosis|Nonspecific reaction to tuberculin skin test without active tuberculosis
C3161127|T033|AB|795.51|ICD9CM|Nonsp rea skn test wo tb|Nonsp rea skn test wo tb
C3161127|T033|PT|795.51|ICD9CM|Nonspecific reaction to tuberculin skin test without active tuberculosis|Nonspecific reaction to tuberculin skin test without active tuberculosis
C3161128|T033|AB|795.52|ICD9CM|Nonsp rea gma interferon|Nonsp rea gma interferon
C0159128|T033|AB|795.6|ICD9CM|False pos sero test-syph|False pos sero test-syph
C0159128|T033|PT|795.6|ICD9CM|False positive serological test for syphilis|False positive serological test for syphilis
C0375580|T033|HT|795.7|ICD9CM|Other nonspecific immunological findings|Other nonspecific immunological findings
C0375580|T033|AB|795.79|ICD9CM|Oth unspcf nspf imun fnd|Oth unspcf nspf imun fnd
C0375580|T033|PT|795.79|ICD9CM|Other and unspecified nonspecific immunological findings|Other and unspecified nonspecific immunological findings
C1719651|T033|HT|795.8|ICD9CM|Abnormal tumor markers|Abnormal tumor markers
C1719649|T033|AB|795.81|ICD9CM|Elev ca-embryoic antigen|Elev ca-embryoic antigen
C1719649|T033|PT|795.81|ICD9CM|Elevated carcinoembryonic antigen [CEA]|Elevated carcinoembryonic antigen [CEA]
C0238875|T033|AB|795.82|ICD9CM|Elev ca antigen 125|Elev ca antigen 125
C0238875|T033|PT|795.82|ICD9CM|Elevated cancer antigen 125 [CA 125]|Elevated cancer antigen 125 [CA 125]
C1719650|T033|AB|795.89|ICD9CM|Abnorml tumor marker NEC|Abnorml tumor marker NEC
C1719650|T033|PT|795.89|ICD9CM|Other abnormal tumor markers|Other abnormal tumor markers
C0159131|T033|HT|796|ICD9CM|Other nonspecific abnormal findings|Other nonspecific abnormal findings
C0159132|T033|AB|796.0|ICD9CM|Abn toxicologic finding|Abn toxicologic finding
C0159132|T033|PT|796.0|ICD9CM|Nonspecific abnormal toxicological findings|Nonspecific abnormal toxicological findings
C0034933|T033|AB|796.1|ICD9CM|Abnormal reflex|Abnormal reflex
C0034933|T033|PT|796.1|ICD9CM|Abnormal reflex|Abnormal reflex
C0392682|T033|AB|796.2|ICD9CM|Elev bl pres w/o hypertn|Elev bl pres w/o hypertn
C0392682|T033|PT|796.2|ICD9CM|Elevated blood pressure reading without diagnosis of hypertension|Elevated blood pressure reading without diagnosis of hypertension
C0476454|T033|AB|796.3|ICD9CM|Low blood press reading|Low blood press reading
C0476454|T033|PT|796.3|ICD9CM|Nonspecific low blood pressure reading|Nonspecific low blood pressure reading
C0159135|T033|AB|796.4|ICD9CM|Abn clinical finding NEC|Abn clinical finding NEC
C0159135|T033|PT|796.4|ICD9CM|Other abnormal clinical findings|Other abnormal clinical findings
C0490012|T033|AB|796.5|ICD9CM|Abn find antenatl screen|Abn find antenatl screen
C0490012|T033|PT|796.5|ICD9CM|Abnormal finding on antenatal screening|Abnormal finding on antenatal screening
C1455903|T033|AB|796.6|ICD9CM|Abnorm neonate screening|Abnorm neonate screening
C1455903|T033|PT|796.6|ICD9CM|Abnormal findings on neonatal screening|Abnormal findings on neonatal screening
C2349713|T033|HT|796.7|ICD9CM|Abnormal cytologic smear of anus and anal HPV|Abnormal cytologic smear of anus and anal HPV
C2349699|T033|AB|796.70|ICD9CM|Abn gland pap smear anus|Abn gland pap smear anus
C2349699|T033|PT|796.70|ICD9CM|Abnormal glandular Papanicolaou smear of anus|Abnormal glandular Papanicolaou smear of anus
C2349701|T033|AB|796.71|ICD9CM|Pap smear anus w ASC-US|Pap smear anus w ASC-US
C2349701|T033|PT|796.71|ICD9CM|Papanicolaou smear of anus with atypical squamous cells of undetermined significance (ASC-US)|Papanicolaou smear of anus with atypical squamous cells of undetermined significance (ASC-US)
C2349702|T033|AB|796.72|ICD9CM|Pap smear anus w ASC-H|Pap smear anus w ASC-H
C2349703|T033|AB|796.73|ICD9CM|Pap smear anus w LGSIL|Pap smear anus w LGSIL
C2349703|T033|PT|796.73|ICD9CM|Papanicolaou smear of anus with low grade squamous intraepithelial lesion (LGSIL)|Papanicolaou smear of anus with low grade squamous intraepithelial lesion (LGSIL)
C2349704|T033|AB|796.74|ICD9CM|Pap smear anus w HGSIL|Pap smear anus w HGSIL
C2349704|T033|PT|796.74|ICD9CM|Papanicolaou smear of anus with high grade squamous intraepithelial lesion (HGSIL)|Papanicolaou smear of anus with high grade squamous intraepithelial lesion (HGSIL)
C2349705|T033|AB|796.75|ICD9CM|Anal hi risk HPV-DNA pos|Anal hi risk HPV-DNA pos
C2349705|T033|PT|796.75|ICD9CM|Anal high risk human papillomavirus (HPV) DNA test positive|Anal high risk human papillomavirus (HPV) DNA test positive
C2349706|T033|AB|796.76|ICD9CM|Pap smr anus-cytol malig|Pap smr anus-cytol malig
C2349706|T033|PT|796.76|ICD9CM|Papanicolaou smear of anus with cytologic evidence of malignancy|Papanicolaou smear of anus with cytologic evidence of malignancy
C2349707|T033|AB|796.77|ICD9CM|Sat anal smr-no trnsfrm|Sat anal smr-no trnsfrm
C2349707|T033|PT|796.77|ICD9CM|Satisfactory anal smear but lacking transformation zone|Satisfactory anal smear but lacking transformation zone
C2349708|T033|AB|796.78|ICD9CM|Anal cytolgy smr unsatis|Anal cytolgy smr unsatis
C2349708|T033|PT|796.78|ICD9CM|Unsatisfactory anal cytology smear|Unsatisfactory anal cytology smear
C2349710|T033|AB|796.79|ICD9CM|Oth abn Pap smr anus/HPV|Oth abn Pap smr anus/HPV
C2349710|T033|PT|796.79|ICD9CM|Other abnormal Papanicolaou smear of anus and anal HPV|Other abnormal Papanicolaou smear of anus and anal HPV
C0159131|T033|AB|796.9|ICD9CM|Abnormal findings NEC|Abnormal findings NEC
C0159131|T033|PT|796.9|ICD9CM|Other nonspecific abnormal findings|Other nonspecific abnormal findings
C0036654|T048|AB|797|ICD9CM|Senility w/o psychosis|Senility w/o psychosis
C0036654|T048|PT|797|ICD9CM|Senility without mention of psychosis|Senility without mention of psychosis
C0362047|T033|HT|797-799.99|ICD9CM|ILL-DEFINED AND UNKNOWN CAUSES OF MORBIDITY AND MORTALITY|ILL-DEFINED AND UNKNOWN CAUSES OF MORBIDITY AND MORTALITY
C0520806|T033|HT|798|ICD9CM|Sudden death, cause unknown|Sudden death, cause unknown
C0038644|T047|AB|798.0|ICD9CM|Sudden infant death synd|Sudden infant death synd
C0038644|T047|PT|798.0|ICD9CM|Sudden infant death syndrome|Sudden infant death syndrome
C0021614|T046|AB|798.1|ICD9CM|Instantaneous death|Instantaneous death
C0021614|T046|PT|798.1|ICD9CM|Instantaneous death|Instantaneous death
C0277590|T033|PT|798.2|ICD9CM|Death occurring in less than 24 hours from onset of symptoms, not otherwise explained|Death occurring in less than 24 hours from onset of symptoms, not otherwise explained
C0277590|T033|AB|798.2|ICD9CM|Death within 24 hr sympt|Death within 24 hr sympt
C0152229|T033|AB|798.9|ICD9CM|Unattended death|Unattended death
C0152229|T033|PT|798.9|ICD9CM|Unattended death|Unattended death
C0159138|T033|HT|799|ICD9CM|Other ill-defined and unknown causes of morbidity and mortality|Other ill-defined and unknown causes of morbidity and mortality
C1561822|T046|HT|799.0|ICD9CM|Asphyxia and hypoxemia|Asphyxia and hypoxemia
C0004044|T046|AB|799.01|ICD9CM|Asphyxia|Asphyxia
C0004044|T046|PT|799.01|ICD9CM|Asphyxia|Asphyxia
C0700292|T033|PT|799.02|ICD9CM|Hypoxemia|Hypoxemia
C0700292|T033|AB|799.02|ICD9CM|Hypoxemia|Hypoxemia
C0162297|T046|AB|799.1|ICD9CM|Respiratory arrest|Respiratory arrest
C0162297|T046|PT|799.1|ICD9CM|Respiratory arrest|Respiratory arrest
C0495691|T184|HT|799.2|ICD9CM|Signs and symptoms involving emotional state|Signs and symptoms involving emotional state
C0027769|T184|AB|799.21|ICD9CM|Nervousness|Nervousness
C0027769|T184|PT|799.21|ICD9CM|Nervousness|Nervousness
C0022107|T033|AB|799.22|ICD9CM|Irritability|Irritability
C0022107|T033|PT|799.22|ICD9CM|Irritability|Irritability
C0564567|T048|AB|799.23|ICD9CM|Impulsiveness|Impulsiveness
C0564567|T048|PT|799.23|ICD9CM|Impulsiveness|Impulsiveness
C0085633|T048|AB|799.24|ICD9CM|Emotional lability|Emotional lability
C0085633|T048|PT|799.24|ICD9CM|Emotional lability|Emotional lability
C0476478|T184|AB|799.25|ICD9CM|Demoralization & apathy|Demoralization & apathy
C0476478|T184|PT|799.25|ICD9CM|Demoralization and apathy|Demoralization and apathy
C0478140|T184|AB|799.29|ICD9CM|Emotional state sym NEC|Emotional state sym NEC
C0478140|T184|PT|799.29|ICD9CM|Other signs and symptoms involving emotional state|Other signs and symptoms involving emotional state
C3714552|T184|AB|799.3|ICD9CM|Debility NOS|Debility NOS
C3714552|T184|PT|799.3|ICD9CM|Debility, unspecified|Debility, unspecified
C0006625|T184|AB|799.4|ICD9CM|Cachexia|Cachexia
C0006625|T184|PT|799.4|ICD9CM|Cachexia|Cachexia
C2921135|T184|HT|799.5|ICD9CM|Signs and symptoms involving cognition|Signs and symptoms involving cognition
C2921136|T184|PT|799.51|ICD9CM|Attention or concentration deficit|Attention or concentration deficit
C2921136|T184|AB|799.51|ICD9CM|Attn/concentrate deficit|Attn/concentrate deficit
C2921137|T184|AB|799.52|ICD9CM|Cog communicate deficit|Cog communicate deficit
C2921137|T184|PT|799.52|ICD9CM|Cognitive communication deficit|Cognitive communication deficit
C2921138|T184|AB|799.53|ICD9CM|Visuospatial deficit|Visuospatial deficit
C2921138|T184|PT|799.53|ICD9CM|Visuospatial deficit|Visuospatial deficit
C2921139|T033|PT|799.54|ICD9CM|Psychomotor deficit|Psychomotor deficit
C2921139|T033|AB|799.54|ICD9CM|Psychomotor deficit|Psychomotor deficit
C2921140|T184|PT|799.55|ICD9CM|Frontal lobe and executive function deficit|Frontal lobe and executive function deficit
C2921140|T184|AB|799.55|ICD9CM|Frontal lobe deficit|Frontal lobe deficit
C2921141|T184|AB|799.59|ICD9CM|Cognition sign/sympt NEC|Cognition sign/sympt NEC
C2921141|T184|PT|799.59|ICD9CM|Other signs and symptoms involving cognition|Other signs and symptoms involving cognition
C0277538|T046|HT|799.8|ICD9CM|Other ill-defined conditions|Other ill-defined conditions
C0011124|T033|AB|799.81|ICD9CM|Decreased libido|Decreased libido
C0011124|T033|PT|799.81|ICD9CM|Decreased libido|Decreased libido
C2712370|T047|AB|799.82|ICD9CM|Appar life threat-infant|Appar life threat-infant
C2712370|T047|PT|799.82|ICD9CM|Apparent life threatening event in infant|Apparent life threatening event in infant
C0277538|T046|AB|799.89|ICD9CM|Ill-define condition NEC|Ill-define condition NEC
C0277538|T046|PT|799.89|ICD9CM|Other ill-defined conditions|Other ill-defined conditions
C0476465|T033|PT|799.9|ICD9CM|Other unknown and unspecified cause of morbidity and mortality|Other unknown and unspecified cause of morbidity and mortality
C0476465|T033|AB|799.9|ICD9CM|Unkn cause morb/mort NEC|Unkn cause morb/mort NEC
C0159139|T037|HT|800|ICD9CM|Fracture of vault of skull|Fracture of vault of skull
C0037304|T037|HT|800-804.99|ICD9CM|FRACTURE OF SKULL|FRACTURE OF SKULL
C0016658|T037|HT|800-829.99|ICD9CM|FRACTURES|FRACTURES
C0178314|T037|HT|800-999.99|ICD9CM|INJURY AND POISONING|INJURY AND POISONING
C0159140|T037|HT|800.0|ICD9CM|Closed fracture of vault of skull without mention of intracranial injury|Closed fracture of vault of skull without mention of intracranial injury
C0159141|T037|AB|800.00|ICD9CM|Closed skull vault fx|Closed skull vault fx
C0159142|T037|AB|800.01|ICD9CM|Cl skull vlt fx w/o coma|Cl skull vlt fx w/o coma
C0159143|T037|AB|800.02|ICD9CM|Cl skull vlt fx-brf coma|Cl skull vlt fx-brf coma
C0159144|T037|AB|800.03|ICD9CM|Cl skull vlt fx-mod coma|Cl skull vlt fx-mod coma
C0159145|T037|AB|800.04|ICD9CM|Cl skl vlt fx-proln coma|Cl skl vlt fx-proln coma
C0159146|T037|AB|800.05|ICD9CM|Cl skul vlt fx-deep coma|Cl skul vlt fx-deep coma
C0159147|T037|AB|800.06|ICD9CM|Cl skull vlt fx-coma NOS|Cl skull vlt fx-coma NOS
C0159148|T037|AB|800.09|ICD9CM|Cl skl vlt fx-concus NOS|Cl skl vlt fx-concus NOS
C0159149|T037|HT|800.1|ICD9CM|Closed fracture of vault of skull with cerebral laceration and contusion|Closed fracture of vault of skull with cerebral laceration and contusion
C0159150|T037|AB|800.10|ICD9CM|Cl skl vlt fx/cerebr lac|Cl skl vlt fx/cerebr lac
C0159151|T037|AB|800.11|ICD9CM|Cl skull vlt fx w/o coma|Cl skull vlt fx w/o coma
C0159152|T037|AB|800.12|ICD9CM|Cl skull vlt fx-brf coma|Cl skull vlt fx-brf coma
C0159153|T037|AB|800.13|ICD9CM|Cl skull vlt fx-mod coma|Cl skull vlt fx-mod coma
C0159154|T037|AB|800.14|ICD9CM|Cl skl vlt fx-proln coma|Cl skl vlt fx-proln coma
C0159155|T037|AB|800.15|ICD9CM|Cl skul vlt fx-deep coma|Cl skul vlt fx-deep coma
C0159156|T037|AB|800.16|ICD9CM|Cl skull vlt fx-coma NOS|Cl skull vlt fx-coma NOS
C0375581|T037|AB|800.19|ICD9CM|Cl skl vlt fx-concus NOS|Cl skl vlt fx-concus NOS
C0159158|T037|HT|800.2|ICD9CM|Closed fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage|Closed fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage
C0159159|T037|AB|800.20|ICD9CM|Cl skl vlt fx/mening hem|Cl skl vlt fx/mening hem
C0159160|T037|AB|800.21|ICD9CM|Cl skull vlt fx w/o coma|Cl skull vlt fx w/o coma
C0159161|T037|AB|800.22|ICD9CM|Cl skull vlt fx-brf coma|Cl skull vlt fx-brf coma
C0159162|T037|AB|800.23|ICD9CM|Cl skull vlt fx-mod coma|Cl skull vlt fx-mod coma
C0159163|T037|AB|800.24|ICD9CM|Cl skl vlt fx-proln coma|Cl skl vlt fx-proln coma
C0159164|T037|AB|800.25|ICD9CM|Cl skul vlt fx-deep coma|Cl skul vlt fx-deep coma
C0159165|T037|AB|800.26|ICD9CM|Cl skull vlt fx-coma NOS|Cl skull vlt fx-coma NOS
C0375582|T037|AB|800.29|ICD9CM|Cl skl vlt fx-concus NOS|Cl skl vlt fx-concus NOS
C0159167|T037|HT|800.3|ICD9CM|Closed fracture of vault of skull with other and unspecified intracranial hemorrhage|Closed fracture of vault of skull with other and unspecified intracranial hemorrhage
C0159168|T037|AB|800.30|ICD9CM|Cl skull vlt fx/hem NEC|Cl skull vlt fx/hem NEC
C0159169|T037|AB|800.31|ICD9CM|Cl skull vlt fx w/o coma|Cl skull vlt fx w/o coma
C0159170|T037|AB|800.32|ICD9CM|Cl skull vlt fx-brf coma|Cl skull vlt fx-brf coma
C0159171|T037|AB|800.33|ICD9CM|Cl skull vlt fx-mod coma|Cl skull vlt fx-mod coma
C0159172|T037|AB|800.34|ICD9CM|Cl skl vlt fx-proln coma|Cl skl vlt fx-proln coma
C0159173|T037|AB|800.35|ICD9CM|Cl skul vlt fx-deep coma|Cl skul vlt fx-deep coma
C0159174|T037|AB|800.36|ICD9CM|Cl skull vlt fx-coma NOS|Cl skull vlt fx-coma NOS
C0375583|T037|AB|800.39|ICD9CM|Cl skl vlt fx-concus NOS|Cl skl vlt fx-concus NOS
C0159176|T037|HT|800.4|ICD9CM|Closed fracture of vault of skull with intracranial injury of other and unspecified nature|Closed fracture of vault of skull with intracranial injury of other and unspecified nature
C0159177|T037|AB|800.40|ICD9CM|Cl skl vlt fx/br inj NEC|Cl skl vlt fx/br inj NEC
C0159178|T037|AB|800.41|ICD9CM|Cl skull vlt fx w/o coma|Cl skull vlt fx w/o coma
C0159179|T037|AB|800.42|ICD9CM|Cl skull vlt fx-brf coma|Cl skull vlt fx-brf coma
C0159180|T037|AB|800.43|ICD9CM|Cl skull vlt fx-mod coma|Cl skull vlt fx-mod coma
C0159181|T037|AB|800.44|ICD9CM|Cl skl vlt fx-proln coma|Cl skl vlt fx-proln coma
C0159182|T037|AB|800.45|ICD9CM|Cl skul vlt fx-deep coma|Cl skul vlt fx-deep coma
C0159183|T037|AB|800.46|ICD9CM|Cl skull vlt fx-coma NOS|Cl skull vlt fx-coma NOS
C0159184|T037|AB|800.49|ICD9CM|Cl skl vlt fx-concus NOS|Cl skl vlt fx-concus NOS
C0159185|T037|HT|800.5|ICD9CM|Open fracture of vault of skull without mention of intracranial injury|Open fracture of vault of skull without mention of intracranial injury
C0159186|T037|AB|800.50|ICD9CM|Opn skull vault fracture|Opn skull vault fracture
C0159187|T037|AB|800.51|ICD9CM|Opn skul vlt fx w/o coma|Opn skul vlt fx w/o coma
C0159188|T037|AB|800.52|ICD9CM|Opn skul vlt fx-brf coma|Opn skul vlt fx-brf coma
C0159189|T037|AB|800.53|ICD9CM|Opn skul vlt fx-mod coma|Opn skul vlt fx-mod coma
C0159190|T037|AB|800.54|ICD9CM|Opn skl vlt fx-proln com|Opn skl vlt fx-proln com
C0159191|T037|AB|800.55|ICD9CM|Opn skl vlt fx-deep coma|Opn skl vlt fx-deep coma
C0159192|T037|AB|800.56|ICD9CM|Opn skul vlt fx-coma NOS|Opn skul vlt fx-coma NOS
C0159193|T037|AB|800.59|ICD9CM|Op skl vlt fx-concus NOS|Op skl vlt fx-concus NOS
C0159193|T037|PT|800.59|ICD9CM|Open fracture of vault of skull without mention of intracranial injury, with concussion, unspecified|Open fracture of vault of skull without mention of intracranial injury, with concussion, unspecified
C0159194|T037|HT|800.6|ICD9CM|Open fracture of vault of skull with cerebral laceration and contusion|Open fracture of vault of skull with cerebral laceration and contusion
C0159195|T037|AB|800.60|ICD9CM|Opn skl vlt fx/cereb lac|Opn skl vlt fx/cereb lac
C0159196|T037|AB|800.61|ICD9CM|Opn skul vlt fx w/o coma|Opn skul vlt fx w/o coma
C0159197|T037|AB|800.62|ICD9CM|Opn skul vlt fx-brf coma|Opn skul vlt fx-brf coma
C0159198|T037|AB|800.63|ICD9CM|Opn skul vlt fx-mod coma|Opn skul vlt fx-mod coma
C0159199|T037|AB|800.64|ICD9CM|Opn skl vlt fx-proln com|Opn skl vlt fx-proln com
C0159200|T037|AB|800.65|ICD9CM|Opn skl vlt fx-deep coma|Opn skl vlt fx-deep coma
C0159201|T037|AB|800.66|ICD9CM|Opn skul vlt fx-coma NOS|Opn skul vlt fx-coma NOS
C0375585|T037|AB|800.69|ICD9CM|Op skl vlt fx-concus NOS|Op skl vlt fx-concus NOS
C0375585|T037|PT|800.69|ICD9CM|Open fracture of vault of skull with cerebral laceration and contusion, with concussion, unspecified|Open fracture of vault of skull with cerebral laceration and contusion, with concussion, unspecified
C0159203|T037|HT|800.7|ICD9CM|Open fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage|Open fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage
C0159204|T037|AB|800.70|ICD9CM|Opn skl vlt fx/menin hem|Opn skl vlt fx/menin hem
C0159205|T037|AB|800.71|ICD9CM|Opn skul vlt fx w/o coma|Opn skul vlt fx w/o coma
C0159206|T037|AB|800.72|ICD9CM|Opn skul vlt fx-brf coma|Opn skul vlt fx-brf coma
C0159207|T037|AB|800.73|ICD9CM|Opn skul vlt fx-mod coma|Opn skul vlt fx-mod coma
C0159208|T037|AB|800.74|ICD9CM|Opn skl vlt fx-proln com|Opn skl vlt fx-proln com
C0159209|T037|AB|800.75|ICD9CM|Opn skl vlt fx-deep coma|Opn skl vlt fx-deep coma
C0159210|T037|AB|800.76|ICD9CM|Opn skul vlt fx-coma NOS|Opn skul vlt fx-coma NOS
C0375586|T037|AB|800.79|ICD9CM|Op skl vlt fx-concus NOS|Op skl vlt fx-concus NOS
C0159212|T037|HT|800.8|ICD9CM|Open fracture of vault of skull with other and unspecified intracranial hemorrhage|Open fracture of vault of skull with other and unspecified intracranial hemorrhage
C0159213|T037|AB|800.80|ICD9CM|Opn skull vlt fx/hem NEC|Opn skull vlt fx/hem NEC
C0159214|T037|AB|800.81|ICD9CM|Opn skul vlt fx w/o coma|Opn skul vlt fx w/o coma
C0159215|T037|AB|800.82|ICD9CM|Opn skul vlt fx-brf coma|Opn skul vlt fx-brf coma
C0159216|T037|AB|800.83|ICD9CM|Opn skul vlt fx-mod coma|Opn skul vlt fx-mod coma
C0159217|T037|AB|800.84|ICD9CM|Opn skl vlt fx-proln com|Opn skl vlt fx-proln com
C0159218|T037|AB|800.85|ICD9CM|Opn skl vlt fx-deep coma|Opn skl vlt fx-deep coma
C0159219|T037|AB|800.86|ICD9CM|Opn skul vlt fx-coma NOS|Opn skul vlt fx-coma NOS
C0375587|T037|AB|800.89|ICD9CM|Op skl vlt fx-concus NOS|Op skl vlt fx-concus NOS
C0159221|T037|HT|800.9|ICD9CM|Open fracture of vault of skull with intracranial injury of other and unspecified nature|Open fracture of vault of skull with intracranial injury of other and unspecified nature
C0159222|T037|AB|800.90|ICD9CM|Op skl vlt fx/br inj NEC|Op skl vlt fx/br inj NEC
C0159223|T037|AB|800.91|ICD9CM|Opn skul vlt fx w/o coma|Opn skul vlt fx w/o coma
C0159224|T037|AB|800.92|ICD9CM|Opn skul vlt fx-brf coma|Opn skul vlt fx-brf coma
C0159225|T037|AB|800.93|ICD9CM|Opn skul vlt fx-mod coma|Opn skul vlt fx-mod coma
C0159226|T037|AB|800.94|ICD9CM|Opn skl vlt fx-proln com|Opn skl vlt fx-proln com
C0159227|T037|AB|800.95|ICD9CM|Op skul vlt fx-deep coma|Op skul vlt fx-deep coma
C0159228|T037|AB|800.96|ICD9CM|Opn skul vlt fx-coma NOS|Opn skul vlt fx-coma NOS
C0159229|T037|AB|800.99|ICD9CM|Op skl vlt fx-concus NOS|Op skl vlt fx-concus NOS
C0748830|T037|HT|801|ICD9CM|Fracture of base of skull|Fracture of base of skull
C0435271|T037|HT|801.0|ICD9CM|Closed fracture of base of skull without mention of intracranial injury|Closed fracture of base of skull without mention of intracranial injury
C0159232|T037|AB|801.00|ICD9CM|Clos skull base fracture|Clos skull base fracture
C0159233|T037|AB|801.01|ICD9CM|Cl skul base fx w/o coma|Cl skul base fx w/o coma
C0159234|T037|AB|801.02|ICD9CM|Cl skul base fx-brf coma|Cl skul base fx-brf coma
C0159235|T037|AB|801.03|ICD9CM|Cl skul base fx-mod coma|Cl skul base fx-mod coma
C0159236|T037|AB|801.04|ICD9CM|Cl skl base fx-prol coma|Cl skl base fx-prol coma
C0159237|T037|AB|801.05|ICD9CM|Cl skl base fx-deep coma|Cl skl base fx-deep coma
C0159238|T037|AB|801.06|ICD9CM|Cl skul base fx-coma NOS|Cl skul base fx-coma NOS
C0159239|T037|AB|801.09|ICD9CM|Cl skull base fx-concuss|Cl skull base fx-concuss
C0159240|T037|HT|801.1|ICD9CM|Closed fracture of base of skull with cerebral laceration and contusion|Closed fracture of base of skull with cerebral laceration and contusion
C0159241|T037|AB|801.10|ICD9CM|Cl skl base fx/cereb lac|Cl skl base fx/cereb lac
C0159242|T037|AB|801.11|ICD9CM|Cl skul base fx w/o coma|Cl skul base fx w/o coma
C0159243|T037|AB|801.12|ICD9CM|Cl skul base fx-brf coma|Cl skul base fx-brf coma
C0159244|T037|AB|801.13|ICD9CM|Cl skul base fx-mod coma|Cl skul base fx-mod coma
C0159245|T037|AB|801.14|ICD9CM|Cl skl base fx-prol coma|Cl skl base fx-prol coma
C0159246|T037|AB|801.15|ICD9CM|Cl skl base fx-deep coma|Cl skl base fx-deep coma
C0159247|T037|AB|801.16|ICD9CM|Cl skul base fx-coma NOS|Cl skul base fx-coma NOS
C0375589|T037|AB|801.19|ICD9CM|Cl skull base fx-concuss|Cl skull base fx-concuss
C0159249|T037|HT|801.2|ICD9CM|Closed fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage|Closed fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage
C0159250|T037|AB|801.20|ICD9CM|Cl skl base fx/menin hem|Cl skl base fx/menin hem
C0159251|T037|AB|801.21|ICD9CM|Cl skul base fx w/o coma|Cl skul base fx w/o coma
C0159252|T037|AB|801.22|ICD9CM|Cl skul base fx/brf coma|Cl skul base fx/brf coma
C0159253|T037|AB|801.23|ICD9CM|Cl skul base fx-mod coma|Cl skul base fx-mod coma
C0159254|T037|AB|801.24|ICD9CM|Cl skl base fx-prol coma|Cl skl base fx-prol coma
C0159255|T037|AB|801.25|ICD9CM|Cl skl base fx-deep coma|Cl skl base fx-deep coma
C0159256|T037|AB|801.26|ICD9CM|Cl skul base fx-coma NOS|Cl skul base fx-coma NOS
C0375590|T037|AB|801.29|ICD9CM|Cl skull base fx-concuss|Cl skull base fx-concuss
C0159258|T037|HT|801.3|ICD9CM|Closed fracture of base of skull with other and unspecified intracranial hemorrhage|Closed fracture of base of skull with other and unspecified intracranial hemorrhage
C0159259|T037|AB|801.30|ICD9CM|Cl skull base fx/hem NEC|Cl skull base fx/hem NEC
C0159260|T037|AB|801.31|ICD9CM|Cl skul base fx w/o coma|Cl skul base fx w/o coma
C0159261|T037|AB|801.32|ICD9CM|Cl skul base fx-brf coma|Cl skul base fx-brf coma
C0159262|T037|AB|801.33|ICD9CM|Cl skul base fx-mod coma|Cl skul base fx-mod coma
C0159263|T037|AB|801.34|ICD9CM|Cl skl base fx-prol coma|Cl skl base fx-prol coma
C0159264|T037|AB|801.35|ICD9CM|Cl skl base fx-deep coma|Cl skl base fx-deep coma
C0159265|T037|AB|801.36|ICD9CM|Cl skul base fx-coma NOS|Cl skul base fx-coma NOS
C0375591|T037|AB|801.39|ICD9CM|Cl skull base fx-concuss|Cl skull base fx-concuss
C0159267|T037|HT|801.4|ICD9CM|Closed fracture of base of skull with intracranial injury of other and unspecified nature|Closed fracture of base of skull with intracranial injury of other and unspecified nature
C0159268|T037|AB|801.40|ICD9CM|Cl sk base fx/br inj NEC|Cl sk base fx/br inj NEC
C0159269|T037|AB|801.41|ICD9CM|Cl skul base fx w/o coma|Cl skul base fx w/o coma
C0159270|T037|AB|801.42|ICD9CM|Cl skul base fx-brf coma|Cl skul base fx-brf coma
C0159271|T037|AB|801.43|ICD9CM|Cl skul base fx-mod coma|Cl skul base fx-mod coma
C0159272|T037|AB|801.44|ICD9CM|Cl skl base fx-prol coma|Cl skl base fx-prol coma
C0159273|T037|AB|801.45|ICD9CM|Cl skl base fx-deep coma|Cl skl base fx-deep coma
C0159274|T037|AB|801.46|ICD9CM|Cl skul base fx-coma NOS|Cl skul base fx-coma NOS
C0159275|T037|AB|801.49|ICD9CM|Cl skull base fx-concuss|Cl skull base fx-concuss
C0159276|T037|HT|801.5|ICD9CM|Open fracture of base of skull without mention of intracranial injury|Open fracture of base of skull without mention of intracranial injury
C0159277|T037|AB|801.50|ICD9CM|Open skull base fracture|Open skull base fracture
C0159278|T037|PT|801.51|ICD9CM|Open fracture of base of skull without mention of intracranial injury, with no loss of consciousness|Open fracture of base of skull without mention of intracranial injury, with no loss of consciousness
C0159278|T037|AB|801.51|ICD9CM|Opn skl base fx w/o coma|Opn skl base fx w/o coma
C0159279|T037|AB|801.52|ICD9CM|Opn skl base fx-brf coma|Opn skl base fx-brf coma
C0159280|T037|AB|801.53|ICD9CM|Opn skl base fx-mod coma|Opn skl base fx-mod coma
C0159281|T037|AB|801.54|ICD9CM|Op skl base fx-prol coma|Op skl base fx-prol coma
C0159282|T037|AB|801.55|ICD9CM|Op skl base fx-deep coma|Op skl base fx-deep coma
C0159283|T037|AB|801.56|ICD9CM|Opn skl base fx-coma NOS|Opn skl base fx-coma NOS
C0159284|T037|PT|801.59|ICD9CM|Open fracture of base of skull without mention of intracranial injury, with concussion, unspecified|Open fracture of base of skull without mention of intracranial injury, with concussion, unspecified
C0159284|T037|AB|801.59|ICD9CM|Opn skul base fx-concuss|Opn skul base fx-concuss
C0159285|T037|HT|801.6|ICD9CM|Open fracture of base of skull with cerebral laceration and contusion|Open fracture of base of skull with cerebral laceration and contusion
C0159286|T037|AB|801.60|ICD9CM|Op skl base fx/cereb lac|Op skl base fx/cereb lac
C0159287|T037|PT|801.61|ICD9CM|Open fracture of base of skull with cerebral laceration and contusion, with no loss of consciousness|Open fracture of base of skull with cerebral laceration and contusion, with no loss of consciousness
C0159287|T037|AB|801.61|ICD9CM|Opn skl base fx w/o coma|Opn skl base fx w/o coma
C0159288|T037|AB|801.62|ICD9CM|Opn skl base fx-brf coma|Opn skl base fx-brf coma
C0159289|T037|AB|801.63|ICD9CM|Opn skl base fx-mod coma|Opn skl base fx-mod coma
C0159290|T037|AB|801.64|ICD9CM|Op skl base fx-prol coma|Op skl base fx-prol coma
C0159291|T037|AB|801.65|ICD9CM|Op skl base fx-deep coma|Op skl base fx-deep coma
C0159292|T037|AB|801.66|ICD9CM|Opn skl base fx-coma NOS|Opn skl base fx-coma NOS
C0375593|T037|PT|801.69|ICD9CM|Open fracture of base of skull with cerebral laceration and contusion, with concussion, unspecified|Open fracture of base of skull with cerebral laceration and contusion, with concussion, unspecified
C0375593|T037|AB|801.69|ICD9CM|Opn skul base fx-concuss|Opn skul base fx-concuss
C0159294|T037|HT|801.7|ICD9CM|Open fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage|Open fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage
C0159295|T037|AB|801.70|ICD9CM|Op skl base fx/menin hem|Op skl base fx/menin hem
C0159296|T037|AB|801.71|ICD9CM|Opn skl base fx w/o coma|Opn skl base fx w/o coma
C0159297|T037|AB|801.72|ICD9CM|Opn skl base fx-brf coma|Opn skl base fx-brf coma
C0159298|T037|AB|801.73|ICD9CM|Opn skl base fx-mod coma|Opn skl base fx-mod coma
C0159299|T037|AB|801.74|ICD9CM|Op skl base fx-prol coma|Op skl base fx-prol coma
C0159300|T037|AB|801.75|ICD9CM|Op skl base fx-deep coma|Op skl base fx-deep coma
C0159301|T037|AB|801.76|ICD9CM|Opn skl base fx-coma NOS|Opn skl base fx-coma NOS
C0375594|T037|AB|801.79|ICD9CM|Opn skul base fx-concuss|Opn skul base fx-concuss
C0159303|T037|HT|801.8|ICD9CM|Open fracture of base of skull with other and unspecified intracranial hemorrhage|Open fracture of base of skull with other and unspecified intracranial hemorrhage
C0159304|T037|AB|801.80|ICD9CM|Opn skul base fx/hem NEC|Opn skul base fx/hem NEC
C0159305|T037|AB|801.81|ICD9CM|Opn skl base fx w/o coma|Opn skl base fx w/o coma
C0159306|T037|AB|801.82|ICD9CM|Opn skl base fx-brf coma|Opn skl base fx-brf coma
C0159307|T037|AB|801.83|ICD9CM|Opn skl base fx-mod coma|Opn skl base fx-mod coma
C0159308|T037|AB|801.84|ICD9CM|Op skl base fx-prol coma|Op skl base fx-prol coma
C0159309|T037|AB|801.85|ICD9CM|Op skl base fx-deep coma|Op skl base fx-deep coma
C0159310|T037|AB|801.86|ICD9CM|Opn skl base fx-coma NOS|Opn skl base fx-coma NOS
C0375595|T037|AB|801.89|ICD9CM|Opn skul base fx-concuss|Opn skul base fx-concuss
C0159312|T037|HT|801.9|ICD9CM|Open fracture of base of skull with intracranial injury of other and unspecified nature|Open fracture of base of skull with intracranial injury of other and unspecified nature
C0159313|T037|AB|801.90|ICD9CM|Op sk base fx/br inj NEC|Op sk base fx/br inj NEC
C0159314|T037|AB|801.91|ICD9CM|Op skul base fx w/o coma|Op skul base fx w/o coma
C0159315|T037|AB|801.92|ICD9CM|Opn skl base fx-brf coma|Opn skl base fx-brf coma
C0159316|T037|AB|801.93|ICD9CM|Opn skl base fx-mod coma|Opn skl base fx-mod coma
C0159317|T037|AB|801.94|ICD9CM|Op skl base fx-prol coma|Op skl base fx-prol coma
C0159318|T037|AB|801.95|ICD9CM|Op skl base fx-deep coma|Op skl base fx-deep coma
C0159319|T037|AB|801.96|ICD9CM|Opn skl base fx-coma NOS|Opn skl base fx-coma NOS
C0159320|T037|AB|801.99|ICD9CM|Opn skul base fx-concuss|Opn skul base fx-concuss
C0159321|T037|HT|802|ICD9CM|Fracture of face bones|Fracture of face bones
C0159322|T037|PT|802.0|ICD9CM|Closed fracture of nasal bones|Closed fracture of nasal bones
C0159322|T037|AB|802.0|ICD9CM|Nasal bone fx-closed|Nasal bone fx-closed
C0159323|T037|AB|802.1|ICD9CM|Nasal bone fx-open|Nasal bone fx-open
C0159323|T037|PT|802.1|ICD9CM|Open fracture of nasal bones|Open fracture of nasal bones
C0159324|T037|HT|802.2|ICD9CM|Mandible closed fracture|Mandible closed fracture
C0159324|T037|PT|802.20|ICD9CM|Closed fracture of mandible, unspecified site|Closed fracture of mandible, unspecified site
C0159324|T037|AB|802.20|ICD9CM|Mandible fx NOS-closed|Mandible fx NOS-closed
C0159325|T037|PT|802.21|ICD9CM|Closed fracture of mandible, condylar process|Closed fracture of mandible, condylar process
C0159325|T037|AB|802.21|ICD9CM|Fx condyl proc mandib-cl|Fx condyl proc mandib-cl
C0272468|T037|PT|802.22|ICD9CM|Closed fracture of mandible, subcondylar|Closed fracture of mandible, subcondylar
C0272468|T037|AB|802.22|ICD9CM|Subcondylar fx mandib-cl|Subcondylar fx mandib-cl
C0159327|T037|PT|802.23|ICD9CM|Closed fracture of mandible, coronoid process|Closed fracture of mandible, coronoid process
C0159327|T037|AB|802.23|ICD9CM|Fx coron proc mandib-cl|Fx coron proc mandib-cl
C0272469|T037|PT|802.24|ICD9CM|Closed fracture of mandible, ramus, unspecified|Closed fracture of mandible, ramus, unspecified
C0272469|T037|AB|802.24|ICD9CM|Fx ramus NOS-closed|Fx ramus NOS-closed
C0435334|T037|PT|802.25|ICD9CM|Closed fracture of mandible, angle of jaw|Closed fracture of mandible, angle of jaw
C0435334|T037|AB|802.25|ICD9CM|Fx angle of jaw-closed|Fx angle of jaw-closed
C0159330|T037|PT|802.26|ICD9CM|Closed fracture of mandible, symphysis of body|Closed fracture of mandible, symphysis of body
C0159330|T037|AB|802.26|ICD9CM|Fx symphy mandib body-cl|Fx symphy mandib body-cl
C0159331|T037|PT|802.27|ICD9CM|Closed fracture of mandible, alveolar border of body|Closed fracture of mandible, alveolar border of body
C0159331|T037|AB|802.27|ICD9CM|Fx alveolar bord mand-cl|Fx alveolar bord mand-cl
C0435335|T037|PT|802.28|ICD9CM|Closed fracture of mandible, body, other and unspecified|Closed fracture of mandible, body, other and unspecified
C0435335|T037|AB|802.28|ICD9CM|Fx mandible body NEC-cl|Fx mandible body NEC-cl
C0159333|T037|PT|802.29|ICD9CM|Closed fracture of mandible, multiple sites|Closed fracture of mandible, multiple sites
C0159333|T037|AB|802.29|ICD9CM|Mult fx mandible-closed|Mult fx mandible-closed
C0159334|T037|HT|802.3|ICD9CM|Mandible open fracture|Mandible open fracture
C0159334|T037|AB|802.30|ICD9CM|Mandible fx NOS-open|Mandible fx NOS-open
C0159334|T037|PT|802.30|ICD9CM|Open fracture of mandible, unspecified site|Open fracture of mandible, unspecified site
C0159336|T037|AB|802.31|ICD9CM|Fx condyl proc mand-open|Fx condyl proc mand-open
C0159336|T037|PT|802.31|ICD9CM|Open fracture of mandible, condylar process|Open fracture of mandible, condylar process
C0272471|T037|PT|802.32|ICD9CM|Open fracture of mandible, subcondylar|Open fracture of mandible, subcondylar
C0272471|T037|AB|802.32|ICD9CM|Subcondyl fx mandib-open|Subcondyl fx mandib-open
C0159338|T037|AB|802.33|ICD9CM|Fx coron proc mandib-opn|Fx coron proc mandib-opn
C0159338|T037|PT|802.33|ICD9CM|Open fracture of mandible, coronoid process|Open fracture of mandible, coronoid process
C0272472|T037|AB|802.34|ICD9CM|Fx ramus NOS-open|Fx ramus NOS-open
C0272472|T037|PT|802.34|ICD9CM|Open fracture of mandible, ramus, unspecified|Open fracture of mandible, ramus, unspecified
C0435337|T037|AB|802.35|ICD9CM|Fx angle of jaw-open|Fx angle of jaw-open
C0435337|T037|PT|802.35|ICD9CM|Open fracture of mandible, angle of jaw|Open fracture of mandible, angle of jaw
C0159341|T037|AB|802.36|ICD9CM|Fx symphy mandib bdy-opn|Fx symphy mandib bdy-opn
C0159341|T037|PT|802.36|ICD9CM|Open fracture of mandible, symphysis of body|Open fracture of mandible, symphysis of body
C0159342|T037|AB|802.37|ICD9CM|Fx alv bord mand bdy-opn|Fx alv bord mand bdy-opn
C0159342|T037|PT|802.37|ICD9CM|Open fracture of mandible, alveolar border of body|Open fracture of mandible, alveolar border of body
C0435338|T037|AB|802.38|ICD9CM|Fx mandible body NEC-opn|Fx mandible body NEC-opn
C0435338|T037|PT|802.38|ICD9CM|Open fracture of mandible, body, other and unspecified|Open fracture of mandible, body, other and unspecified
C0159344|T037|AB|802.39|ICD9CM|Mult fx mandible-open|Mult fx mandible-open
C0159344|T037|PT|802.39|ICD9CM|Open fracture of mandible, multiple sites|Open fracture of mandible, multiple sites
C0009045|T037|PT|802.4|ICD9CM|Closed fracture of malar and maxillary bones|Closed fracture of malar and maxillary bones
C0009045|T037|AB|802.4|ICD9CM|Fx malar/maxillary-close|Fx malar/maxillary-close
C0159345|T037|AB|802.5|ICD9CM|Fx malar/maxillary-open|Fx malar/maxillary-open
C0159345|T037|PT|802.5|ICD9CM|Open fracture of malar and maxillary bones|Open fracture of malar and maxillary bones
C0339150|T037|PT|802.6|ICD9CM|Closed fracture of orbital floor (blow-out)|Closed fracture of orbital floor (blow-out)
C0339150|T037|AB|802.6|ICD9CM|Fx orbital floor-closed|Fx orbital floor-closed
C0339151|T037|AB|802.7|ICD9CM|Fx orbital floor-open|Fx orbital floor-open
C0339151|T037|PT|802.7|ICD9CM|Open fracture of orbital floor (blow-out)|Open fracture of orbital floor (blow-out)
C0159348|T037|PT|802.8|ICD9CM|Closed fracture of other facial bones|Closed fracture of other facial bones
C0159348|T037|AB|802.8|ICD9CM|Fx facial bone NEC-close|Fx facial bone NEC-close
C0159349|T037|AB|802.9|ICD9CM|Fx facial bone NEC-open|Fx facial bone NEC-open
C0159349|T037|PT|802.9|ICD9CM|Open fracture of other facial bones|Open fracture of other facial bones
C0159350|T037|HT|803|ICD9CM|Other and unqualified skull fractures|Other and unqualified skull fractures
C0029547|T037|HT|803.0|ICD9CM|Other closed skull fracture without mention of intracranial injury|Other closed skull fracture without mention of intracranial injury
C0159351|T037|AB|803.00|ICD9CM|Close skull fracture NEC|Close skull fracture NEC
C0159352|T037|AB|803.01|ICD9CM|Cl skull fx NEC w/o coma|Cl skull fx NEC w/o coma
C0159352|T037|PT|803.01|ICD9CM|Other closed skull fracture without mention of intracranial injury, with no loss of consciousness|Other closed skull fracture without mention of intracranial injury, with no loss of consciousness
C0159353|T037|AB|803.02|ICD9CM|Cl skull fx NEC-brf coma|Cl skull fx NEC-brf coma
C0159354|T037|AB|803.03|ICD9CM|Cl skull fx NEC-mod coma|Cl skull fx NEC-mod coma
C0159355|T037|AB|803.04|ICD9CM|Cl skl fx NEC-proln coma|Cl skl fx NEC-proln coma
C0159356|T037|AB|803.05|ICD9CM|Cl skul fx NEC-deep coma|Cl skul fx NEC-deep coma
C0159357|T037|AB|803.06|ICD9CM|Cl skull fx NEC-coma NOS|Cl skull fx NEC-coma NOS
C0159358|T037|AB|803.09|ICD9CM|Cl skull fx NEC-concuss|Cl skull fx NEC-concuss
C0159358|T037|PT|803.09|ICD9CM|Other closed skull fracture without mention of intracranial injury, with concussion, unspecified|Other closed skull fracture without mention of intracranial injury, with concussion, unspecified
C0159359|T037|HT|803.1|ICD9CM|Other closed skull fracture with cerebral laceration and contusion|Other closed skull fracture with cerebral laceration and contusion
C0159360|T037|AB|803.10|ICD9CM|Cl skl fx NEC/cerebr lac|Cl skl fx NEC/cerebr lac
C0159361|T037|AB|803.11|ICD9CM|Cl skull fx NEC w/o coma|Cl skull fx NEC w/o coma
C0159361|T037|PT|803.11|ICD9CM|Other closed skull fracture with cerebral laceration and contusion, with no loss of consciousness|Other closed skull fracture with cerebral laceration and contusion, with no loss of consciousness
C0159362|T037|AB|803.12|ICD9CM|Cl skull fx NEC-brf coma|Cl skull fx NEC-brf coma
C0159363|T037|AB|803.13|ICD9CM|Cl skull fx NEC-mod coma|Cl skull fx NEC-mod coma
C0159364|T037|AB|803.14|ICD9CM|Cl skl fx NEC-proln coma|Cl skl fx NEC-proln coma
C0159365|T037|AB|803.15|ICD9CM|Cl skul fx NEC-deep coma|Cl skul fx NEC-deep coma
C0159366|T037|AB|803.16|ICD9CM|Cl skull fx NEC-coma NOS|Cl skull fx NEC-coma NOS
C0375598|T037|AB|803.19|ICD9CM|Cl skull fx NEC-concuss|Cl skull fx NEC-concuss
C0375598|T037|PT|803.19|ICD9CM|Other closed skull fracture with cerebral laceration and contusion, with concussion, unspecified|Other closed skull fracture with cerebral laceration and contusion, with concussion, unspecified
C0159368|T037|HT|803.2|ICD9CM|Other closed skull fracture with subarachnoid, subdural, and extradural hemorrhage|Other closed skull fracture with subarachnoid, subdural, and extradural hemorrhage
C0159369|T037|AB|803.20|ICD9CM|Cl skl fx NEC/mening hem|Cl skl fx NEC/mening hem
C0159370|T037|AB|803.21|ICD9CM|Cl skull fx NEC w/o coma|Cl skull fx NEC w/o coma
C0159371|T037|AB|803.22|ICD9CM|Cl skull fx NEC-brf coma|Cl skull fx NEC-brf coma
C0159372|T037|AB|803.23|ICD9CM|Cl skull fx NEC-mod coma|Cl skull fx NEC-mod coma
C0159373|T037|AB|803.24|ICD9CM|Cl skl fx NEC-proln coma|Cl skl fx NEC-proln coma
C0159374|T037|AB|803.25|ICD9CM|Cl skul fx NEC-deep coma|Cl skul fx NEC-deep coma
C0159375|T037|AB|803.26|ICD9CM|Cl skull fx NEC-coma NOS|Cl skull fx NEC-coma NOS
C0375599|T037|AB|803.29|ICD9CM|Cl skull fx NEC-concuss|Cl skull fx NEC-concuss
C0159377|T037|HT|803.3|ICD9CM|Closed skull fracture with other and unspecified intracranial hemorrhage|Closed skull fracture with other and unspecified intracranial hemorrhage
C0159378|T037|AB|803.30|ICD9CM|Cl skull fx NEC/hem NEC|Cl skull fx NEC/hem NEC
C0159379|T037|AB|803.31|ICD9CM|Cl skull fx NEC w/o coma|Cl skull fx NEC w/o coma
C0159380|T037|AB|803.32|ICD9CM|Cl skull fx NEC-brf coma|Cl skull fx NEC-brf coma
C0159381|T037|AB|803.33|ICD9CM|Cl skull fx NEC-mod coma|Cl skull fx NEC-mod coma
C0159382|T037|AB|803.34|ICD9CM|Cl skl fx NEC-proln coma|Cl skl fx NEC-proln coma
C0159383|T037|AB|803.35|ICD9CM|Cl skul fx NEC-deep coma|Cl skul fx NEC-deep coma
C0159384|T037|AB|803.36|ICD9CM|Cl skull fx NEC-coma NOS|Cl skull fx NEC-coma NOS
C0375600|T037|AB|803.39|ICD9CM|Cl skull fx NEC-concuss|Cl skull fx NEC-concuss
C0159386|T037|HT|803.4|ICD9CM|Other closed skull fracture with intracranial injury of other and unspecified nature|Other closed skull fracture with intracranial injury of other and unspecified nature
C0159387|T037|AB|803.40|ICD9CM|Cl skl fx NEC/br inj NEC|Cl skl fx NEC/br inj NEC
C0159388|T037|AB|803.41|ICD9CM|Cl skull fx NEC w/o coma|Cl skull fx NEC w/o coma
C0159389|T037|AB|803.42|ICD9CM|Cl skull fx NEC-brf coma|Cl skull fx NEC-brf coma
C0159390|T037|AB|803.43|ICD9CM|Cl skull fx NEC-mod coma|Cl skull fx NEC-mod coma
C0159391|T037|AB|803.44|ICD9CM|Cl skl fx NEC-proln coma|Cl skl fx NEC-proln coma
C0159392|T037|AB|803.45|ICD9CM|Cl skul fx NEC-deep coma|Cl skul fx NEC-deep coma
C0159393|T037|AB|803.46|ICD9CM|Cl skull fx NEC-coma NOS|Cl skull fx NEC-coma NOS
C0159394|T037|AB|803.49|ICD9CM|Cl skull fx NEC-concuss|Cl skull fx NEC-concuss
C0159395|T037|HT|803.5|ICD9CM|Other open skull fracture without mention of intracranial injury|Other open skull fracture without mention of intracranial injury
C0159396|T037|AB|803.50|ICD9CM|Open skull fracture NEC|Open skull fracture NEC
C0159396|T037|PT|803.50|ICD9CM|Other open skull fracture without mention of injury, unspecified state of consciousness|Other open skull fracture without mention of injury, unspecified state of consciousness
C0159397|T037|AB|803.51|ICD9CM|Opn skul fx NEC w/o coma|Opn skul fx NEC w/o coma
C0159397|T037|PT|803.51|ICD9CM|Other open skull fracture without mention of intracranial injury, with no loss of consciousness|Other open skull fracture without mention of intracranial injury, with no loss of consciousness
C0159398|T037|AB|803.52|ICD9CM|Opn skul fx NEC-brf coma|Opn skul fx NEC-brf coma
C0159399|T037|AB|803.53|ICD9CM|Opn skul fx NEC-mod coma|Opn skul fx NEC-mod coma
C0159400|T037|AB|803.54|ICD9CM|Opn skl fx NEC-prol coma|Opn skl fx NEC-prol coma
C0159401|T037|AB|803.55|ICD9CM|Opn skl fx NEC-deep coma|Opn skl fx NEC-deep coma
C0159402|T037|AB|803.56|ICD9CM|Opn skul fx NEC-coma NOS|Opn skul fx NEC-coma NOS
C0159403|T037|AB|803.59|ICD9CM|Opn skull fx NEC-concuss|Opn skull fx NEC-concuss
C0159403|T037|PT|803.59|ICD9CM|Other open skull fracture without mention of intracranial injury, with concussion, unspecified|Other open skull fracture without mention of intracranial injury, with concussion, unspecified
C0159404|T037|HT|803.6|ICD9CM|Other open skull fracture with cerebral laceration and contusion|Other open skull fracture with cerebral laceration and contusion
C0159405|T037|AB|803.60|ICD9CM|Opn skl fx NEC/cereb lac|Opn skl fx NEC/cereb lac
C0159405|T037|PT|803.60|ICD9CM|Other open skull fracture with cerebral laceration and contusion, unspecified state of consciousness|Other open skull fracture with cerebral laceration and contusion, unspecified state of consciousness
C0159406|T037|AB|803.61|ICD9CM|Opn skul fx NEC w/o coma|Opn skul fx NEC w/o coma
C0159406|T037|PT|803.61|ICD9CM|Other open skull fracture with cerebral laceration and contusion, with no loss of consciousness|Other open skull fracture with cerebral laceration and contusion, with no loss of consciousness
C0159407|T037|AB|803.62|ICD9CM|Opn skul fx NEC-brf coma|Opn skul fx NEC-brf coma
C0159408|T037|AB|803.63|ICD9CM|Opn skul fx NEC-mod coma|Opn skul fx NEC-mod coma
C0159409|T037|AB|803.64|ICD9CM|Opn skl fx NEC-proln com|Opn skl fx NEC-proln com
C0159410|T037|AB|803.65|ICD9CM|Opn skl fx NEC-deep coma|Opn skl fx NEC-deep coma
C0159411|T037|AB|803.66|ICD9CM|Opn skul fx NEC-coma NOS|Opn skul fx NEC-coma NOS
C0375603|T037|AB|803.69|ICD9CM|Opn skull fx NEC-concuss|Opn skull fx NEC-concuss
C0375603|T037|PT|803.69|ICD9CM|Other open skull fracture with cerebral laceration and contusion, with concussion, unspecified|Other open skull fracture with cerebral laceration and contusion, with concussion, unspecified
C0159413|T037|HT|803.7|ICD9CM|Other open skull fracture with subarachnoid, subdural, and extradural hemorrhage|Other open skull fracture with subarachnoid, subdural, and extradural hemorrhage
C0159414|T037|AB|803.70|ICD9CM|Opn skl fx NEC/menin hem|Opn skl fx NEC/menin hem
C0159415|T037|AB|803.71|ICD9CM|Opn skul fx NEC w/o coma|Opn skul fx NEC w/o coma
C0159416|T037|AB|803.72|ICD9CM|Opn skul fx NEC-brf coma|Opn skul fx NEC-brf coma
C0159417|T037|AB|803.73|ICD9CM|Opn skul fx NEC-mod coma|Opn skul fx NEC-mod coma
C0159418|T037|AB|803.74|ICD9CM|Opn skl fx NEC-prol coma|Opn skl fx NEC-prol coma
C0159419|T037|AB|803.75|ICD9CM|Opn skl fx NEC-deep coma|Opn skl fx NEC-deep coma
C0159420|T037|AB|803.76|ICD9CM|Opn skul fx NEC-coma NOS|Opn skul fx NEC-coma NOS
C0375604|T037|AB|803.79|ICD9CM|Opn skull fx NEC-concuss|Opn skull fx NEC-concuss
C0159422|T037|HT|803.8|ICD9CM|Other open skull fracture with other and unspecified intracranial hemorrhage|Other open skull fracture with other and unspecified intracranial hemorrhage
C0159423|T037|AB|803.80|ICD9CM|Opn skull fx NEC/hem NEC|Opn skull fx NEC/hem NEC
C0159424|T037|AB|803.81|ICD9CM|Opn skul fx NEC w/o coma|Opn skul fx NEC w/o coma
C0159425|T037|AB|803.82|ICD9CM|Opn skul fx NEC-brf coma|Opn skul fx NEC-brf coma
C0159426|T037|AB|803.83|ICD9CM|Opn skul fx NEC-mod coma|Opn skul fx NEC-mod coma
C0159427|T037|AB|803.84|ICD9CM|Opn skl fx NEC-prol coma|Opn skl fx NEC-prol coma
C0159428|T037|AB|803.85|ICD9CM|Opn skl fx NEC-deep coma|Opn skl fx NEC-deep coma
C0159429|T037|AB|803.86|ICD9CM|Opn skul fx NEC-coma NOS|Opn skul fx NEC-coma NOS
C0375605|T037|AB|803.89|ICD9CM|Opn skull fx NEC-concuss|Opn skull fx NEC-concuss
C0159431|T037|HT|803.9|ICD9CM|Other open skull fracture with intracranial injury of other and unspecified nature|Other open skull fracture with intracranial injury of other and unspecified nature
C0159432|T037|AB|803.90|ICD9CM|Op skl fx NEC/br inj NEC|Op skl fx NEC/br inj NEC
C0159433|T037|AB|803.91|ICD9CM|Opn skul fx NEC w/o coma|Opn skul fx NEC w/o coma
C0159434|T037|AB|803.92|ICD9CM|Opn skul fx NEC-brf coma|Opn skul fx NEC-brf coma
C0159435|T037|AB|803.93|ICD9CM|Opn skul fx NEC-mod coma|Opn skul fx NEC-mod coma
C0159436|T037|AB|803.94|ICD9CM|Opn skl fx NEC-prol coma|Opn skl fx NEC-prol coma
C0159437|T037|AB|803.95|ICD9CM|Opn skl fx NEC-deep coma|Opn skl fx NEC-deep coma
C0159438|T037|AB|803.96|ICD9CM|Opn skul fx NEC-coma NOS|Opn skul fx NEC-coma NOS
C0159439|T037|AB|803.99|ICD9CM|Opn skull fx NEC-concuss|Opn skull fx NEC-concuss
C0159440|T037|HT|804|ICD9CM|Multiple fractures involving skull or face with other bones|Multiple fractures involving skull or face with other bones
C0159441|T037|HT|804.0|ICD9CM|Closed fractures involving skull or face with other bones, without mention of intracranial injury|Closed fractures involving skull or face with other bones, without mention of intracranial injury
C0159442|T037|AB|804.00|ICD9CM|Cl skul fx w oth bone fx|Cl skul fx w oth bone fx
C0159443|T037|AB|804.01|ICD9CM|Cl skl w oth fx w/o coma|Cl skl w oth fx w/o coma
C0159444|T037|AB|804.02|ICD9CM|Cl skl w oth fx-brf coma|Cl skl w oth fx-brf coma
C0159445|T037|AB|804.03|ICD9CM|Cl skl w oth fx-mod coma|Cl skl w oth fx-mod coma
C0159446|T037|AB|804.04|ICD9CM|Cl skl/oth fx-proln coma|Cl skl/oth fx-proln coma
C0159447|T037|AB|804.05|ICD9CM|Cl skul/oth fx-deep coma|Cl skul/oth fx-deep coma
C0159448|T037|AB|804.06|ICD9CM|Cl skl w oth fx-coma NOS|Cl skl w oth fx-coma NOS
C0159449|T037|AB|804.09|ICD9CM|Cl skul w oth fx-concuss|Cl skul w oth fx-concuss
C0159450|T037|HT|804.1|ICD9CM|Closed fractures involving skull or face with other bones, with cerebral laceration and contusion|Closed fractures involving skull or face with other bones, with cerebral laceration and contusion
C0159451|T037|AB|804.10|ICD9CM|Cl sk w oth fx/cereb lac|Cl sk w oth fx/cereb lac
C0159452|T037|AB|804.11|ICD9CM|Cl skl w oth fx w/o coma|Cl skl w oth fx w/o coma
C0159453|T037|AB|804.12|ICD9CM|Cl skl w oth fx-brf coma|Cl skl w oth fx-brf coma
C0159454|T037|AB|804.13|ICD9CM|Cl skl w oth fx-mod coma|Cl skl w oth fx-mod coma
C0159455|T037|AB|804.14|ICD9CM|Cl skl/oth fx-proln coma|Cl skl/oth fx-proln coma
C0159456|T037|AB|804.15|ICD9CM|Cl skul/oth fx-deep coma|Cl skul/oth fx-deep coma
C0159457|T037|AB|804.16|ICD9CM|Cl skl w oth fx-coma NOS|Cl skl w oth fx-coma NOS
C0375608|T037|AB|804.19|ICD9CM|Cl skul w oth fx-concuss|Cl skul w oth fx-concuss
C0159460|T037|AB|804.20|ICD9CM|Cl skl/oth fx/mening hem|Cl skl/oth fx/mening hem
C0159461|T037|AB|804.21|ICD9CM|Cl skl w oth fx w/o coma|Cl skl w oth fx w/o coma
C0159462|T037|AB|804.22|ICD9CM|Cl skl w oth fx-brf coma|Cl skl w oth fx-brf coma
C0159463|T037|AB|804.23|ICD9CM|Cl skl w oth fx-mod coma|Cl skl w oth fx-mod coma
C0159464|T037|AB|804.24|ICD9CM|Cl skl/oth fx-proln coma|Cl skl/oth fx-proln coma
C0159465|T037|AB|804.25|ICD9CM|Cl skul/oth fx-deep coma|Cl skul/oth fx-deep coma
C0159466|T037|AB|804.26|ICD9CM|Cl skl w oth fx-coma NOS|Cl skl w oth fx-coma NOS
C0375609|T037|AB|804.29|ICD9CM|Cl skul w oth fx-concuss|Cl skul w oth fx-concuss
C0159469|T037|AB|804.30|ICD9CM|Cl skul w oth fx/hem NEC|Cl skul w oth fx/hem NEC
C0159470|T037|AB|804.31|ICD9CM|Cl skl w oth fx w/o coma|Cl skl w oth fx w/o coma
C0159471|T037|AB|804.32|ICD9CM|Cl skl w oth fx-brf coma|Cl skl w oth fx-brf coma
C0159472|T037|AB|804.33|ICD9CM|Cl skl w oth fx-mod coma|Cl skl w oth fx-mod coma
C0159473|T037|AB|804.34|ICD9CM|Cl skl/oth fx-proln coma|Cl skl/oth fx-proln coma
C0159474|T037|AB|804.35|ICD9CM|Cl skul/oth fx-deep coma|Cl skul/oth fx-deep coma
C0159475|T037|AB|804.36|ICD9CM|Cl skl w oth fx-coma NOS|Cl skl w oth fx-coma NOS
C0375610|T037|AB|804.39|ICD9CM|Cl skul w oth fx-concuss|Cl skul w oth fx-concuss
C0159478|T037|AB|804.40|ICD9CM|Cl skl/oth fx/br inj NEC|Cl skl/oth fx/br inj NEC
C0159479|T037|AB|804.41|ICD9CM|Cl skl w oth fx w/o coma|Cl skl w oth fx w/o coma
C0159480|T037|AB|804.42|ICD9CM|Cl skl w oth fx-brf coma|Cl skl w oth fx-brf coma
C0159481|T037|AB|804.43|ICD9CM|Cl skl w oth fx-mod coma|Cl skl w oth fx-mod coma
C0159482|T037|AB|804.44|ICD9CM|Cl skl/oth fx-proln coma|Cl skl/oth fx-proln coma
C0159483|T037|AB|804.45|ICD9CM|Cl skul/oth fx-deep coma|Cl skul/oth fx-deep coma
C0159484|T037|AB|804.46|ICD9CM|Cl skl w oth fx-coma NOS|Cl skl w oth fx-coma NOS
C0159485|T037|AB|804.49|ICD9CM|Cl skul w oth fx-concuss|Cl skul w oth fx-concuss
C0159486|T037|HT|804.5|ICD9CM|Open fractures involving skull or face with other bones, without mention of intracranial injury|Open fractures involving skull or face with other bones, without mention of intracranial injury
C0159487|T037|AB|804.50|ICD9CM|Opn skull fx/oth bone fx|Opn skull fx/oth bone fx
C0159488|T037|AB|804.51|ICD9CM|Opn skul/oth fx w/o coma|Opn skul/oth fx w/o coma
C0159489|T037|AB|804.52|ICD9CM|Opn skul/oth fx-brf coma|Opn skul/oth fx-brf coma
C0159490|T037|AB|804.53|ICD9CM|Opn skul/oth fx-mod coma|Opn skul/oth fx-mod coma
C0159491|T037|AB|804.54|ICD9CM|Opn skl/oth fx-prol coma|Opn skl/oth fx-prol coma
C0159492|T037|AB|804.55|ICD9CM|Opn skl/oth fx-deep coma|Opn skl/oth fx-deep coma
C0159493|T037|AB|804.56|ICD9CM|Opn skul/oth fx-coma NOS|Opn skul/oth fx-coma NOS
C0159494|T037|AB|804.59|ICD9CM|Opn skull/oth fx-concuss|Opn skull/oth fx-concuss
C0159495|T037|HT|804.6|ICD9CM|Open fractures involving skull or face with other bones, with cerebral laceration and contusion|Open fractures involving skull or face with other bones, with cerebral laceration and contusion
C0159496|T037|AB|804.60|ICD9CM|Opn skl/oth fx/cereb lac|Opn skl/oth fx/cereb lac
C0159497|T037|AB|804.61|ICD9CM|Opn skul/oth fx w/o coma|Opn skul/oth fx w/o coma
C0159498|T037|AB|804.62|ICD9CM|Opn skul/oth fx-brf coma|Opn skul/oth fx-brf coma
C0159499|T037|AB|804.63|ICD9CM|Opn skul/oth fx-mod coma|Opn skul/oth fx-mod coma
C0159500|T037|AB|804.64|ICD9CM|Opn skl/oth fx-prol coma|Opn skl/oth fx-prol coma
C0159501|T037|AB|804.65|ICD9CM|Opn skl/oth fx-deep coma|Opn skl/oth fx-deep coma
C0159502|T037|AB|804.66|ICD9CM|Opn skul/oth fx-coma NOS|Opn skul/oth fx-coma NOS
C0375613|T037|AB|804.69|ICD9CM|Opn skull/oth fx-concuss|Opn skull/oth fx-concuss
C0159505|T037|AB|804.70|ICD9CM|Opn skl/oth fx/menin hem|Opn skl/oth fx/menin hem
C0159506|T037|AB|804.71|ICD9CM|Opn skul/oth fx w/o coma|Opn skul/oth fx w/o coma
C0159507|T037|AB|804.72|ICD9CM|Opn skul/oth fx-brf coma|Opn skul/oth fx-brf coma
C0159508|T037|AB|804.73|ICD9CM|Opn skul/oth fx-mod coma|Opn skul/oth fx-mod coma
C0159509|T037|AB|804.74|ICD9CM|Opn skl/oth fx-prol coma|Opn skl/oth fx-prol coma
C0159510|T037|AB|804.75|ICD9CM|Opn skl/oth fx-deep coma|Opn skl/oth fx-deep coma
C0159511|T037|AB|804.76|ICD9CM|Opn skul/oth fx-coma NOS|Opn skul/oth fx-coma NOS
C0375614|T037|AB|804.79|ICD9CM|Opn skull/oth fx-concuss|Opn skull/oth fx-concuss
C0159514|T037|AB|804.80|ICD9CM|Opn skl w oth fx/hem NEC|Opn skl w oth fx/hem NEC
C0159515|T037|AB|804.81|ICD9CM|Opn skul/oth fx w/o coma|Opn skul/oth fx w/o coma
C0159516|T037|AB|804.82|ICD9CM|Opn skul/oth fx-brf coma|Opn skul/oth fx-brf coma
C0159517|T037|AB|804.83|ICD9CM|Opn skul/oth fx-mod coma|Opn skul/oth fx-mod coma
C0159518|T037|AB|804.84|ICD9CM|Opn skl/oth fx-prol coma|Opn skl/oth fx-prol coma
C0159519|T037|AB|804.85|ICD9CM|Opn skl/oth fx-deep coma|Opn skl/oth fx-deep coma
C0159520|T037|AB|804.86|ICD9CM|Opn skul/oth fx-coma NOS|Opn skul/oth fx-coma NOS
C0375615|T037|AB|804.89|ICD9CM|Opn skull/oth fx-concuss|Opn skull/oth fx-concuss
C0159523|T037|AB|804.90|ICD9CM|Op skl/oth fx/br inj NEC|Op skl/oth fx/br inj NEC
C0159524|T037|AB|804.91|ICD9CM|Opn skul/oth fx w/o coma|Opn skul/oth fx w/o coma
C0159525|T037|AB|804.92|ICD9CM|Opn skul/oth fx-brf coma|Opn skul/oth fx-brf coma
C0159526|T037|AB|804.93|ICD9CM|Opn skul/oth fx-mod coma|Opn skul/oth fx-mod coma
C0159527|T037|AB|804.94|ICD9CM|Opn skl/oth fx-prol coma|Opn skl/oth fx-prol coma
C0159528|T037|AB|804.95|ICD9CM|Opn skl/oth fx-deep coma|Opn skl/oth fx-deep coma
C0159529|T037|AB|804.96|ICD9CM|Opn skul/oth fx-coma NOS|Opn skul/oth fx-coma NOS
C0159530|T037|AB|804.99|ICD9CM|Opn skull/oth fx-concuss|Opn skull/oth fx-concuss
C0559043|T037|HT|805|ICD9CM|Fracture of vertebral column without mention of spinal cord injury|Fracture of vertebral column without mention of spinal cord injury
C0178315|T037|HT|805-809.99|ICD9CM|FRACTURE OF NECK AND TRUNK|FRACTURE OF NECK AND TRUNK
C0859693|T037|HT|805.0|ICD9CM|Closed fracture of cervical vertebra without mention of spinal cord injury|Closed fracture of cervical vertebra without mention of spinal cord injury
C0375617|T037|PT|805.00|ICD9CM|Closed fracture of cervical vertebra, unspecified level|Closed fracture of cervical vertebra, unspecified level
C0375617|T037|AB|805.00|ICD9CM|Fx cervical vert NOS-cl|Fx cervical vert NOS-cl
C0159533|T037|PT|805.01|ICD9CM|Closed fracture of first cervical vertebra|Closed fracture of first cervical vertebra
C0159533|T037|AB|805.01|ICD9CM|Fx c1 vertebra-closed|Fx c1 vertebra-closed
C0159534|T037|PT|805.02|ICD9CM|Closed fracture of second cervical vertebra|Closed fracture of second cervical vertebra
C0159534|T037|AB|805.02|ICD9CM|Fx c2 vertebra-closed|Fx c2 vertebra-closed
C0159535|T037|PT|805.03|ICD9CM|Closed fracture of third cervical vertebra|Closed fracture of third cervical vertebra
C0159535|T037|AB|805.03|ICD9CM|Fx c3 vertebra-closed|Fx c3 vertebra-closed
C0159536|T037|PT|805.04|ICD9CM|Closed fracture of fourth cervical vertebra|Closed fracture of fourth cervical vertebra
C0159536|T037|AB|805.04|ICD9CM|Fx c4 vertebra-closed|Fx c4 vertebra-closed
C0159537|T037|PT|805.05|ICD9CM|Closed fracture of fifth cervical vertebra|Closed fracture of fifth cervical vertebra
C0159537|T037|AB|805.05|ICD9CM|Fx c5 vertebra-closed|Fx c5 vertebra-closed
C0159538|T037|PT|805.06|ICD9CM|Closed fracture of sixth cervical vertebra|Closed fracture of sixth cervical vertebra
C0159538|T037|AB|805.06|ICD9CM|Fx c6 vertebra-closed|Fx c6 vertebra-closed
C0159539|T037|PT|805.07|ICD9CM|Closed fracture of seventh cervical vertebra|Closed fracture of seventh cervical vertebra
C0159539|T037|AB|805.07|ICD9CM|Fx c7 vertebra-closed|Fx c7 vertebra-closed
C0159540|T037|PT|805.08|ICD9CM|Closed fracture of multiple cervical vertebrae|Closed fracture of multiple cervical vertebrae
C0159540|T037|AB|805.08|ICD9CM|Fx mult cervical vert-cl|Fx mult cervical vert-cl
C0859694|T037|HT|805.1|ICD9CM|Open fracture of cervical vertebra without mention of spinal cord injury|Open fracture of cervical vertebra without mention of spinal cord injury
C0375618|T037|AB|805.10|ICD9CM|Fx cervical vert NOS-opn|Fx cervical vert NOS-opn
C0375618|T037|PT|805.10|ICD9CM|Open fracture of cervical vertebra, unspecified level|Open fracture of cervical vertebra, unspecified level
C0159543|T037|AB|805.11|ICD9CM|Fx c1 vertebra-open|Fx c1 vertebra-open
C0159543|T037|PT|805.11|ICD9CM|Open fracture of first cervical vertebra|Open fracture of first cervical vertebra
C0159544|T037|AB|805.12|ICD9CM|Fx c2 vertebra-open|Fx c2 vertebra-open
C0159544|T037|PT|805.12|ICD9CM|Open fracture of second cervical vertebra|Open fracture of second cervical vertebra
C0159545|T037|AB|805.13|ICD9CM|Fx c3 vertebra-open|Fx c3 vertebra-open
C0159545|T037|PT|805.13|ICD9CM|Open fracture of third cervical vertebra|Open fracture of third cervical vertebra
C0159546|T037|AB|805.14|ICD9CM|Fx c4 vertebra-open|Fx c4 vertebra-open
C0159546|T037|PT|805.14|ICD9CM|Open fracture of fourth cervical vertebra|Open fracture of fourth cervical vertebra
C0159547|T037|AB|805.15|ICD9CM|Fx c5 vertebra-open|Fx c5 vertebra-open
C0159547|T037|PT|805.15|ICD9CM|Open fracture of fifth cervical vertebra|Open fracture of fifth cervical vertebra
C0159548|T037|AB|805.16|ICD9CM|Fx c6 vertebra-open|Fx c6 vertebra-open
C0159548|T037|PT|805.16|ICD9CM|Open fracture of sixth cervical vertebra|Open fracture of sixth cervical vertebra
C0159549|T037|AB|805.17|ICD9CM|Fx c7 vertebra-open|Fx c7 vertebra-open
C0159549|T037|PT|805.17|ICD9CM|Open fracture of seventh cervical vertebra|Open fracture of seventh cervical vertebra
C0159550|T037|AB|805.18|ICD9CM|Fx mlt cervical vert-opn|Fx mlt cervical vert-opn
C0159550|T037|PT|805.18|ICD9CM|Open fracture of multiple cervical vertebrae|Open fracture of multiple cervical vertebrae
C0159551|T037|PT|805.2|ICD9CM|Closed fracture of dorsal [thoracic] vertebra without mention of spinal cord injury|Closed fracture of dorsal [thoracic] vertebra without mention of spinal cord injury
C0159551|T037|AB|805.2|ICD9CM|Fx dorsal vertebra-close|Fx dorsal vertebra-close
C0159552|T037|AB|805.3|ICD9CM|Fx dorsal vertebra-open|Fx dorsal vertebra-open
C0159552|T037|PT|805.3|ICD9CM|Open fracture of dorsal [thoracic] vertebra without mention of spinal cord injury|Open fracture of dorsal [thoracic] vertebra without mention of spinal cord injury
C0859697|T037|PT|805.4|ICD9CM|Closed fracture of lumbar vertebra without mention of spinal cord injury|Closed fracture of lumbar vertebra without mention of spinal cord injury
C0859697|T037|AB|805.4|ICD9CM|Fx lumbar vertebra-close|Fx lumbar vertebra-close
C0859698|T037|AB|805.5|ICD9CM|Fx lumbar vertebra-open|Fx lumbar vertebra-open
C0859698|T037|PT|805.5|ICD9CM|Open fracture of lumbar vertebra without mention of spinal cord injury|Open fracture of lumbar vertebra without mention of spinal cord injury
C0159555|T037|PT|805.6|ICD9CM|Closed fracture of sacrum and coccyx without mention of spinal cord injury|Closed fracture of sacrum and coccyx without mention of spinal cord injury
C0159555|T037|AB|805.6|ICD9CM|Fx sacrum/coccyx-closed|Fx sacrum/coccyx-closed
C0159556|T037|AB|805.7|ICD9CM|Fx sacrum/coccyx-open|Fx sacrum/coccyx-open
C0159556|T037|PT|805.7|ICD9CM|Open fracture of sacrum and coccyx without mention of spinal cord injury|Open fracture of sacrum and coccyx without mention of spinal cord injury
C0009048|T037|PT|805.8|ICD9CM|Closed fracture of unspecified vertebral column without mention of spinal cord injury|Closed fracture of unspecified vertebral column without mention of spinal cord injury
C0009048|T037|AB|805.8|ICD9CM|Vertebral fx NOS-closed|Vertebral fx NOS-closed
C0159557|T037|PT|805.9|ICD9CM|Open fracture of unspecified vertebral column without mention of spinal cord injury|Open fracture of unspecified vertebral column without mention of spinal cord injury
C0159557|T037|AB|805.9|ICD9CM|Vertebral fx NOS-open|Vertebral fx NOS-open
C0435349|T037|HT|806|ICD9CM|Fracture of vertebral column with spinal cord injury|Fracture of vertebral column with spinal cord injury
C0859703|T037|HT|806.0|ICD9CM|Closed fracture of cervical vertebra with spinal cord injury|Closed fracture of cervical vertebra with spinal cord injury
C0159560|T037|AB|806.00|ICD9CM|C1-c4 fx-cl/cord inj NOS|C1-c4 fx-cl/cord inj NOS
C0159560|T037|PT|806.00|ICD9CM|Closed fracture of C1-C4 level with unspecified spinal cord injury|Closed fracture of C1-C4 level with unspecified spinal cord injury
C0435397|T037|AB|806.01|ICD9CM|C1-c4 fx-cl/com cord les|C1-c4 fx-cl/com cord les
C0435397|T037|PT|806.01|ICD9CM|Closed fracture of C1-C4 level with complete lesion of cord|Closed fracture of C1-C4 level with complete lesion of cord
C0159562|T037|AB|806.02|ICD9CM|C1-c4 fx-cl/ant cord syn|C1-c4 fx-cl/ant cord syn
C0159562|T037|PT|806.02|ICD9CM|Closed fracture of C1-C4 level with anterior cord syndrome|Closed fracture of C1-C4 level with anterior cord syndrome
C0159563|T037|AB|806.03|ICD9CM|C1-c4 fx-cl/cen cord syn|C1-c4 fx-cl/cen cord syn
C0159563|T037|PT|806.03|ICD9CM|Closed fracture of C1-C4 level with central cord syndrome|Closed fracture of C1-C4 level with central cord syndrome
C0159564|T037|AB|806.04|ICD9CM|C1-c4 fx-cl/cord inj NEC|C1-c4 fx-cl/cord inj NEC
C0159564|T037|PT|806.04|ICD9CM|Closed fracture of C1-C4 level with other specified spinal cord injury|Closed fracture of C1-C4 level with other specified spinal cord injury
C0159565|T037|AB|806.05|ICD9CM|C5-c7 fx-cl/cord inj NOS|C5-c7 fx-cl/cord inj NOS
C0159565|T037|PT|806.05|ICD9CM|Closed fracture of C5-C7 level with unspecified spinal cord injury|Closed fracture of C5-C7 level with unspecified spinal cord injury
C0435403|T037|AB|806.06|ICD9CM|C5-c7 fx-cl/com cord les|C5-c7 fx-cl/com cord les
C0435403|T037|PT|806.06|ICD9CM|Closed fracture of C5-C7 level with complete lesion of cord|Closed fracture of C5-C7 level with complete lesion of cord
C0159567|T037|AB|806.07|ICD9CM|C5-c7 fx-cl/ant cord syn|C5-c7 fx-cl/ant cord syn
C0159567|T037|PT|806.07|ICD9CM|Closed fracture of C5-C7 level with anterior cord syndrome|Closed fracture of C5-C7 level with anterior cord syndrome
C0159568|T037|AB|806.08|ICD9CM|C5-c7 fx-cl/cen cord syn|C5-c7 fx-cl/cen cord syn
C0159568|T037|PT|806.08|ICD9CM|Closed fracture of C5-C7 level with central cord syndrome|Closed fracture of C5-C7 level with central cord syndrome
C0159569|T037|AB|806.09|ICD9CM|C5-c7 fx-cl/cord inj NEC|C5-c7 fx-cl/cord inj NEC
C0159569|T037|PT|806.09|ICD9CM|Closed fracture of C5-C7 level with other specified spinal cord injury|Closed fracture of C5-C7 level with other specified spinal cord injury
C0859704|T037|HT|806.1|ICD9CM|Open fracture of cervical vertebra with spinal cord injury|Open fracture of cervical vertebra with spinal cord injury
C0159571|T037|AB|806.10|ICD9CM|C1-c4 fx-op/cord inj NOS|C1-c4 fx-op/cord inj NOS
C0159571|T037|PT|806.10|ICD9CM|Open fracture of C1-C4 level with unspecified spinal cord injury|Open fracture of C1-C4 level with unspecified spinal cord injury
C0435410|T037|AB|806.11|ICD9CM|C1-c4 fx-op/com cord les|C1-c4 fx-op/com cord les
C0435410|T037|PT|806.11|ICD9CM|Open fracture of C1-C4 level with complete lesion of cord|Open fracture of C1-C4 level with complete lesion of cord
C0159573|T037|AB|806.12|ICD9CM|C1-c4 fx-op/ant cord syn|C1-c4 fx-op/ant cord syn
C0159573|T037|PT|806.12|ICD9CM|Open fracture of C1-C4 level with anterior cord syndrome|Open fracture of C1-C4 level with anterior cord syndrome
C0159574|T037|AB|806.13|ICD9CM|C1-c4 fx-op/cen cord syn|C1-c4 fx-op/cen cord syn
C0159574|T037|PT|806.13|ICD9CM|Open fracture of C1-C4 level with central cord syndrome|Open fracture of C1-C4 level with central cord syndrome
C0159575|T037|AB|806.14|ICD9CM|C1-c4 fx-op/cord inj NEC|C1-c4 fx-op/cord inj NEC
C0159575|T037|PT|806.14|ICD9CM|Open fracture of C1-C4 level with other specified spinal cord injury|Open fracture of C1-C4 level with other specified spinal cord injury
C0159576|T037|AB|806.15|ICD9CM|C5-c7 fx-op/cord inj NOS|C5-c7 fx-op/cord inj NOS
C0159576|T037|PT|806.15|ICD9CM|Open fracture of C5-C7 level with unspecified spinal cord injury|Open fracture of C5-C7 level with unspecified spinal cord injury
C0435416|T037|AB|806.16|ICD9CM|C5-c7 fx-op/com cord les|C5-c7 fx-op/com cord les
C0435416|T037|PT|806.16|ICD9CM|Open fracture of C5-C7 level with complete lesion of cord|Open fracture of C5-C7 level with complete lesion of cord
C0159578|T037|AB|806.17|ICD9CM|C5-c7 fx-op/ant cord syn|C5-c7 fx-op/ant cord syn
C0159578|T037|PT|806.17|ICD9CM|Open fracture of C5-C7 level with anterior cord syndrome|Open fracture of C5-C7 level with anterior cord syndrome
C0159579|T037|AB|806.18|ICD9CM|C5-c7 fx-op/cen cord syn|C5-c7 fx-op/cen cord syn
C0159579|T037|PT|806.18|ICD9CM|Open fracture of C5-C7 level with central cord syndrome|Open fracture of C5-C7 level with central cord syndrome
C0159580|T037|AB|806.19|ICD9CM|C5-c7 fx-op/cord inj NEC|C5-c7 fx-op/cord inj NEC
C0159580|T037|PT|806.19|ICD9CM|Open fracture of C5-C7 level with other specified spinal cord injury|Open fracture of C5-C7 level with other specified spinal cord injury
C0859705|T037|HT|806.2|ICD9CM|Closed fracture of dorsal vertebra with spinal cord injury|Closed fracture of dorsal vertebra with spinal cord injury
C0159582|T037|PT|806.20|ICD9CM|Closed fracture of T1-T6 level with unspecified spinal cord injury|Closed fracture of T1-T6 level with unspecified spinal cord injury
C0159582|T037|AB|806.20|ICD9CM|T1-t6 fx-cl/cord inj NOS|T1-t6 fx-cl/cord inj NOS
C0435439|T037|PT|806.21|ICD9CM|Closed fracture of T1-T6 level with complete lesion of cord|Closed fracture of T1-T6 level with complete lesion of cord
C0435439|T037|AB|806.21|ICD9CM|T1-t6 fx-cl/com cord les|T1-t6 fx-cl/com cord les
C0159584|T037|PT|806.22|ICD9CM|Closed fracture of T1-T6 level with anterior cord syndrome|Closed fracture of T1-T6 level with anterior cord syndrome
C0159584|T037|AB|806.22|ICD9CM|T1-t6 fx-cl/ant cord syn|T1-t6 fx-cl/ant cord syn
C0159585|T037|PT|806.23|ICD9CM|Closed fracture of T1-T6 level with central cord syndrome|Closed fracture of T1-T6 level with central cord syndrome
C0159585|T037|AB|806.23|ICD9CM|T1-t6 fx-cl/cen cord syn|T1-t6 fx-cl/cen cord syn
C0159586|T037|PT|806.24|ICD9CM|Closed fracture of T1-T6 level with other specified spinal cord injury|Closed fracture of T1-T6 level with other specified spinal cord injury
C0159586|T037|AB|806.24|ICD9CM|T1-t6 fx-cl/cord inj NEC|T1-t6 fx-cl/cord inj NEC
C0159587|T037|PT|806.25|ICD9CM|Closed fracture of T7-T12 level with unspecified spinal cord injury|Closed fracture of T7-T12 level with unspecified spinal cord injury
C0159587|T037|AB|806.25|ICD9CM|T7-t12 fx-cl/crd inj NOS|T7-t12 fx-cl/crd inj NOS
C0435445|T037|PT|806.26|ICD9CM|Closed fracture of T7-T12 level with complete lesion of cord|Closed fracture of T7-T12 level with complete lesion of cord
C0435445|T037|AB|806.26|ICD9CM|T7-t12 fx-cl/com crd les|T7-t12 fx-cl/com crd les
C0159589|T037|PT|806.27|ICD9CM|Closed fracture of T7-T12 level with anterior cord syndrome|Closed fracture of T7-T12 level with anterior cord syndrome
C0159589|T037|AB|806.27|ICD9CM|T7-t12 fx-cl/ant crd syn|T7-t12 fx-cl/ant crd syn
C0159590|T037|PT|806.28|ICD9CM|Closed fracture of T7-T12 level with central cord syndrome|Closed fracture of T7-T12 level with central cord syndrome
C0159590|T037|AB|806.28|ICD9CM|T7-t12 fx-cl/cen crd syn|T7-t12 fx-cl/cen crd syn
C0159591|T037|PT|806.29|ICD9CM|Closed fracture of T7-T12 level with other specified spinal cord injury|Closed fracture of T7-T12 level with other specified spinal cord injury
C0159591|T037|AB|806.29|ICD9CM|T7-t12 fx-cl/crd inj NEC|T7-t12 fx-cl/crd inj NEC
C0859706|T037|HT|806.3|ICD9CM|Open fracture of dorsal vertebra with spinal cord injury|Open fracture of dorsal vertebra with spinal cord injury
C0159593|T037|PT|806.30|ICD9CM|Open fracture of T1-T6 level with unspecified spinal cord injury|Open fracture of T1-T6 level with unspecified spinal cord injury
C0159593|T037|AB|806.30|ICD9CM|T1-t6 fx-op/cord inj NOS|T1-t6 fx-op/cord inj NOS
C0435452|T037|PT|806.31|ICD9CM|Open fracture of T1-T6 level with complete lesion of cord|Open fracture of T1-T6 level with complete lesion of cord
C0435452|T037|AB|806.31|ICD9CM|T1-t6 fx-op/com cord les|T1-t6 fx-op/com cord les
C0159595|T037|PT|806.32|ICD9CM|Open fracture of T1-T6 level with anterior cord syndrome|Open fracture of T1-T6 level with anterior cord syndrome
C0159595|T037|AB|806.32|ICD9CM|T1-t6 fx-op/ant cord syn|T1-t6 fx-op/ant cord syn
C0159596|T037|PT|806.33|ICD9CM|Open fracture of T1-T6 level with central cord syndrome|Open fracture of T1-T6 level with central cord syndrome
C0159596|T037|AB|806.33|ICD9CM|T1-t6 fx-op/cen cord syn|T1-t6 fx-op/cen cord syn
C0159597|T037|PT|806.34|ICD9CM|Open fracture of T1-T6 level with other specified spinal cord injury|Open fracture of T1-T6 level with other specified spinal cord injury
C0159597|T037|AB|806.34|ICD9CM|T1-t6 fx-op/cord inj NEC|T1-t6 fx-op/cord inj NEC
C0159598|T037|PT|806.35|ICD9CM|Open fracture of T7-T12 level with unspecified spinal cord injury|Open fracture of T7-T12 level with unspecified spinal cord injury
C0159598|T037|AB|806.35|ICD9CM|T7-t12 fx-op/crd inj NOS|T7-t12 fx-op/crd inj NOS
C0435457|T037|PT|806.36|ICD9CM|Open fracture of T7-T12 level with complete lesion of cord|Open fracture of T7-T12 level with complete lesion of cord
C0435457|T037|AB|806.36|ICD9CM|T7-t12 fx-op/com crd les|T7-t12 fx-op/com crd les
C0159600|T037|PT|806.37|ICD9CM|Open fracture of T7-T12 level with anterior cord syndrome|Open fracture of T7-T12 level with anterior cord syndrome
C0159600|T037|AB|806.37|ICD9CM|T7-t12 fx-op/ant crd syn|T7-t12 fx-op/ant crd syn
C0159601|T037|PT|806.38|ICD9CM|Open fracture of T7-T12 level with central cord syndrome|Open fracture of T7-T12 level with central cord syndrome
C0159601|T037|AB|806.38|ICD9CM|T7-t12 fx-op/cen crd syn|T7-t12 fx-op/cen crd syn
C0159602|T037|PT|806.39|ICD9CM|Open fracture of T7-T12 level with other specified spinal cord injury|Open fracture of T7-T12 level with other specified spinal cord injury
C0159602|T037|AB|806.39|ICD9CM|T7-t12 fx-op/crd inj NEC|T7-t12 fx-op/crd inj NEC
C3665459|T037|AB|806.4|ICD9CM|Cl lumbar fx w cord inj|Cl lumbar fx w cord inj
C3665459|T037|PT|806.4|ICD9CM|Closed fracture of lumbar spine with spinal cord injury|Closed fracture of lumbar spine with spinal cord injury
C0435484|T037|PT|806.5|ICD9CM|Open fracture of lumbar spine with spinal cord injury|Open fracture of lumbar spine with spinal cord injury
C0435484|T037|AB|806.5|ICD9CM|Opn lumbar fx w cord inj|Opn lumbar fx w cord inj
C0159606|T037|HT|806.6|ICD9CM|Closed fracture of sacrum and coccyx with spinal cord injury|Closed fracture of sacrum and coccyx with spinal cord injury
C0159606|T037|PT|806.60|ICD9CM|Closed fracture of sacrum and coccyx with unspecified spinal cord injury|Closed fracture of sacrum and coccyx with unspecified spinal cord injury
C0159606|T037|AB|806.60|ICD9CM|Fx sacrum-cl/crd inj NOS|Fx sacrum-cl/crd inj NOS
C0159607|T037|PT|806.61|ICD9CM|Closed fracture of sacrum and coccyx with complete cauda equina lesion|Closed fracture of sacrum and coccyx with complete cauda equina lesion
C0159607|T037|AB|806.61|ICD9CM|Fx sacr-cl/cauda equ les|Fx sacr-cl/cauda equ les
C0159608|T037|PT|806.62|ICD9CM|Closed fracture of sacrum and coccyx with other cauda equina injury|Closed fracture of sacrum and coccyx with other cauda equina injury
C0159608|T037|AB|806.62|ICD9CM|Fx sacr-cl/cauda inj NEC|Fx sacr-cl/cauda inj NEC
C0159609|T037|PT|806.69|ICD9CM|Closed fracture of sacrum and coccyx with other spinal cord injury|Closed fracture of sacrum and coccyx with other spinal cord injury
C0159609|T037|AB|806.69|ICD9CM|Fx sacrum-cl/crd inj NEC|Fx sacrum-cl/crd inj NEC
C0159611|T037|HT|806.7|ICD9CM|Open fracture of sacrum and coccyx with spinal cord injury|Open fracture of sacrum and coccyx with spinal cord injury
C0159611|T037|AB|806.70|ICD9CM|Fx sacrum-op/crd inj NOS|Fx sacrum-op/crd inj NOS
C0159611|T037|PT|806.70|ICD9CM|Open fracture of sacrum and coccyx with unspecified spinal cord injury|Open fracture of sacrum and coccyx with unspecified spinal cord injury
C0159612|T037|AB|806.71|ICD9CM|Fx sacr-op/cauda equ les|Fx sacr-op/cauda equ les
C0159612|T037|PT|806.71|ICD9CM|Open fracture of sacrum and coccyx with complete cauda equina lesion|Open fracture of sacrum and coccyx with complete cauda equina lesion
C0159613|T037|AB|806.72|ICD9CM|Fx sacr-op/cauda inj NEC|Fx sacr-op/cauda inj NEC
C0159613|T037|PT|806.72|ICD9CM|Open fracture of sacrum and coccyx with other cauda equina injury|Open fracture of sacrum and coccyx with other cauda equina injury
C0159614|T037|AB|806.79|ICD9CM|Fx sacrum-op/crd inj NEC|Fx sacrum-op/crd inj NEC
C0159614|T037|PT|806.79|ICD9CM|Open fracture of sacrum and coccyx with other spinal cord injury|Open fracture of sacrum and coccyx with other spinal cord injury
C0159615|T037|PT|806.8|ICD9CM|Closed fracture of unspecified vertebral column with spinal cord injury|Closed fracture of unspecified vertebral column with spinal cord injury
C0159615|T037|AB|806.8|ICD9CM|Vert fx NOS-cl w crd inj|Vert fx NOS-cl w crd inj
C0159616|T037|PT|806.9|ICD9CM|Open fracture of unspecified vertebral column with spinal cord injury|Open fracture of unspecified vertebral column with spinal cord injury
C0159616|T037|AB|806.9|ICD9CM|Vert fx NOS-op w crd inj|Vert fx NOS-op w crd inj
C0159617|T037|HT|807|ICD9CM|Fracture of rib(s), sternum, larynx, and trachea|Fracture of rib(s), sternum, larynx, and trachea
C0435750|T037|HT|807.0|ICD9CM|Closed fracture of rib(s)|Closed fracture of rib(s)
C0435750|T037|PT|807.00|ICD9CM|Closed fracture of rib(s), unspecified|Closed fracture of rib(s), unspecified
C0435750|T037|AB|807.00|ICD9CM|Fracture rib NOS-closed|Fracture rib NOS-closed
C0159618|T037|PT|807.01|ICD9CM|Closed fracture of one rib|Closed fracture of one rib
C0159618|T037|AB|807.01|ICD9CM|Fracture one rib-closed|Fracture one rib-closed
C0159619|T037|PT|807.02|ICD9CM|Closed fracture of two ribs|Closed fracture of two ribs
C0159619|T037|AB|807.02|ICD9CM|Fracture two ribs-closed|Fracture two ribs-closed
C0159620|T037|PT|807.03|ICD9CM|Closed fracture of three ribs|Closed fracture of three ribs
C0159620|T037|AB|807.03|ICD9CM|Fracture three ribs-clos|Fracture three ribs-clos
C0159621|T037|PT|807.04|ICD9CM|Closed fracture of four ribs|Closed fracture of four ribs
C0159621|T037|AB|807.04|ICD9CM|Fracture four ribs-close|Fracture four ribs-close
C0159622|T037|PT|807.05|ICD9CM|Closed fracture of five ribs|Closed fracture of five ribs
C0159622|T037|AB|807.05|ICD9CM|Fracture five ribs-close|Fracture five ribs-close
C0159623|T037|PT|807.06|ICD9CM|Closed fracture of six ribs|Closed fracture of six ribs
C0159623|T037|AB|807.06|ICD9CM|Fracture six ribs-closed|Fracture six ribs-closed
C0159624|T037|PT|807.07|ICD9CM|Closed fracture of seven ribs|Closed fracture of seven ribs
C0159624|T037|AB|807.07|ICD9CM|Fracture seven ribs-clos|Fracture seven ribs-clos
C0159625|T037|PT|807.08|ICD9CM|Closed fracture of eight or more ribs|Closed fracture of eight or more ribs
C0159625|T037|AB|807.08|ICD9CM|Fx eight/more rib-closed|Fx eight/more rib-closed
C0159626|T037|PT|807.09|ICD9CM|Closed fracture of multiple ribs, unspecified|Closed fracture of multiple ribs, unspecified
C0159626|T037|AB|807.09|ICD9CM|Fx mult ribs NOS-closed|Fx mult ribs NOS-closed
C0435751|T037|HT|807.1|ICD9CM|Open fracture of rib(s)|Open fracture of rib(s)
C0435751|T037|AB|807.10|ICD9CM|Fracture rib NOS-open|Fracture rib NOS-open
C0435751|T037|PT|807.10|ICD9CM|Open fracture of rib(s), unspecified|Open fracture of rib(s), unspecified
C0159628|T037|AB|807.11|ICD9CM|Fracture one rib-open|Fracture one rib-open
C0159628|T037|PT|807.11|ICD9CM|Open fracture of one rib|Open fracture of one rib
C0159629|T037|AB|807.12|ICD9CM|Fracture two ribs-open|Fracture two ribs-open
C0159629|T037|PT|807.12|ICD9CM|Open fracture of two ribs|Open fracture of two ribs
C0159630|T037|AB|807.13|ICD9CM|Fracture three ribs-open|Fracture three ribs-open
C0159630|T037|PT|807.13|ICD9CM|Open fracture of three ribs|Open fracture of three ribs
C0159631|T037|AB|807.14|ICD9CM|Fracture four ribs-open|Fracture four ribs-open
C0159631|T037|PT|807.14|ICD9CM|Open fracture of four ribs|Open fracture of four ribs
C0159632|T037|AB|807.15|ICD9CM|Fracture five ribs-open|Fracture five ribs-open
C0159632|T037|PT|807.15|ICD9CM|Open fracture of five ribs|Open fracture of five ribs
C0159633|T037|AB|807.16|ICD9CM|Fracture six ribs-open|Fracture six ribs-open
C0159633|T037|PT|807.16|ICD9CM|Open fracture of six ribs|Open fracture of six ribs
C0159634|T037|AB|807.17|ICD9CM|Fracture seven ribs-open|Fracture seven ribs-open
C0159634|T037|PT|807.17|ICD9CM|Open fracture of seven ribs|Open fracture of seven ribs
C0159635|T037|AB|807.18|ICD9CM|Fx eight/more ribs-open|Fx eight/more ribs-open
C0159635|T037|PT|807.18|ICD9CM|Open fracture of eight or more ribs|Open fracture of eight or more ribs
C0159636|T037|AB|807.19|ICD9CM|Fx mult ribs NOS-open|Fx mult ribs NOS-open
C0159636|T037|PT|807.19|ICD9CM|Open fracture of multiple ribs, unspecified|Open fracture of multiple ribs, unspecified
C0159637|T037|PT|807.2|ICD9CM|Closed fracture of sternum|Closed fracture of sternum
C0159637|T037|AB|807.2|ICD9CM|Fracture of sternum-clos|Fracture of sternum-clos
C0159638|T037|AB|807.3|ICD9CM|Fracture of sternum-open|Fracture of sternum-open
C0159638|T037|PT|807.3|ICD9CM|Open fracture of sternum|Open fracture of sternum
C0016196|T037|AB|807.4|ICD9CM|Flail chest|Flail chest
C0016196|T037|PT|807.4|ICD9CM|Flail chest|Flail chest
C0159639|T037|PT|807.5|ICD9CM|Closed fracture of larynx and trachea|Closed fracture of larynx and trachea
C0159639|T037|AB|807.5|ICD9CM|Fx larynx/trachea-closed|Fx larynx/trachea-closed
C0159640|T037|AB|807.6|ICD9CM|Fx larynx/trachea-open|Fx larynx/trachea-open
C0159640|T037|PT|807.6|ICD9CM|Open fracture of larynx and trachea|Open fracture of larynx and trachea
C0149531|T037|HT|808|ICD9CM|Fracture of pelvis|Fracture of pelvis
C0159641|T037|PT|808.0|ICD9CM|Closed fracture of acetabulum|Closed fracture of acetabulum
C0159641|T037|AB|808.0|ICD9CM|Fracture acetabulum-clos|Fracture acetabulum-clos
C0159642|T037|AB|808.1|ICD9CM|Fracture acetabulum-open|Fracture acetabulum-open
C0159642|T037|PT|808.1|ICD9CM|Open fracture of acetabulum|Open fracture of acetabulum
C0159643|T037|PT|808.2|ICD9CM|Closed fracture of pubis|Closed fracture of pubis
C0159643|T037|AB|808.2|ICD9CM|Fracture of pubis-closed|Fracture of pubis-closed
C0159644|T037|AB|808.3|ICD9CM|Fracture of pubis-open|Fracture of pubis-open
C0159644|T037|PT|808.3|ICD9CM|Open fracture of pubis|Open fracture of pubis
C0159645|T037|HT|808.4|ICD9CM|Closed fracture of other specified part of pelvis|Closed fracture of other specified part of pelvis
C0159646|T037|PT|808.41|ICD9CM|Closed fracture of ilium|Closed fracture of ilium
C0159646|T037|AB|808.41|ICD9CM|Fracture of ilium-closed|Fracture of ilium-closed
C0159647|T037|PT|808.42|ICD9CM|Closed fracture of ischium|Closed fracture of ischium
C0159647|T037|AB|808.42|ICD9CM|Fracture ischium-closed|Fracture ischium-closed
C0272580|T037|PT|808.43|ICD9CM|Multiple closed pelvic fractures with disruption of pelvic circle|Multiple closed pelvic fractures with disruption of pelvic circle
C0272580|T037|AB|808.43|ICD9CM|Pelv fx-clos/pelv disrup|Pelv fx-clos/pelv disrup
C3161129|T037|PT|808.44|ICD9CM|Multiple closed pelvic fractures without disruption of pelvic circle|Multiple closed pelvic fractures without disruption of pelvic circle
C3161129|T037|AB|808.44|ICD9CM|Pelv fx-cl w/o plv disrp|Pelv fx-cl w/o plv disrp
C0159645|T037|PT|808.49|ICD9CM|Closed fracture of other specified part of pelvis|Closed fracture of other specified part of pelvis
C0159645|T037|AB|808.49|ICD9CM|Pelvic fracture NEC-clos|Pelvic fracture NEC-clos
C0159649|T037|HT|808.5|ICD9CM|Open fracture of other specified part of pelvis|Open fracture of other specified part of pelvis
C0435771|T037|AB|808.51|ICD9CM|Fracture of ilium-open|Fracture of ilium-open
C0435771|T037|PT|808.51|ICD9CM|Open fracture of ilium|Open fracture of ilium
C0159651|T037|AB|808.52|ICD9CM|Fracture of ischium-open|Fracture of ischium-open
C0159651|T037|PT|808.52|ICD9CM|Open fracture of ischium|Open fracture of ischium
C0272582|T037|PT|808.53|ICD9CM|Multiple open pelvic fractures with disruption of pelvic circle|Multiple open pelvic fractures with disruption of pelvic circle
C0272582|T037|AB|808.53|ICD9CM|Pelv fx-open/pelv disrup|Pelv fx-open/pelv disrup
C3161130|T037|PT|808.54|ICD9CM|Multiple open pelvic fractures without disruption of pelvic circle|Multiple open pelvic fractures without disruption of pelvic circle
C3161130|T037|AB|808.54|ICD9CM|Pelv fx-opn w/o pelv dis|Pelv fx-opn w/o pelv dis
C0159649|T037|PT|808.59|ICD9CM|Open fracture of other specified part of pelvis|Open fracture of other specified part of pelvis
C0159649|T037|AB|808.59|ICD9CM|Pelvic fracture NEC-open|Pelvic fracture NEC-open
C0272576|T037|PT|808.8|ICD9CM|Closed unspecified fracture of pelvis|Closed unspecified fracture of pelvis
C0272576|T037|AB|808.8|ICD9CM|Pelvic fracture NOS-clos|Pelvic fracture NOS-clos
C0272577|T037|PT|808.9|ICD9CM|Open unspecified fracture of pelvis|Open unspecified fracture of pelvis
C0272577|T037|AB|808.9|ICD9CM|Pelvic fracture NOS-open|Pelvic fracture NOS-open
C0159655|T037|HT|809|ICD9CM|Ill-defined fractures of bones of trunk|Ill-defined fractures of bones of trunk
C0159656|T037|PT|809.0|ICD9CM|Fracture of bones of trunk, closed|Fracture of bones of trunk, closed
C0159656|T037|AB|809.0|ICD9CM|Fracture trunk bone-clos|Fracture trunk bone-clos
C0159657|T037|PT|809.1|ICD9CM|Fracture of bones of trunk, open|Fracture of bones of trunk, open
C0159657|T037|AB|809.1|ICD9CM|Fracture trunk bone-open|Fracture trunk bone-open
C0159658|T037|HT|810|ICD9CM|Fracture of clavicle|Fracture of clavicle
C0178316|T037|HT|810-819.99|ICD9CM|FRACTURE OF UPPER LIMB|FRACTURE OF UPPER LIMB
C0159659|T037|HT|810.0|ICD9CM|Closed fracture of clavicle|Closed fracture of clavicle
C0159659|T037|PT|810.00|ICD9CM|Closed fracture of clavicle, unspecified part|Closed fracture of clavicle, unspecified part
C0159659|T037|AB|810.00|ICD9CM|Fx clavicle NOS-closed|Fx clavicle NOS-closed
C0435521|T037|PT|810.01|ICD9CM|Closed fracture of sternal end of clavicle|Closed fracture of sternal end of clavicle
C0435521|T037|AB|810.01|ICD9CM|Fx clavicl, stern end-cl|Fx clavicl, stern end-cl
C0159661|T037|PT|810.02|ICD9CM|Closed fracture of shaft of clavicle|Closed fracture of shaft of clavicle
C0159661|T037|AB|810.02|ICD9CM|Fx clavicle shaft-closed|Fx clavicle shaft-closed
C0435522|T037|PT|810.03|ICD9CM|Closed fracture of acromial end of clavicle|Closed fracture of acromial end of clavicle
C0435522|T037|AB|810.03|ICD9CM|Fx clavicl, acrom end-cl|Fx clavicl, acrom end-cl
C0159663|T037|HT|810.1|ICD9CM|Open fracture of clavicle|Open fracture of clavicle
C0159663|T037|AB|810.10|ICD9CM|Fx clavicle NOS-open|Fx clavicle NOS-open
C0159663|T037|PT|810.10|ICD9CM|Open fracture of clavicle, unspecified part|Open fracture of clavicle, unspecified part
C0435523|T037|AB|810.11|ICD9CM|Fx clavic, stern end-opn|Fx clavic, stern end-opn
C0435523|T037|PT|810.11|ICD9CM|Open fracture of sternal end of clavicle|Open fracture of sternal end of clavicle
C0159665|T037|AB|810.12|ICD9CM|Fx clavicle shaft-open|Fx clavicle shaft-open
C0159665|T037|PT|810.12|ICD9CM|Open fracture of shaft of clavicle|Open fracture of shaft of clavicle
C0435524|T037|AB|810.13|ICD9CM|Fx clavic, acrom end-opn|Fx clavic, acrom end-opn
C0435524|T037|PT|810.13|ICD9CM|Open fracture of acromial end of clavicle|Open fracture of acromial end of clavicle
C0159667|T037|HT|811|ICD9CM|Fracture of scapula|Fracture of scapula
C0159668|T037|HT|811.0|ICD9CM|Closed fracture of scapula|Closed fracture of scapula
C0159668|T037|PT|811.00|ICD9CM|Closed fracture of scapula, unspecified part|Closed fracture of scapula, unspecified part
C0159668|T037|AB|811.00|ICD9CM|Fx scapula NOS-closed|Fx scapula NOS-closed
C0159669|T037|PT|811.01|ICD9CM|Closed fracture of acromial process of scapula|Closed fracture of acromial process of scapula
C0159669|T037|AB|811.01|ICD9CM|Fx scapul, acrom proc-cl|Fx scapul, acrom proc-cl
C0435525|T037|PT|811.02|ICD9CM|Closed fracture of coracoid process of scapula|Closed fracture of coracoid process of scapula
C0435525|T037|AB|811.02|ICD9CM|Fx scapul, corac proc-cl|Fx scapul, corac proc-cl
C0159671|T037|PT|811.03|ICD9CM|Closed fracture of glenoid cavity and neck of scapula|Closed fracture of glenoid cavity and neck of scapula
C0159671|T037|AB|811.03|ICD9CM|Fx scap, glen cav/nck-cl|Fx scap, glen cav/nck-cl
C0159672|T037|PT|811.09|ICD9CM|Closed fracture of scapula, other|Closed fracture of scapula, other
C0159672|T037|AB|811.09|ICD9CM|Fx scapula NEC-closed|Fx scapula NEC-closed
C0159673|T037|HT|811.1|ICD9CM|Open fracture of scapula|Open fracture of scapula
C0159673|T037|AB|811.10|ICD9CM|Fx scapula NOS-open|Fx scapula NOS-open
C0159673|T037|PT|811.10|ICD9CM|Open fracture of scapula, unspecified part|Open fracture of scapula, unspecified part
C0159674|T037|AB|811.11|ICD9CM|Fx scapul, acrom proc-op|Fx scapul, acrom proc-op
C0159674|T037|PT|811.11|ICD9CM|Open fracture of acromial process of scapula|Open fracture of acromial process of scapula
C0159675|T037|AB|811.12|ICD9CM|Fx scapul, corac proc-op|Fx scapul, corac proc-op
C0159675|T037|PT|811.12|ICD9CM|Open fracture of coracoid process|Open fracture of coracoid process
C1306154|T037|AB|811.13|ICD9CM|Fx scap, glen cav/nck-op|Fx scap, glen cav/nck-op
C1306154|T037|PT|811.13|ICD9CM|Open fracture of glenoid cavity and neck of scapula|Open fracture of glenoid cavity and neck of scapula
C0159677|T037|AB|811.19|ICD9CM|Fx scapula NEC-open|Fx scapula NEC-open
C0159677|T037|PT|811.19|ICD9CM|Open fracture of scapula, other|Open fracture of scapula, other
C0020162|T037|HT|812|ICD9CM|Fracture of humerus|Fracture of humerus
C0159678|T037|HT|812.0|ICD9CM|Fracture of upper end of humerus, closed|Fracture of upper end of humerus, closed
C0159679|T037|PT|812.00|ICD9CM|Closed fracture of unspecified part of upper end of humerus|Closed fracture of unspecified part of upper end of humerus
C0159679|T037|AB|812.00|ICD9CM|Fx up end humerus NOS-cl|Fx up end humerus NOS-cl
C0159680|T037|PT|812.01|ICD9CM|Closed fracture of surgical neck of humerus|Closed fracture of surgical neck of humerus
C0159680|T037|AB|812.01|ICD9CM|Fx surg nck humerus-clos|Fx surg nck humerus-clos
C0435532|T037|PT|812.02|ICD9CM|Closed fracture of anatomical neck of humerus|Closed fracture of anatomical neck of humerus
C0435532|T037|AB|812.02|ICD9CM|Fx anatom nck humerus-cl|Fx anatom nck humerus-cl
C0435533|T037|PT|812.03|ICD9CM|Closed fracture of greater tuberosity of humerus|Closed fracture of greater tuberosity of humerus
C0435533|T037|AB|812.03|ICD9CM|Fx gr tuberos humerus-cl|Fx gr tuberos humerus-cl
C0159683|T037|AB|812.09|ICD9CM|Fx upper humerus NEC-cl|Fx upper humerus NEC-cl
C0159683|T037|PT|812.09|ICD9CM|Other closed fracture of upper end of humerus|Other closed fracture of upper end of humerus
C0159684|T037|HT|812.1|ICD9CM|Fracture of upper end of humerus, open|Fracture of upper end of humerus, open
C0159685|T037|AB|812.10|ICD9CM|Fx upper humerus NOS-opn|Fx upper humerus NOS-opn
C0159685|T037|PT|812.10|ICD9CM|Open fracture of unspecified part of upper end of humerus|Open fracture of unspecified part of upper end of humerus
C0159686|T037|AB|812.11|ICD9CM|Fx surg neck humerus-opn|Fx surg neck humerus-opn
C0159686|T037|PT|812.11|ICD9CM|Open fracture of surgical neck of humerus|Open fracture of surgical neck of humerus
C0435539|T037|AB|812.12|ICD9CM|Fx anat neck humerus-opn|Fx anat neck humerus-opn
C0435539|T037|PT|812.12|ICD9CM|Open fracture of anatomical neck of humerus|Open fracture of anatomical neck of humerus
C0435540|T037|AB|812.13|ICD9CM|Fx gr tuberos humer-open|Fx gr tuberos humer-open
C0435540|T037|PT|812.13|ICD9CM|Open fracture of greater tuberosity of humerus|Open fracture of greater tuberosity of humerus
C0159689|T037|AB|812.19|ICD9CM|Fx upper humerus NEC-opn|Fx upper humerus NEC-opn
C0159689|T037|PT|812.19|ICD9CM|Other open fracture of upper end of humerus|Other open fracture of upper end of humerus
C0159690|T037|HT|812.2|ICD9CM|Closed fracture of shaft or unspecified part of humerus|Closed fracture of shaft or unspecified part of humerus
C0272609|T037|PT|812.20|ICD9CM|Closed fracture of unspecified part of humerus|Closed fracture of unspecified part of humerus
C0272609|T037|AB|812.20|ICD9CM|Fx humerus NOS-closed|Fx humerus NOS-closed
C0159692|T037|PT|812.21|ICD9CM|Closed fracture of shaft of humerus|Closed fracture of shaft of humerus
C0159692|T037|AB|812.21|ICD9CM|Fx humerus shaft-closed|Fx humerus shaft-closed
C0159693|T037|HT|812.3|ICD9CM|Fracture of shaft or unspecified part of humerus, open|Fracture of shaft or unspecified part of humerus, open
C0272610|T037|AB|812.30|ICD9CM|Fx humerus NOS-open|Fx humerus NOS-open
C0272610|T037|PT|812.30|ICD9CM|Open fracture of unspecified part of humerus|Open fracture of unspecified part of humerus
C0159695|T037|AB|812.31|ICD9CM|Fx humerus shaft-open|Fx humerus shaft-open
C0159695|T037|PT|812.31|ICD9CM|Open fracture of shaft of humerus|Open fracture of shaft of humerus
C0555330|T037|HT|812.4|ICD9CM|Fracture of lower end of humerus, closed|Fracture of lower end of humerus, closed
C0555330|T037|PT|812.40|ICD9CM|Closed fracture of unspecified part of lower end of humerus|Closed fracture of unspecified part of lower end of humerus
C0555330|T037|AB|812.40|ICD9CM|Fx lower humerus NOS-cl|Fx lower humerus NOS-cl
C0435569|T037|PT|812.41|ICD9CM|Closed supracondylar fracture of humerus|Closed supracondylar fracture of humerus
C0435569|T037|AB|812.41|ICD9CM|Suprcondyl fx humerus-cl|Suprcondyl fx humerus-cl
C0435552|T037|PT|812.42|ICD9CM|Closed fracture of lateral condyle of humerus|Closed fracture of lateral condyle of humerus
C0435552|T037|AB|812.42|ICD9CM|Fx humer, lat condyl-cl|Fx humer, lat condyl-cl
C0435553|T037|PT|812.43|ICD9CM|Closed fracture of medial condyle of humerus|Closed fracture of medial condyle of humerus
C0435553|T037|AB|812.43|ICD9CM|Fx humer, med condyl-cl|Fx humer, med condyl-cl
C0159701|T037|PT|812.44|ICD9CM|Closed fracture of unspecified condyle(s) of humerus|Closed fracture of unspecified condyle(s) of humerus
C0159701|T037|AB|812.44|ICD9CM|Fx humer, condyl NOS-cl|Fx humer, condyl NOS-cl
C0159702|T037|AB|812.49|ICD9CM|Fx lower humerus NEC-cl|Fx lower humerus NEC-cl
C0159702|T037|PT|812.49|ICD9CM|Other closed fracture of lower end of humerus|Other closed fracture of lower end of humerus
C0555332|T037|HT|812.5|ICD9CM|Fracture of lower end of humerus, open|Fracture of lower end of humerus, open
C0555332|T037|AB|812.50|ICD9CM|Fx lower humer NOS-open|Fx lower humer NOS-open
C0555332|T037|PT|812.50|ICD9CM|Open fracture of unspecified part of lower end of humerus|Open fracture of unspecified part of lower end of humerus
C0435570|T037|PT|812.51|ICD9CM|Open supracondylar fracture of humerus|Open supracondylar fracture of humerus
C0435570|T037|AB|812.51|ICD9CM|Supracondyl fx humer-opn|Supracondyl fx humer-opn
C0435563|T037|AB|812.52|ICD9CM|Fx humer, lat condyl-opn|Fx humer, lat condyl-opn
C0435563|T037|PT|812.52|ICD9CM|Open fracture of lateral condyle of humerus|Open fracture of lateral condyle of humerus
C0435564|T037|AB|812.53|ICD9CM|Fx humer, med condyl-opn|Fx humer, med condyl-opn
C0435564|T037|PT|812.53|ICD9CM|Open fracture of medial condyle of humerus|Open fracture of medial condyle of humerus
C0159708|T037|AB|812.54|ICD9CM|Fx humer, condyl NOS-opn|Fx humer, condyl NOS-opn
C0159708|T037|PT|812.54|ICD9CM|Open fracture of unspecified condyle(s) of humerus|Open fracture of unspecified condyle(s) of humerus
C0159709|T037|AB|812.59|ICD9CM|Fx lower humer NEC-open|Fx lower humer NEC-open
C0159709|T037|PT|812.59|ICD9CM|Other open fracture of lower end of humerus|Other open fracture of lower end of humerus
C0159710|T037|HT|813|ICD9CM|Fracture of radius and ulna|Fracture of radius and ulna
C0435623|T037|HT|813.0|ICD9CM|Fracture of upper end of radius and ulna, closed|Fracture of upper end of radius and ulna, closed
C0375623|T037|PT|813.00|ICD9CM|Closed fracture of upper end of forearm, unspecified|Closed fracture of upper end of forearm, unspecified
C0375623|T037|AB|813.00|ICD9CM|Fx upper forearm NOS-cl|Fx upper forearm NOS-cl
C0159713|T037|PT|813.01|ICD9CM|Closed fracture of olecranon process of ulna|Closed fracture of olecranon process of ulna
C0159713|T037|AB|813.01|ICD9CM|Fx olecran proc ulna-cl|Fx olecran proc ulna-cl
C0435603|T037|PT|813.02|ICD9CM|Closed fracture of coronoid process of ulna|Closed fracture of coronoid process of ulna
C0435603|T037|AB|813.02|ICD9CM|Fx coronoid proc ulna-cl|Fx coronoid proc ulna-cl
C0026509|T037|PT|813.03|ICD9CM|Closed Monteggia's fracture|Closed Monteggia's fracture
C0026509|T037|AB|813.03|ICD9CM|Monteggia's fx-closed|Monteggia's fx-closed
C0159715|T037|AB|813.04|ICD9CM|Fx upper ulna NEC/NOS-cl|Fx upper ulna NEC/NOS-cl
C0159715|T037|PT|813.04|ICD9CM|Other and unspecified closed fractures of proximal end of ulna (alone)|Other and unspecified closed fractures of proximal end of ulna (alone)
C0159716|T037|PT|813.05|ICD9CM|Closed fracture of head of radius|Closed fracture of head of radius
C0159716|T037|AB|813.05|ICD9CM|Fx radius head-closed|Fx radius head-closed
C0159717|T037|PT|813.06|ICD9CM|Closed fracture of neck of radius|Closed fracture of neck of radius
C0159717|T037|AB|813.06|ICD9CM|Fx radius neck-closed|Fx radius neck-closed
C0159718|T037|AB|813.07|ICD9CM|Fx up radius NEC/NOS-cl|Fx up radius NEC/NOS-cl
C0159718|T037|PT|813.07|ICD9CM|Other and unspecified closed fractures of proximal end of radius (alone)|Other and unspecified closed fractures of proximal end of radius (alone)
C0435623|T037|PT|813.08|ICD9CM|Closed fracture of radius with ulna, upper end [any part]|Closed fracture of radius with ulna, upper end [any part]
C0435623|T037|AB|813.08|ICD9CM|Fx up radius w ulna-clos|Fx up radius w ulna-clos
C0159720|T037|HT|813.1|ICD9CM|Fracture of upper end of radius and ulna, open|Fracture of upper end of radius and ulna, open
C0375624|T037|AB|813.10|ICD9CM|Fx upper forearm NOS-opn|Fx upper forearm NOS-opn
C0375624|T037|PT|813.10|ICD9CM|Open fracture of upper end of forearm, unspecified|Open fracture of upper end of forearm, unspecified
C0159722|T037|AB|813.11|ICD9CM|Fx olecran proc ulna-opn|Fx olecran proc ulna-opn
C0159722|T037|PT|813.11|ICD9CM|Open fracture of olecranon process of ulna|Open fracture of olecranon process of ulna
C0159723|T037|AB|813.12|ICD9CM|Fx coronoid pro ulna-opn|Fx coronoid pro ulna-opn
C0159723|T037|PT|813.12|ICD9CM|Open fracture of coronoid process of ulna|Open fracture of coronoid process of ulna
C0159724|T037|AB|813.13|ICD9CM|Monteggia's fx-open|Monteggia's fx-open
C0159724|T037|PT|813.13|ICD9CM|Open Monteggia's fracture|Open Monteggia's fracture
C0159725|T037|AB|813.14|ICD9CM|Fx up ulna NEC/NOS-open|Fx up ulna NEC/NOS-open
C0159725|T037|PT|813.14|ICD9CM|Other and unspecified open fractures of proximal end of ulna (alone)|Other and unspecified open fractures of proximal end of ulna (alone)
C0159726|T037|AB|813.15|ICD9CM|Fx radius head-open|Fx radius head-open
C0159726|T037|PT|813.15|ICD9CM|Open fracture of head of radius|Open fracture of head of radius
C0159727|T037|AB|813.16|ICD9CM|Fx radius neck-open|Fx radius neck-open
C0159727|T037|PT|813.16|ICD9CM|Open fracture of neck of radius|Open fracture of neck of radius
C0159728|T037|AB|813.17|ICD9CM|Fx up radius NEC/NOS-opn|Fx up radius NEC/NOS-opn
C0159728|T037|PT|813.17|ICD9CM|Other and unspecified open fractures of proximal end of radius (alone)|Other and unspecified open fractures of proximal end of radius (alone)
C0159720|T037|AB|813.18|ICD9CM|Fx up radius w ulna-open|Fx up radius w ulna-open
C0159720|T037|PT|813.18|ICD9CM|Open fracture of radius with ulna, upper end (any part)|Open fracture of radius with ulna, upper end (any part)
C0159730|T037|HT|813.2|ICD9CM|Fracture of shaft of radius and ulna, closed|Fracture of shaft of radius and ulna, closed
C0159731|T037|PT|813.20|ICD9CM|Closed fracture of shaft of radius or ulna, unspecified|Closed fracture of shaft of radius or ulna, unspecified
C0159731|T037|AB|813.20|ICD9CM|Fx shaft forearm NOS-cl|Fx shaft forearm NOS-cl
C0272638|T037|PT|813.21|ICD9CM|Closed fracture of shaft of radius (alone)|Closed fracture of shaft of radius (alone)
C0272638|T037|AB|813.21|ICD9CM|Fx radius shaft-closed|Fx radius shaft-closed
C0159733|T037|PT|813.22|ICD9CM|Closed fracture of shaft of ulna (alone)|Closed fracture of shaft of ulna (alone)
C0159733|T037|AB|813.22|ICD9CM|Fx ulna shaft-closed|Fx ulna shaft-closed
C0159730|T037|PT|813.23|ICD9CM|Closed fracture of shaft of radius with ulna|Closed fracture of shaft of radius with ulna
C0159730|T037|AB|813.23|ICD9CM|Fx shaft rad w ulna-clos|Fx shaft rad w ulna-clos
C0159734|T037|HT|813.3|ICD9CM|Fracture of shaft of radius and ulna, open|Fracture of shaft of radius and ulna, open
C0159735|T037|AB|813.30|ICD9CM|Fx shaft forearm NOS-opn|Fx shaft forearm NOS-opn
C0159735|T037|PT|813.30|ICD9CM|Open fracture of shaft of radius or ulna, unspecified|Open fracture of shaft of radius or ulna, unspecified
C0272641|T037|AB|813.31|ICD9CM|Fx radius shaft-open|Fx radius shaft-open
C0272641|T037|PT|813.31|ICD9CM|Open fracture of shaft of radius (alone)|Open fracture of shaft of radius (alone)
C0159737|T037|AB|813.32|ICD9CM|Fx ulna shaft-open|Fx ulna shaft-open
C0159737|T037|PT|813.32|ICD9CM|Open fracture of shaft of ulna (alone)|Open fracture of shaft of ulna (alone)
C0159734|T037|AB|813.33|ICD9CM|Fx shaft rad w ulna-open|Fx shaft rad w ulna-open
C0159734|T037|PT|813.33|ICD9CM|Open fracture of shaft of radius with ulna|Open fracture of shaft of radius with ulna
C0159738|T037|HT|813.4|ICD9CM|Fracture of lower end of radius and ulna, closed|Fracture of lower end of radius and ulna, closed
C0159739|T037|PT|813.40|ICD9CM|Closed fracture of lower end of forearm, unspecified|Closed fracture of lower end of forearm, unspecified
C0159739|T037|AB|813.40|ICD9CM|Fx lower forearm NOS-cl|Fx lower forearm NOS-cl
C0009354|T037|PT|813.41|ICD9CM|Closed Colles' fracture|Closed Colles' fracture
C0009354|T037|AB|813.41|ICD9CM|Colles' fracture-closed|Colles' fracture-closed
C0159740|T037|AB|813.42|ICD9CM|Fx distal radius NEC-cl|Fx distal radius NEC-cl
C0159740|T037|PT|813.42|ICD9CM|Other closed fractures of distal end of radius (alone)|Other closed fractures of distal end of radius (alone)
C0272647|T037|PT|813.43|ICD9CM|Closed fracture of distal end of ulna (alone)|Closed fracture of distal end of ulna (alone)
C0272647|T037|AB|813.43|ICD9CM|Fx distal ulna-closed|Fx distal ulna-closed
C0159738|T037|PT|813.44|ICD9CM|Closed fracture of lower end of radius with ulna|Closed fracture of lower end of radius with ulna
C0159738|T037|AB|813.44|ICD9CM|Fx low radius w ulna-cl|Fx low radius w ulna-cl
C2712371|T037|PT|813.45|ICD9CM|Torus fracture of radius (alone)|Torus fracture of radius (alone)
C2712371|T037|AB|813.45|ICD9CM|Torus fx radius-cl/alone|Torus fx radius-cl/alone
C2712372|T037|PT|813.46|ICD9CM|Torus fracture of ulna (alone)|Torus fracture of ulna (alone)
C2712372|T037|AB|813.46|ICD9CM|Torus fx ulna-closed|Torus fx ulna-closed
C2712373|T037|PT|813.47|ICD9CM|Torus fracture of radius and ulna|Torus fracture of radius and ulna
C2712373|T037|AB|813.47|ICD9CM|Torus fx radius/ulna-clo|Torus fx radius/ulna-clo
C0159742|T037|HT|813.5|ICD9CM|Fracture of lower end of radius and ulna, open|Fracture of lower end of radius and ulna, open
C0159743|T037|AB|813.50|ICD9CM|Fx lower forearm NOS-opn|Fx lower forearm NOS-opn
C0159743|T037|PT|813.50|ICD9CM|Open fracture of lower end of forearm, unspecified|Open fracture of lower end of forearm, unspecified
C0159744|T037|AB|813.51|ICD9CM|Colles' fracture-open|Colles' fracture-open
C0159744|T037|PT|813.51|ICD9CM|Open Colles' fracture|Open Colles' fracture
C0159745|T037|AB|813.52|ICD9CM|Fx distal radius NEC-opn|Fx distal radius NEC-opn
C0159745|T037|PT|813.52|ICD9CM|Other open fractures of distal end of radius (alone)|Other open fractures of distal end of radius (alone)
C0159746|T037|AB|813.53|ICD9CM|Fx distal ulna-open|Fx distal ulna-open
C0159746|T037|PT|813.53|ICD9CM|Open fracture of distal end of ulna (alone)|Open fracture of distal end of ulna (alone)
C0159742|T037|AB|813.54|ICD9CM|Fx low radius w ulna-opn|Fx low radius w ulna-opn
C0159742|T037|PT|813.54|ICD9CM|Open fracture of lower end of radius with ulna|Open fracture of lower end of radius with ulna
C0159747|T037|HT|813.8|ICD9CM|Fracture of unspecified part of radius with ulna, closed|Fracture of unspecified part of radius with ulna, closed
C0159748|T037|PT|813.80|ICD9CM|Closed fracture of unspecified part of forearm|Closed fracture of unspecified part of forearm
C0159748|T037|AB|813.80|ICD9CM|Fx forearm NOS-closed|Fx forearm NOS-closed
C0016652|T037|PT|813.81|ICD9CM|Closed fracture of unspecified part of radius (alone)|Closed fracture of unspecified part of radius (alone)
C0016652|T037|AB|813.81|ICD9CM|Fx radius NOS-closed|Fx radius NOS-closed
C0016653|T037|PT|813.82|ICD9CM|Closed fracture of unspecified part of ulna (alone)|Closed fracture of unspecified part of ulna (alone)
C0016653|T037|AB|813.82|ICD9CM|Fracture ulna NOS-closed|Fracture ulna NOS-closed
C0159747|T037|PT|813.83|ICD9CM|Closed fracture of unspecified part of radius with ulna|Closed fracture of unspecified part of radius with ulna
C0159747|T037|AB|813.83|ICD9CM|Fx radius w ulna NOS-cl|Fx radius w ulna NOS-cl
C0159749|T037|HT|813.9|ICD9CM|Fracture of unspecified part of radius with ulna, open|Fracture of unspecified part of radius with ulna, open
C0159750|T037|AB|813.90|ICD9CM|Fx forearm NOS-open|Fx forearm NOS-open
C0159750|T037|PT|813.90|ICD9CM|Open fracture of unspecified part of forearm|Open fracture of unspecified part of forearm
C0159751|T037|AB|813.91|ICD9CM|Fracture radius NOS-open|Fracture radius NOS-open
C0159751|T037|PT|813.91|ICD9CM|Open fracture of unspecified part of radius (alone)|Open fracture of unspecified part of radius (alone)
C0159752|T037|AB|813.92|ICD9CM|Fracture ulna NOS-open|Fracture ulna NOS-open
C0159752|T037|PT|813.92|ICD9CM|Open fracture of unspecified part of ulna (alone)|Open fracture of unspecified part of ulna (alone)
C0159749|T037|AB|813.93|ICD9CM|Fx radius w ulna NOS-opn|Fx radius w ulna NOS-opn
C0159749|T037|PT|813.93|ICD9CM|Open fracture of unspecified part of radius with ulna|Open fracture of unspecified part of radius with ulna
C0016644|T037|HT|814|ICD9CM|Fracture of carpal bone(s)|Fracture of carpal bone(s)
C0009044|T037|HT|814.0|ICD9CM|Closed fractures of carpal bones|Closed fractures of carpal bones
C0009044|T037|PT|814.00|ICD9CM|Closed fracture of carpal bone, unspecified|Closed fracture of carpal bone, unspecified
C0009044|T037|AB|814.00|ICD9CM|Fx carpal bone NOS-close|Fx carpal bone NOS-close
C0435644|T037|PT|814.01|ICD9CM|Closed fracture of navicular [scaphoid] bone of wrist|Closed fracture of navicular [scaphoid] bone of wrist
C0435644|T037|AB|814.01|ICD9CM|Fx navicular, wrist-clos|Fx navicular, wrist-clos
C0435633|T037|PT|814.02|ICD9CM|Closed fracture of lunate [semilunar] bone of wrist|Closed fracture of lunate [semilunar] bone of wrist
C0435633|T037|AB|814.02|ICD9CM|Fx lunate, wrist-closed|Fx lunate, wrist-closed
C0272665|T037|PT|814.03|ICD9CM|Closed fracture of triquetral [cuneiform] bone of wrist|Closed fracture of triquetral [cuneiform] bone of wrist
C0272665|T037|AB|814.03|ICD9CM|Fx triquetral, wrist-cl|Fx triquetral, wrist-cl
C0159758|T037|PT|814.04|ICD9CM|Closed fracture of pisiform bone of wrist|Closed fracture of pisiform bone of wrist
C0159758|T037|AB|814.04|ICD9CM|Fx pisiform-closed|Fx pisiform-closed
C0272666|T037|PT|814.05|ICD9CM|Closed fracture of trapezium bone [larger multangular] of wrist|Closed fracture of trapezium bone [larger multangular] of wrist
C0272666|T037|AB|814.05|ICD9CM|Fx trapezium bone-closed|Fx trapezium bone-closed
C0435634|T037|PT|814.06|ICD9CM|Closed fracture of trapezoid bone [smaller multangular] of wrist|Closed fracture of trapezoid bone [smaller multangular] of wrist
C0435634|T037|AB|814.06|ICD9CM|Fx trapezoid bone-closed|Fx trapezoid bone-closed
C0272668|T037|PT|814.07|ICD9CM|Closed fracture of capitate bone [os magnum] of wrist|Closed fracture of capitate bone [os magnum] of wrist
C0272668|T037|AB|814.07|ICD9CM|Fx capitate bone-closed|Fx capitate bone-closed
C0272669|T037|PT|814.08|ICD9CM|Closed fracture of hamate [unciform] bone of wrist|Closed fracture of hamate [unciform] bone of wrist
C0272669|T037|AB|814.08|ICD9CM|Fx hamate bone-closed|Fx hamate bone-closed
C0159763|T037|PT|814.09|ICD9CM|Closed fracture of other bone of wrist|Closed fracture of other bone of wrist
C0159763|T037|AB|814.09|ICD9CM|Fx carpal bone NEC-close|Fx carpal bone NEC-close
C0159765|T037|HT|814.1|ICD9CM|Open fractures of carpal bones|Open fractures of carpal bones
C0159765|T037|AB|814.10|ICD9CM|Fx carpal bone NOS-open|Fx carpal bone NOS-open
C0159765|T037|PT|814.10|ICD9CM|Open fracture of carpal bone, unspecified|Open fracture of carpal bone, unspecified
C0435650|T037|AB|814.11|ICD9CM|Fx navicular, wrist-open|Fx navicular, wrist-open
C0435650|T037|PT|814.11|ICD9CM|Open fracture of navicular [scaphoid] bone of wrist|Open fracture of navicular [scaphoid] bone of wrist
C0435638|T037|AB|814.12|ICD9CM|Fx lunate, wrist-open|Fx lunate, wrist-open
C0435638|T037|PT|814.12|ICD9CM|Open fracture of lunate [semilunar] bone of wrist|Open fracture of lunate [semilunar] bone of wrist
C0272672|T037|AB|814.13|ICD9CM|Fx triquetral, wrist-opn|Fx triquetral, wrist-opn
C0272672|T037|PT|814.13|ICD9CM|Open fracture of triquetral [cuneiform] bone of wrist|Open fracture of triquetral [cuneiform] bone of wrist
C0159769|T037|AB|814.14|ICD9CM|Fx pisiform-open|Fx pisiform-open
C0159769|T037|PT|814.14|ICD9CM|Open fracture of pisiform bone of wrist|Open fracture of pisiform bone of wrist
C0272673|T037|AB|814.15|ICD9CM|Fx trapezium bone-open|Fx trapezium bone-open
C0272673|T037|PT|814.15|ICD9CM|Open fracture of trapezium bone [larger multangular] of wrist|Open fracture of trapezium bone [larger multangular] of wrist
C0435639|T037|AB|814.16|ICD9CM|Fx trapezoid bone-open|Fx trapezoid bone-open
C0435639|T037|PT|814.16|ICD9CM|Open fracture of trapezoid bone [smaller multangular] of wrist|Open fracture of trapezoid bone [smaller multangular] of wrist
C0272675|T037|AB|814.17|ICD9CM|Fx capitate bone-open|Fx capitate bone-open
C0272675|T037|PT|814.17|ICD9CM|Open fracture of capitate bone [os magnum] of wrist|Open fracture of capitate bone [os magnum] of wrist
C0272676|T037|AB|814.18|ICD9CM|Fx hamate bone-open|Fx hamate bone-open
C0272676|T037|PT|814.18|ICD9CM|Open fracture of hamate [unciform] bone of wrist|Open fracture of hamate [unciform] bone of wrist
C0159774|T037|AB|814.19|ICD9CM|Fx carpal bone NEC-open|Fx carpal bone NEC-open
C0159774|T037|PT|814.19|ICD9CM|Open fracture of other bone of wrist|Open fracture of other bone of wrist
C0272677|T037|HT|815|ICD9CM|Fracture of metacarpal bone(s)|Fracture of metacarpal bone(s)
C0159776|T037|HT|815.0|ICD9CM|Closed fracture of metacarpal bones|Closed fracture of metacarpal bones
C0159776|T037|PT|815.00|ICD9CM|Closed fracture of metacarpal bone(s), site unspecified|Closed fracture of metacarpal bone(s), site unspecified
C0159776|T037|AB|815.00|ICD9CM|Fx metacarpal NOS-closed|Fx metacarpal NOS-closed
C0272684|T037|PT|815.01|ICD9CM|Closed fracture of base of thumb [first] metacarpal|Closed fracture of base of thumb [first] metacarpal
C0272684|T037|AB|815.01|ICD9CM|Fx 1st metacarp base-cl|Fx 1st metacarp base-cl
C0272686|T037|PT|815.02|ICD9CM|Closed fracture of base of other metacarpal bone(s)|Closed fracture of base of other metacarpal bone(s)
C0272686|T037|AB|815.02|ICD9CM|Fx metacarp base NEC-cl|Fx metacarp base NEC-cl
C0272687|T037|PT|815.03|ICD9CM|Closed fracture of shaft of metacarpal bone(s)|Closed fracture of shaft of metacarpal bone(s)
C0272687|T037|AB|815.03|ICD9CM|Fx metacarpal shaft-clos|Fx metacarpal shaft-clos
C0272688|T037|PT|815.04|ICD9CM|Closed fracture of neck of metacarpal bone(s)|Closed fracture of neck of metacarpal bone(s)
C0272688|T037|AB|815.04|ICD9CM|Fx metacarpal neck-close|Fx metacarpal neck-close
C0435669|T037|PT|815.09|ICD9CM|Closed fracture of multiple sites of metacarpus|Closed fracture of multiple sites of metacarpus
C0435669|T037|AB|815.09|ICD9CM|Mult fx metacarpus-close|Mult fx metacarpus-close
C0159783|T037|HT|815.1|ICD9CM|Open fracture of metacarpal bones|Open fracture of metacarpal bones
C0159783|T037|AB|815.10|ICD9CM|Fx metacarpal NOS-open|Fx metacarpal NOS-open
C0159783|T037|PT|815.10|ICD9CM|Open fracture of metacarpal bone(s), site unspecified|Open fracture of metacarpal bone(s), site unspecified
C0272689|T037|AB|815.11|ICD9CM|Fx 1st metacarp base-opn|Fx 1st metacarp base-opn
C0272689|T037|PT|815.11|ICD9CM|Open fracture of base of thumb [first] metacarpal|Open fracture of base of thumb [first] metacarpal
C0272691|T037|AB|815.12|ICD9CM|Fx metacarp base NEC-opn|Fx metacarp base NEC-opn
C0272691|T037|PT|815.12|ICD9CM|Open fracture of base of other metacarpal bone(s)|Open fracture of base of other metacarpal bone(s)
C0272692|T037|AB|815.13|ICD9CM|Fx metacarpal shaft-open|Fx metacarpal shaft-open
C0272692|T037|PT|815.13|ICD9CM|Open fracture of shaft of metacarpal bone(s)|Open fracture of shaft of metacarpal bone(s)
C0272693|T037|AB|815.14|ICD9CM|Fx metacarpal neck-open|Fx metacarpal neck-open
C0272693|T037|PT|815.14|ICD9CM|Open fracture of neck of metacarpal bone(s)|Open fracture of neck of metacarpal bone(s)
C0435656|T037|AB|815.19|ICD9CM|Mult fx metacarpus-open|Mult fx metacarpus-open
C0435656|T037|PT|815.19|ICD9CM|Open fracture of multiple sites of metacarpus|Open fracture of multiple sites of metacarpus
C0159790|T037|HT|816|ICD9CM|Fracture of one or more phalanges of hand|Fracture of one or more phalanges of hand
C0159791|T037|HT|816.0|ICD9CM|Closed fracture of one or more phalanges of hand|Closed fracture of one or more phalanges of hand
C0159791|T037|PT|816.00|ICD9CM|Closed fracture of phalanx or phalanges of hand, unspecified|Closed fracture of phalanx or phalanges of hand, unspecified
C0159791|T037|AB|816.00|ICD9CM|Fx phalanx, hand NOS-cl|Fx phalanx, hand NOS-cl
C0159793|T037|PT|816.01|ICD9CM|Closed fracture of middle or proximal phalanx or phalanges of hand|Closed fracture of middle or proximal phalanx or phalanges of hand
C0159793|T037|AB|816.01|ICD9CM|Fx mid/prx phal, hand-cl|Fx mid/prx phal, hand-cl
C0159794|T037|PT|816.02|ICD9CM|Closed fracture of distal phalanx or phalanges of hand|Closed fracture of distal phalanx or phalanges of hand
C0159794|T037|AB|816.02|ICD9CM|Fx dist phalanx, hand-cl|Fx dist phalanx, hand-cl
C0159795|T037|PT|816.03|ICD9CM|Closed fracture of multiple sites of phalanx or phalanges of hand|Closed fracture of multiple sites of phalanx or phalanges of hand
C0159795|T037|AB|816.03|ICD9CM|Fx mult phalan, hand-cl|Fx mult phalan, hand-cl
C0159796|T037|HT|816.1|ICD9CM|Open fracture of one or more phalanges of hand|Open fracture of one or more phalanges of hand
C0159796|T037|AB|816.10|ICD9CM|Fx phalanx, hand NOS-opn|Fx phalanx, hand NOS-opn
C0159796|T037|PT|816.10|ICD9CM|Open fracture of phalanx or phalanges of hand, unspecified|Open fracture of phalanx or phalanges of hand, unspecified
C0159798|T037|AB|816.11|ICD9CM|Fx mid/prx phal, hand-op|Fx mid/prx phal, hand-op
C0159798|T037|PT|816.11|ICD9CM|Open fracture of middle or proximal phalanx or phalanges of hand|Open fracture of middle or proximal phalanx or phalanges of hand
C0159799|T037|AB|816.12|ICD9CM|Fx distal phal, hand-opn|Fx distal phal, hand-opn
C0159799|T037|PT|816.12|ICD9CM|Open fracture of distal phalanx or phalanges of hand|Open fracture of distal phalanx or phalanges of hand
C0159800|T037|AB|816.13|ICD9CM|Fx mult phalan, hand-opn|Fx mult phalan, hand-opn
C0159800|T037|PT|816.13|ICD9CM|Open fracture of multiple sites of phalanx or phalanges of hand|Open fracture of multiple sites of phalanx or phalanges of hand
C0159801|T037|HT|817|ICD9CM|Multiple fractures of hand bones|Multiple fractures of hand bones
C0159802|T037|PT|817.0|ICD9CM|Multiple closed fractures of hand bones|Multiple closed fractures of hand bones
C0159802|T037|AB|817.0|ICD9CM|Multiple fx hand-closed|Multiple fx hand-closed
C0159803|T037|AB|817.1|ICD9CM|Multiple fx hand-open|Multiple fx hand-open
C0159803|T037|PT|817.1|ICD9CM|Multiple open fractures of hand bones|Multiple open fractures of hand bones
C0159804|T037|HT|818|ICD9CM|Ill-defined fractures of upper limb|Ill-defined fractures of upper limb
C0159805|T037|AB|818.0|ICD9CM|Fx arm mult/NOS-closed|Fx arm mult/NOS-closed
C0159805|T037|PT|818.0|ICD9CM|Ill-defined closed fractures of upper limb|Ill-defined closed fractures of upper limb
C0159806|T037|AB|818.1|ICD9CM|Fx arm mult/NOS-open|Fx arm mult/NOS-open
C0159806|T037|PT|818.1|ICD9CM|Ill-defined open fractures of upper limb|Ill-defined open fractures of upper limb
C0159807|T037|HT|819|ICD9CM|Multiple fractures involving both upper limbs, and upper limb with rib(s) and sternum|Multiple fractures involving both upper limbs, and upper limb with rib(s) and sternum
C0159808|T037|AB|819.0|ICD9CM|Fx arms w rib/sternum-cl|Fx arms w rib/sternum-cl
C0159808|T037|PT|819.0|ICD9CM|Multiple closed fractures involving both upper limbs, and upper limb with rib(s) and sternum|Multiple closed fractures involving both upper limbs, and upper limb with rib(s) and sternum
C0159809|T037|AB|819.1|ICD9CM|Fx arms w rib/stern-open|Fx arms w rib/stern-open
C0159809|T037|PT|819.1|ICD9CM|Multiple open fractures involving both upper limbs, and upper limb with rib(s) and sternum|Multiple open fractures involving both upper limbs, and upper limb with rib(s) and sternum
C0015806|T037|HT|820|ICD9CM|Fracture of neck of femur|Fracture of neck of femur
C1542178|T037|HT|820-829.99|ICD9CM|FRACTURE OF LOWER LIMB|FRACTURE OF LOWER LIMB
C0159810|T037|HT|820.0|ICD9CM|Transcervical fracture, closed|Transcervical fracture, closed
C0159811|T037|PT|820.00|ICD9CM|Closed fracture of intracapsular section of neck of femur, unspecified|Closed fracture of intracapsular section of neck of femur, unspecified
C0159811|T037|AB|820.00|ICD9CM|Fx femur intrcaps NOS-cl|Fx femur intrcaps NOS-cl
C0159812|T037|PT|820.01|ICD9CM|Closed fracture of epiphysis (separation) (upper) of neck of femur|Closed fracture of epiphysis (separation) (upper) of neck of femur
C0159812|T037|AB|820.01|ICD9CM|Fx up femur epiphy-clos|Fx up femur epiphy-clos
C0159813|T037|PT|820.02|ICD9CM|Closed fracture of midcervical section of neck of femur|Closed fracture of midcervical section of neck of femur
C0159813|T037|AB|820.02|ICD9CM|Fx femur, midcervic-clos|Fx femur, midcervic-clos
C0159814|T037|PT|820.03|ICD9CM|Closed fracture of base of neck of femur|Closed fracture of base of neck of femur
C0159814|T037|AB|820.03|ICD9CM|Fx base femoral nck-clos|Fx base femoral nck-clos
C0159815|T037|AB|820.09|ICD9CM|Fx femur intrcaps NEC-cl|Fx femur intrcaps NEC-cl
C0159815|T037|PT|820.09|ICD9CM|Other closed transcervical fracture of neck of femur|Other closed transcervical fracture of neck of femur
C0159816|T037|HT|820.1|ICD9CM|Transcervical fracture, open|Transcervical fracture, open
C0159817|T037|AB|820.10|ICD9CM|Fx femur intrcap NOS-opn|Fx femur intrcap NOS-opn
C0159817|T037|PT|820.10|ICD9CM|Open fracture of intracapsular section of neck of femur, unspecified|Open fracture of intracapsular section of neck of femur, unspecified
C0159818|T037|AB|820.11|ICD9CM|Fx up femur epiphy-open|Fx up femur epiphy-open
C0159818|T037|PT|820.11|ICD9CM|Open fracture of epiphysis (separation) (upper) of neck of femur|Open fracture of epiphysis (separation) (upper) of neck of femur
C0159819|T037|AB|820.12|ICD9CM|Fx femur, midcervic-open|Fx femur, midcervic-open
C0159819|T037|PT|820.12|ICD9CM|Open fracture of midcervical section of neck of femur|Open fracture of midcervical section of neck of femur
C0159820|T037|AB|820.13|ICD9CM|Fx base femoral nck-open|Fx base femoral nck-open
C0159820|T037|PT|820.13|ICD9CM|Open fracture of base of neck of femur|Open fracture of base of neck of femur
C0159821|T037|AB|820.19|ICD9CM|Fx femur intrcap NEC-opn|Fx femur intrcap NEC-opn
C0159821|T037|PT|820.19|ICD9CM|Other open transcervical fracture of neck of femur|Other open transcervical fracture of neck of femur
C0159822|T037|HT|820.2|ICD9CM|Pertrochanteric fracture of femur, closed|Pertrochanteric fracture of femur, closed
C0159823|T037|PT|820.20|ICD9CM|Closed fracture of trochanteric section of neck of femur|Closed fracture of trochanteric section of neck of femur
C0159823|T037|AB|820.20|ICD9CM|Trochanteric fx NOS-clos|Trochanteric fx NOS-clos
C0159824|T037|PT|820.21|ICD9CM|Closed fracture of intertrochanteric section of neck of femur|Closed fracture of intertrochanteric section of neck of femur
C0159824|T037|AB|820.21|ICD9CM|Intertrochanteric fx-cl|Intertrochanteric fx-cl
C0435830|T037|PT|820.22|ICD9CM|Closed fracture of subtrochanteric section of neck of femur|Closed fracture of subtrochanteric section of neck of femur
C0435830|T037|AB|820.22|ICD9CM|Subtrochanteric fx-close|Subtrochanteric fx-close
C0159826|T037|HT|820.3|ICD9CM|Pertrochanteric fracture of femur, open|Pertrochanteric fracture of femur, open
C0159827|T037|PT|820.30|ICD9CM|Open fracture of trochanteric section of neck of femur, unspecified|Open fracture of trochanteric section of neck of femur, unspecified
C0159827|T037|AB|820.30|ICD9CM|Trochanteric fx NOS-open|Trochanteric fx NOS-open
C0159828|T037|AB|820.31|ICD9CM|Intertrochanteric fx-opn|Intertrochanteric fx-opn
C0159828|T037|PT|820.31|ICD9CM|Open fracture of intertrochanteric section of neck of femur|Open fracture of intertrochanteric section of neck of femur
C0435834|T037|PT|820.32|ICD9CM|Open fracture of subtrochanteric section of neck of femur|Open fracture of subtrochanteric section of neck of femur
C0435834|T037|AB|820.32|ICD9CM|Subtrochanteric fx-open|Subtrochanteric fx-open
C0272751|T037|PT|820.8|ICD9CM|Closed fracture of unspecified part of neck of femur|Closed fracture of unspecified part of neck of femur
C0272751|T037|AB|820.8|ICD9CM|Fx neck of femur NOS-cl|Fx neck of femur NOS-cl
C0272752|T037|AB|820.9|ICD9CM|Fx neck of femur NOS-opn|Fx neck of femur NOS-opn
C0272752|T037|PT|820.9|ICD9CM|Open fracture of unspecified part of neck of femur|Open fracture of unspecified part of neck of femur
C0159831|T037|HT|821|ICD9CM|Fracture of other and unspecified parts of femur|Fracture of other and unspecified parts of femur
C0159832|T037|HT|821.0|ICD9CM|Fracture of shaft or unspecified part of femur, closed|Fracture of shaft or unspecified part of femur, closed
C0272729|T037|PT|821.00|ICD9CM|Closed fracture of unspecified part of femur|Closed fracture of unspecified part of femur
C0272729|T037|AB|821.00|ICD9CM|Fx femur NOS-closed|Fx femur NOS-closed
C0159833|T037|PT|821.01|ICD9CM|Closed fracture of shaft of femur|Closed fracture of shaft of femur
C0159833|T037|AB|821.01|ICD9CM|Fx femur shaft-closed|Fx femur shaft-closed
C0159834|T037|HT|821.1|ICD9CM|Fracture of shaft or unspecified part of femur, open|Fracture of shaft or unspecified part of femur, open
C0159835|T037|AB|821.10|ICD9CM|Fx femur NOS-open|Fx femur NOS-open
C0159835|T037|PT|821.10|ICD9CM|Open fracture of unspecified part of femur|Open fracture of unspecified part of femur
C0159836|T037|AB|821.11|ICD9CM|Fx femur shaft-open|Fx femur shaft-open
C0159836|T037|PT|821.11|ICD9CM|Open fracture of shaft of femur|Open fracture of shaft of femur
C0159837|T037|HT|821.2|ICD9CM|Fracture of lower end of femur, closed|Fracture of lower end of femur, closed
C0159838|T037|PT|821.20|ICD9CM|Closed fracture of lower end of femur, unspecified part|Closed fracture of lower end of femur, unspecified part
C0159838|T037|AB|821.20|ICD9CM|Fx low end femur NOS-cl|Fx low end femur NOS-cl
C0272754|T037|PT|821.21|ICD9CM|Closed fracture of condyle, femoral|Closed fracture of condyle, femoral
C0272754|T037|AB|821.21|ICD9CM|Fx femoral condyle-close|Fx femoral condyle-close
C0159840|T037|PT|821.22|ICD9CM|Closed fracture of epiphysis, lower (separation) of femur|Closed fracture of epiphysis, lower (separation) of femur
C0159840|T037|AB|821.22|ICD9CM|Fx low femur epiphy-clos|Fx low femur epiphy-clos
C0435844|T037|PT|821.23|ICD9CM|Closed supracondylar fracture of femur|Closed supracondylar fracture of femur
C0435844|T037|AB|821.23|ICD9CM|Supracondyl fx femur-cl|Supracondyl fx femur-cl
C0159842|T037|AB|821.29|ICD9CM|Fx low end femur NEC-cl|Fx low end femur NEC-cl
C0159842|T037|PT|821.29|ICD9CM|Other closed fracture of lower end of femur|Other closed fracture of lower end of femur
C0159843|T037|HT|821.3|ICD9CM|Fracture of lower end of femur, open|Fracture of lower end of femur, open
C0159844|T037|AB|821.30|ICD9CM|Fx low end femur NOS-opn|Fx low end femur NOS-opn
C0159844|T037|PT|821.30|ICD9CM|Open fracture of lower end of femur, unspecified part|Open fracture of lower end of femur, unspecified part
C0272757|T037|AB|821.31|ICD9CM|Fx femoral condyle-open|Fx femoral condyle-open
C0272757|T037|PT|821.31|ICD9CM|Open fracture of condyle, femoral|Open fracture of condyle, femoral
C0159846|T037|AB|821.32|ICD9CM|Fx low femur epiphy-open|Fx low femur epiphy-open
C0159846|T037|PT|821.32|ICD9CM|Open fracture of epiphysis. Lower (separation) of femur|Open fracture of epiphysis. Lower (separation) of femur
C0435845|T037|PT|821.33|ICD9CM|Open supracondylar fracture of femur|Open supracondylar fracture of femur
C0435845|T037|AB|821.33|ICD9CM|Supracondyl fx femur-opn|Supracondyl fx femur-opn
C0159848|T037|AB|821.39|ICD9CM|Fx low end femur NEC-opn|Fx low end femur NEC-opn
C0159848|T037|PT|821.39|ICD9CM|Other open fracture of lower end of femur|Other open fracture of lower end of femur
C0159849|T037|HT|822|ICD9CM|Fracture of patella|Fracture of patella
C0159850|T037|PT|822.0|ICD9CM|Closed fracture of patella|Closed fracture of patella
C0159850|T037|AB|822.0|ICD9CM|Fracture patella-closed|Fracture patella-closed
C0159851|T037|AB|822.1|ICD9CM|Fracture patella-open|Fracture patella-open
C0159851|T037|PT|822.1|ICD9CM|Open fracture of patella|Open fracture of patella
C0159852|T037|HT|823|ICD9CM|Fracture of tibia and fibula|Fracture of tibia and fibula
C0435903|T037|HT|823.0|ICD9CM|Fracture of upper end of tibia and fibula, closed|Fracture of upper end of tibia and fibula, closed
C0159854|T037|PT|823.00|ICD9CM|Closed fracture of upper end of tibia alone|Closed fracture of upper end of tibia alone
C0159854|T037|AB|823.00|ICD9CM|Fx upper end tibia-close|Fx upper end tibia-close
C0435898|T037|PT|823.01|ICD9CM|Closed fracture of upper end of fibula alone|Closed fracture of upper end of fibula alone
C0435898|T037|AB|823.01|ICD9CM|Fx upper end fibula-clos|Fx upper end fibula-clos
C0435903|T037|PT|823.02|ICD9CM|Closed fracture of upper end of fibula with tibia|Closed fracture of upper end of fibula with tibia
C0435903|T037|AB|823.02|ICD9CM|Fx up tibia w fibula-cl|Fx up tibia w fibula-cl
C0435905|T037|HT|823.1|ICD9CM|Fracture of upper end of tibia and fibula, open|Fracture of upper end of tibia and fibula, open
C0159858|T037|AB|823.10|ICD9CM|Fx upper end tibia-open|Fx upper end tibia-open
C0159858|T037|PT|823.10|ICD9CM|Open fracture of upper end of tibia alone|Open fracture of upper end of tibia alone
C0435876|T037|AB|823.11|ICD9CM|Fx upper end fibula-open|Fx upper end fibula-open
C0435876|T037|PT|823.11|ICD9CM|Open fracture of upper end of fibula alone|Open fracture of upper end of fibula alone
C0435905|T037|AB|823.12|ICD9CM|Fx up tibia w fibula-opn|Fx up tibia w fibula-opn
C0435905|T037|PT|823.12|ICD9CM|Open fracture of upper end of fibula with tibia|Open fracture of upper end of fibula with tibia
C0159864|T037|HT|823.2|ICD9CM|Fracture of shaft of tibia and fibula, closed|Fracture of shaft of tibia and fibula, closed
C0159862|T037|PT|823.20|ICD9CM|Closed fracture of shaft of tibia alone|Closed fracture of shaft of tibia alone
C0159862|T037|AB|823.20|ICD9CM|Fx shaft tibia-closed|Fx shaft tibia-closed
C0159863|T037|PT|823.21|ICD9CM|Closed fracture of shaft of fibula alone|Closed fracture of shaft of fibula alone
C0159863|T037|AB|823.21|ICD9CM|Fx shaft fibula-closed|Fx shaft fibula-closed
C0159864|T037|PT|823.22|ICD9CM|Closed fracture of shaft of fibula with tibia|Closed fracture of shaft of fibula with tibia
C0159864|T037|AB|823.22|ICD9CM|Fx shaft fib w tib-clos|Fx shaft fib w tib-clos
C0159868|T037|HT|823.3|ICD9CM|Fracture of shaft of tibia and fibula, open|Fracture of shaft of tibia and fibula, open
C0159866|T037|AB|823.30|ICD9CM|Fx tibia shaft-open|Fx tibia shaft-open
C0159866|T037|PT|823.30|ICD9CM|Open fracture of shaft of tibia alone|Open fracture of shaft of tibia alone
C0159867|T037|AB|823.31|ICD9CM|Fx fibula shaft-open|Fx fibula shaft-open
C0159867|T037|PT|823.31|ICD9CM|Open fracture of shaft of fibula alone|Open fracture of shaft of fibula alone
C0159868|T037|AB|823.32|ICD9CM|Fx shaft tibia w fib-opn|Fx shaft tibia w fib-opn
C0159868|T037|PT|823.32|ICD9CM|Open fracture of shaft of fibula with tibia|Open fracture of shaft of fibula with tibia
C1146542|T037|HT|823.4|ICD9CM|Torus fracture|Torus fracture
C1176359|T037|AB|823.40|ICD9CM|Torus fracture of tibia|Torus fracture of tibia
C1176359|T037|PT|823.40|ICD9CM|Torus fracture, tibia alone|Torus fracture, tibia alone
C1176360|T037|AB|823.41|ICD9CM|Torus fracture of fibula|Torus fracture of fibula
C1176360|T037|PT|823.41|ICD9CM|Torus fracture, fibula alone|Torus fracture, fibula alone
C1176361|T037|PT|823.42|ICD9CM|Torus fracture, fibula with tibia|Torus fracture, fibula with tibia
C1176361|T037|AB|823.42|ICD9CM|Torus fx tibia/fibula|Torus fx tibia/fibula
C0555347|T037|HT|823.8|ICD9CM|Fracture of unspecified part of tibia and fibula, closed|Fracture of unspecified part of tibia and fibula, closed
C0159870|T037|PT|823.80|ICD9CM|Closed fracture of unspecified part of tibia alone|Closed fracture of unspecified part of tibia alone
C0159870|T037|AB|823.80|ICD9CM|Fx tibia NOS-closed|Fx tibia NOS-closed
C0159871|T037|PT|823.81|ICD9CM|Closed fracture of unspecified part of fibula alone|Closed fracture of unspecified part of fibula alone
C0159871|T037|AB|823.81|ICD9CM|Fx fibula NOS-closed|Fx fibula NOS-closed
C0555347|T037|PT|823.82|ICD9CM|Closed fracture of unspecified part of fibula with tibia|Closed fracture of unspecified part of fibula with tibia
C0555347|T037|AB|823.82|ICD9CM|Fx tibia w fibula NOS-cl|Fx tibia w fibula NOS-cl
C0159876|T037|HT|823.9|ICD9CM|Fracture of unspecified part of tibia and fibula, open|Fracture of unspecified part of tibia and fibula, open
C0159874|T037|AB|823.90|ICD9CM|Fx tibia NOS-open|Fx tibia NOS-open
C0159874|T037|PT|823.90|ICD9CM|Open fracture of unspecified part of tibia alone|Open fracture of unspecified part of tibia alone
C0159875|T037|AB|823.91|ICD9CM|Fx fibula NOS-open|Fx fibula NOS-open
C0159875|T037|PT|823.91|ICD9CM|Open fracture of unspecified part of fibula alone|Open fracture of unspecified part of fibula alone
C0159876|T037|AB|823.92|ICD9CM|Fx tibia w fib NOS-open|Fx tibia w fib NOS-open
C0159876|T037|PT|823.92|ICD9CM|Open fracture of unspecified part of fibula with tibia|Open fracture of unspecified part of fibula with tibia
C0159877|T037|HT|824|ICD9CM|Fracture of ankle|Fracture of ankle
C0435890|T037|PT|824.0|ICD9CM|Fracture of medial malleolus, closed|Fracture of medial malleolus, closed
C0435890|T037|AB|824.0|ICD9CM|Fx medial malleolus-clos|Fx medial malleolus-clos
C0435891|T037|PT|824.1|ICD9CM|Fracture of medial malleolus, open|Fracture of medial malleolus, open
C0435891|T037|AB|824.1|ICD9CM|Fx medial malleolus-open|Fx medial malleolus-open
C0435892|T037|PT|824.2|ICD9CM|Fracture of lateral malleolus, closed|Fracture of lateral malleolus, closed
C0435892|T037|AB|824.2|ICD9CM|Fx lateral malleolus-cl|Fx lateral malleolus-cl
C0435900|T037|PT|824.3|ICD9CM|Fracture of lateral malleolus, open|Fracture of lateral malleolus, open
C0435900|T037|AB|824.3|ICD9CM|Fx lateral malleolus-opn|Fx lateral malleolus-opn
C0392611|T037|PT|824.4|ICD9CM|Bimalleolar fracture, closed|Bimalleolar fracture, closed
C0392611|T037|AB|824.4|ICD9CM|Fx bimalleolar-closed|Fx bimalleolar-closed
C0159882|T037|PT|824.5|ICD9CM|Bimalleolar fracture, open|Bimalleolar fracture, open
C0159882|T037|AB|824.5|ICD9CM|Fx bimalleolar-open|Fx bimalleolar-open
C0159883|T037|AB|824.6|ICD9CM|Fx trimalleolar-closed|Fx trimalleolar-closed
C0159883|T037|PT|824.6|ICD9CM|Trimalleolar fracture, closed|Trimalleolar fracture, closed
C0159884|T037|AB|824.7|ICD9CM|Fx trimalleolar-open|Fx trimalleolar-open
C0159884|T037|PT|824.7|ICD9CM|Trimalleolar fracture, open|Trimalleolar fracture, open
C0272769|T037|AB|824.8|ICD9CM|Fx ankle NOS-closed|Fx ankle NOS-closed
C0272769|T037|PT|824.8|ICD9CM|Unspecified fracture of ankle, closed|Unspecified fracture of ankle, closed
C0272770|T037|AB|824.9|ICD9CM|Fx ankle NOS-open|Fx ankle NOS-open
C0272770|T037|PT|824.9|ICD9CM|Unspecified fracture of ankle, open|Unspecified fracture of ankle, open
C1963546|T037|HT|825|ICD9CM|Fracture of one or more tarsal and metatarsal bones|Fracture of one or more tarsal and metatarsal bones
C0159888|T037|AB|825.0|ICD9CM|Fracture calcaneus-close|Fracture calcaneus-close
C0159888|T037|PT|825.0|ICD9CM|Fracture of calcaneus, closed|Fracture of calcaneus, closed
C0159889|T037|AB|825.1|ICD9CM|Fracture calcaneus-open|Fracture calcaneus-open
C0159889|T037|PT|825.1|ICD9CM|Fracture of calcaneus, open|Fracture of calcaneus, open
C0159890|T037|HT|825.2|ICD9CM|Fracture of other tarsal and metatarsal bones, closed|Fracture of other tarsal and metatarsal bones, closed
C0272776|T037|PT|825.20|ICD9CM|Closed fracture of unspecified bone(s) of foot [except toes]|Closed fracture of unspecified bone(s) of foot [except toes]
C0272776|T037|AB|825.20|ICD9CM|Fx foot bone NOS-closed|Fx foot bone NOS-closed
C0159892|T037|PT|825.21|ICD9CM|Closed fracture of astragalus|Closed fracture of astragalus
C0159892|T037|AB|825.21|ICD9CM|Fx astragalus-closed|Fx astragalus-closed
C0435940|T037|PT|825.22|ICD9CM|Closed fracture of navicular [scaphoid], foot|Closed fracture of navicular [scaphoid], foot
C0435940|T037|AB|825.22|ICD9CM|Fx navicular, foot-clos|Fx navicular, foot-clos
C0347815|T037|PT|825.23|ICD9CM|Closed fracture of cuboid|Closed fracture of cuboid
C0347815|T037|AB|825.23|ICD9CM|Fx cuboid-closed|Fx cuboid-closed
C0435924|T037|PT|825.24|ICD9CM|Closed fracture of cuneiform, foot|Closed fracture of cuneiform, foot
C0435924|T037|AB|825.24|ICD9CM|Fx cuneiform, foot-clos|Fx cuneiform, foot-clos
C0435944|T037|PT|825.25|ICD9CM|Closed fracture of metatarsal bone(s)|Closed fracture of metatarsal bone(s)
C0435944|T037|AB|825.25|ICD9CM|Fx metatarsal-closed|Fx metatarsal-closed
C0159890|T037|AB|825.29|ICD9CM|Fx foot bone NEC-closed|Fx foot bone NEC-closed
C0159890|T037|PT|825.29|ICD9CM|Other closed fracture of tarsal and metatarsal bones|Other closed fracture of tarsal and metatarsal bones
C0159904|T037|HT|825.3|ICD9CM|Fracture of other tarsal and metatarsal bones, open|Fracture of other tarsal and metatarsal bones, open
C0272778|T037|AB|825.30|ICD9CM|Fx foot bone NOS-open|Fx foot bone NOS-open
C0272778|T037|PT|825.30|ICD9CM|Open fracture of unspecified bone(s) of foot [except toes]|Open fracture of unspecified bone(s) of foot [except toes]
C0159899|T037|AB|825.31|ICD9CM|Fx astragalus-open|Fx astragalus-open
C0159899|T037|PT|825.31|ICD9CM|Open fracture of astragalus|Open fracture of astragalus
C0435941|T037|AB|825.32|ICD9CM|Fx navicular, foot-open|Fx navicular, foot-open
C0435941|T037|PT|825.32|ICD9CM|Open fracture of navicular [scaphoid], foot|Open fracture of navicular [scaphoid], foot
C0347816|T037|AB|825.33|ICD9CM|Fx cuboid-open|Fx cuboid-open
C0347816|T037|PT|825.33|ICD9CM|Open fracture of cuboid|Open fracture of cuboid
C0435920|T037|AB|825.34|ICD9CM|Fx cuneiform, foot-open|Fx cuneiform, foot-open
C0435920|T037|PT|825.34|ICD9CM|Open fracture of cuneiform, foot|Open fracture of cuneiform, foot
C0435950|T037|AB|825.35|ICD9CM|Fx metatarsal-open|Fx metatarsal-open
C0435950|T037|PT|825.35|ICD9CM|Open fracture of metatarsal bone(s)|Open fracture of metatarsal bone(s)
C0159904|T037|AB|825.39|ICD9CM|Fx foot bone NEC-open|Fx foot bone NEC-open
C0159904|T037|PT|825.39|ICD9CM|Other open fracture of tarsal and metatarsal bones|Other open fracture of tarsal and metatarsal bones
C0159905|T037|HT|826|ICD9CM|Fracture of one or more phalanges of foot|Fracture of one or more phalanges of foot
C0159906|T037|PT|826.0|ICD9CM|Closed fracture of one or more phalanges of foot|Closed fracture of one or more phalanges of foot
C0159906|T037|AB|826.0|ICD9CM|Fx phalanx, foot-closed|Fx phalanx, foot-closed
C0159907|T037|AB|826.1|ICD9CM|Fx phalanx, foot-open|Fx phalanx, foot-open
C0159907|T037|PT|826.1|ICD9CM|Open fracture of one or more phalanges of foot|Open fracture of one or more phalanges of foot
C0159908|T037|HT|827|ICD9CM|Other, multiple, and ill-defined fractures of lower limb|Other, multiple, and ill-defined fractures of lower limb
C0159909|T037|AB|827.0|ICD9CM|Fx lower limb NEC-closed|Fx lower limb NEC-closed
C0159909|T037|PT|827.0|ICD9CM|Other, multiple and ill-defined fractures of lower limb, closed|Other, multiple and ill-defined fractures of lower limb, closed
C0159910|T037|AB|827.1|ICD9CM|Fx lower limb NEC-open|Fx lower limb NEC-open
C0159910|T037|PT|827.1|ICD9CM|Other, multiple and ill-defined fractures of lower limb, open|Other, multiple and ill-defined fractures of lower limb, open
C0159912|T037|AB|828.0|ICD9CM|Fx legs w arm/rib-closed|Fx legs w arm/rib-closed
C0159913|T037|AB|828.1|ICD9CM|Fx legs w arm/rib-open|Fx legs w arm/rib-open
C0016658|T037|HT|829|ICD9CM|Fracture of unspecified bones|Fracture of unspecified bones
C0016659|T037|AB|829.0|ICD9CM|Fracture NOS-closed|Fracture NOS-closed
C0016659|T037|PT|829.0|ICD9CM|Fracture of unspecified bone, closed|Fracture of unspecified bone, closed
C0016662|T037|AB|829.1|ICD9CM|Fracture NOS-open|Fracture NOS-open
C0016662|T037|PT|829.1|ICD9CM|Fracture of unspecified bone, open|Fracture of unspecified bone, open
C0159914|T037|HT|830|ICD9CM|Dislocation of jaw|Dislocation of jaw
C0012691|T037|HT|830-839.99|ICD9CM|DISLOCATION|DISLOCATION
C0159915|T037|PT|830.0|ICD9CM|Closed dislocation of jaw|Closed dislocation of jaw
C0159915|T037|AB|830.0|ICD9CM|Dislocation jaw-closed|Dislocation jaw-closed
C0159916|T037|AB|830.1|ICD9CM|Dislocation jaw-open|Dislocation jaw-open
C0159916|T037|PT|830.1|ICD9CM|Open dislocation of jaw|Open dislocation of jaw
C0037005|T037|HT|831|ICD9CM|Dislocation of shoulder|Dislocation of shoulder
C0434579|T037|HT|831.0|ICD9CM|Closed dislocation of shoulder|Closed dislocation of shoulder
C0375625|T037|PT|831.00|ICD9CM|Closed dislocation of shoulder, unspecified|Closed dislocation of shoulder, unspecified
C0375625|T037|AB|831.00|ICD9CM|Disloc shoulder NOS-clos|Disloc shoulder NOS-clos
C0159917|T037|AB|831.01|ICD9CM|Ant disloc humerus-close|Ant disloc humerus-close
C0159917|T037|PT|831.01|ICD9CM|Closed anterior dislocation of humerus|Closed anterior dislocation of humerus
C0159918|T037|PT|831.02|ICD9CM|Closed posterior dislocation of humerus|Closed posterior dislocation of humerus
C0159918|T037|AB|831.02|ICD9CM|Post disloc humerus-clos|Post disloc humerus-clos
C0159919|T037|PT|831.03|ICD9CM|Closed inferior dislocation of humerus|Closed inferior dislocation of humerus
C0159919|T037|AB|831.03|ICD9CM|Infer disloc humerus-cl|Infer disloc humerus-cl
C0159920|T037|PT|831.04|ICD9CM|Closed dislocation of acromioclavicular (joint)|Closed dislocation of acromioclavicular (joint)
C0159920|T037|AB|831.04|ICD9CM|Disloc acromioclavic-cl|Disloc acromioclavic-cl
C0159921|T037|PT|831.09|ICD9CM|Closed dislocation of shoulder, other|Closed dislocation of shoulder, other
C0159921|T037|AB|831.09|ICD9CM|Disloc shoulder NEC-clos|Disloc shoulder NEC-clos
C0434583|T037|HT|831.1|ICD9CM|Open dislocation of shoulder|Open dislocation of shoulder
C0375626|T037|AB|831.10|ICD9CM|Disloc shoulder NOS-open|Disloc shoulder NOS-open
C0375626|T037|PT|831.10|ICD9CM|Open dislocation of shoulder, unspecified|Open dislocation of shoulder, unspecified
C0434585|T037|AB|831.11|ICD9CM|Ant disloc humerus-open|Ant disloc humerus-open
C0434585|T037|PT|831.11|ICD9CM|Open anterior dislocation of humerus|Open anterior dislocation of humerus
C1444204|T037|PT|831.12|ICD9CM|Open posterior dislocation of humerus|Open posterior dislocation of humerus
C1444204|T037|AB|831.12|ICD9CM|Post disloc humerus-open|Post disloc humerus-open
C0434587|T037|AB|831.13|ICD9CM|Infer disloc humerus-opn|Infer disloc humerus-opn
C0434587|T037|PT|831.13|ICD9CM|Open inferior dislocation of humerus|Open inferior dislocation of humerus
C0159926|T037|AB|831.14|ICD9CM|Disloc acromioclavic-opn|Disloc acromioclavic-opn
C0159926|T037|PT|831.14|ICD9CM|Open dislocation of acromioclavicular (joint)|Open dislocation of acromioclavicular (joint)
C0159927|T037|AB|831.19|ICD9CM|Disloc shoulder NEC-open|Disloc shoulder NEC-open
C0159927|T037|PT|831.19|ICD9CM|Open dislocation of shoulder, other|Open dislocation of shoulder, other
C2720437|T037|HT|832|ICD9CM|Dislocation of elbow|Dislocation of elbow
C0434599|T037|HT|832.0|ICD9CM|Closed dislocation of elbow|Closed dislocation of elbow
C0375627|T037|PT|832.00|ICD9CM|Closed dislocation of elbow, unspecified|Closed dislocation of elbow, unspecified
C0375627|T037|AB|832.00|ICD9CM|Dislocat elbow NOS-close|Dislocat elbow NOS-close
C0159930|T037|AB|832.01|ICD9CM|Ant disloc elbow-closed|Ant disloc elbow-closed
C0159930|T037|PT|832.01|ICD9CM|Closed anterior dislocation of elbow|Closed anterior dislocation of elbow
C0159931|T037|PT|832.02|ICD9CM|Closed posterior dislocation of elbow|Closed posterior dislocation of elbow
C0159931|T037|AB|832.02|ICD9CM|Post disloc elbow-closed|Post disloc elbow-closed
C0159932|T037|PT|832.03|ICD9CM|Closed medial dislocation of elbow|Closed medial dislocation of elbow
C0159932|T037|AB|832.03|ICD9CM|Med disloc elbow-closed|Med disloc elbow-closed
C0159933|T037|PT|832.04|ICD9CM|Closed lateral dislocation of elbow|Closed lateral dislocation of elbow
C0159933|T037|AB|832.04|ICD9CM|Lat disloc elbow-closed|Lat disloc elbow-closed
C0159934|T037|PT|832.09|ICD9CM|Closed dislocation of elbow, other|Closed dislocation of elbow, other
C0159934|T037|AB|832.09|ICD9CM|Dislocat elbow NEC-close|Dislocat elbow NEC-close
C0434608|T037|HT|832.1|ICD9CM|Open dislocation of elbow|Open dislocation of elbow
C0434608|T037|AB|832.10|ICD9CM|Dislocat elbow NOS-open|Dislocat elbow NOS-open
C0434608|T037|PT|832.10|ICD9CM|Open dislocation of elbow, unspecified|Open dislocation of elbow, unspecified
C0434601|T037|AB|832.11|ICD9CM|Ant disloc elbow-open|Ant disloc elbow-open
C0434601|T037|PT|832.11|ICD9CM|Open anterior dislocation of elbow|Open anterior dislocation of elbow
C0434602|T037|PT|832.12|ICD9CM|Open posterior dislocation of elbow|Open posterior dislocation of elbow
C0434602|T037|AB|832.12|ICD9CM|Post disloc elbow-open|Post disloc elbow-open
C0434603|T037|AB|832.13|ICD9CM|Med disloc elbow-open|Med disloc elbow-open
C0434603|T037|PT|832.13|ICD9CM|Open medial dislocation of elbow|Open medial dislocation of elbow
C0434604|T037|AB|832.14|ICD9CM|Lat dislocat elbow-open|Lat dislocat elbow-open
C0434604|T037|PT|832.14|ICD9CM|Open lateral dislocation of elbow|Open lateral dislocation of elbow
C0159940|T037|AB|832.19|ICD9CM|Dislocat elbow NEC-open|Dislocat elbow NEC-open
C0159940|T037|PT|832.19|ICD9CM|Open dislocation of elbow, other|Open dislocation of elbow, other
C0149977|T037|AB|832.2|ICD9CM|Nursemaid's elbow|Nursemaid's elbow
C0149977|T037|PT|832.2|ICD9CM|Nursemaid's elbow|Nursemaid's elbow
C0159941|T037|HT|833|ICD9CM|Dislocation of wrist|Dislocation of wrist
C0159942|T037|HT|833.0|ICD9CM|Closed dislocation of wrist|Closed dislocation of wrist
C0159942|T037|PT|833.00|ICD9CM|Closed dislocation of wrist, unspecified part|Closed dislocation of wrist, unspecified part
C0159942|T037|AB|833.00|ICD9CM|Disloc wrist NOS-closed|Disloc wrist NOS-closed
C0159943|T037|PT|833.01|ICD9CM|Closed dislocation of radioulnar (joint), distal|Closed dislocation of radioulnar (joint), distal
C0159943|T037|AB|833.01|ICD9CM|Disloc dist radiouln-cl|Disloc dist radiouln-cl
C0159944|T037|PT|833.02|ICD9CM|Closed dislocation of radiocarpal (joint)|Closed dislocation of radiocarpal (joint)
C0159944|T037|AB|833.02|ICD9CM|Disloc radiocarpal-clos|Disloc radiocarpal-clos
C0159945|T037|PT|833.03|ICD9CM|Closed dislocation of midcarpal (joint)|Closed dislocation of midcarpal (joint)
C0159945|T037|AB|833.03|ICD9CM|Disloca midcarpal-closed|Disloca midcarpal-closed
C0159946|T037|PT|833.04|ICD9CM|Closed dislocation of carpometacarpal (joint)|Closed dislocation of carpometacarpal (joint)
C0159946|T037|AB|833.04|ICD9CM|Disloc carpometacarp-cl|Disloc carpometacarp-cl
C0159947|T037|PT|833.05|ICD9CM|Closed dislocation of metacarpal (bone), proximal end|Closed dislocation of metacarpal (bone), proximal end
C0159947|T037|AB|833.05|ICD9CM|Disloc metacarpal-closed|Disloc metacarpal-closed
C0159948|T037|PT|833.09|ICD9CM|Closed dislocation of wrist, other|Closed dislocation of wrist, other
C0159948|T037|AB|833.09|ICD9CM|Disloc wrist NEC-closed|Disloc wrist NEC-closed
C0434619|T037|HT|833.1|ICD9CM|Open dislocation of wrist|Open dislocation of wrist
C0375629|T037|AB|833.10|ICD9CM|Dislocat wrist NOS-open|Dislocat wrist NOS-open
C0375629|T037|PT|833.10|ICD9CM|Open dislocation of wrist, unspecified part|Open dislocation of wrist, unspecified part
C0159950|T037|AB|833.11|ICD9CM|Disloc dist radiouln-opn|Disloc dist radiouln-opn
C0159950|T037|PT|833.11|ICD9CM|Open dislocation of radioulnar (joint), distal|Open dislocation of radioulnar (joint), distal
C0159951|T037|AB|833.12|ICD9CM|Disloc radiocarpal-open|Disloc radiocarpal-open
C0159951|T037|PT|833.12|ICD9CM|Open dislocation of radiocarpal (joint)|Open dislocation of radiocarpal (joint)
C0159952|T037|AB|833.13|ICD9CM|Dislocat midcarpal-open|Dislocat midcarpal-open
C0159952|T037|PT|833.13|ICD9CM|Open dislocation of midcarpal (joint)|Open dislocation of midcarpal (joint)
C0159953|T037|AB|833.14|ICD9CM|Disloc carpometacarp-opn|Disloc carpometacarp-opn
C0159953|T037|PT|833.14|ICD9CM|Open dislocation of carpometacarpal (joint)|Open dislocation of carpometacarpal (joint)
C0272826|T037|AB|833.15|ICD9CM|Dislocat metacarpal-open|Dislocat metacarpal-open
C0272826|T037|PT|833.15|ICD9CM|Open dislocation of metacarpal (bone), proximal end|Open dislocation of metacarpal (bone), proximal end
C0159955|T037|AB|833.19|ICD9CM|Dislocat wrist NEC-open|Dislocat wrist NEC-open
C0159955|T037|PT|833.19|ICD9CM|Open dislocation of wrist, other|Open dislocation of wrist, other
C0159956|T037|HT|834|ICD9CM|Dislocation of finger|Dislocation of finger
C0159957|T037|HT|834.0|ICD9CM|Closed dislocation of finger|Closed dislocation of finger
C0375630|T037|PT|834.00|ICD9CM|Closed dislocation of finger, unspecified part|Closed dislocation of finger, unspecified part
C0375630|T037|AB|834.00|ICD9CM|Disl finger NOS-closed|Disl finger NOS-closed
C0272828|T037|PT|834.01|ICD9CM|Closed dislocation of metacarpophalangeal (joint)|Closed dislocation of metacarpophalangeal (joint)
C0272828|T037|AB|834.01|ICD9CM|Disloc metacarpophaln-cl|Disloc metacarpophaln-cl
C1264275|T037|PT|834.02|ICD9CM|Closed dislocation of interphalangeal (joint), hand|Closed dislocation of interphalangeal (joint), hand
C1264275|T037|AB|834.02|ICD9CM|Disl interphaln hand-cl|Disl interphaln hand-cl
C0159960|T037|HT|834.1|ICD9CM|Open dislocation of finger|Open dislocation of finger
C0375631|T037|AB|834.10|ICD9CM|Disloc finger NOS-open|Disloc finger NOS-open
C0375631|T037|PT|834.10|ICD9CM|Open dislocation of finger, unspecified part|Open dislocation of finger, unspecified part
C0159961|T037|AB|834.11|ICD9CM|Disl metacarpophalan-opn|Disl metacarpophalan-opn
C0159961|T037|PT|834.11|ICD9CM|Open dislocation of metacarpophalangeal (joint)|Open dislocation of metacarpophalangeal (joint)
C0159962|T037|AB|834.12|ICD9CM|Disl interphaln hand-opn|Disl interphaln hand-opn
C0159962|T037|PT|834.12|ICD9CM|Open dislocation interphalangeal (joint), hand|Open dislocation interphalangeal (joint), hand
C0019554|T037|HT|835|ICD9CM|Dislocation of hip|Dislocation of hip
C0009041|T037|HT|835.0|ICD9CM|Closed dislocation of hip|Closed dislocation of hip
C0375632|T037|PT|835.00|ICD9CM|Closed dislocation of hip, unspecified site|Closed dislocation of hip, unspecified site
C0375632|T037|AB|835.00|ICD9CM|Dislocat hip NOS-closed|Dislocat hip NOS-closed
C0159963|T037|PT|835.01|ICD9CM|Closed posterior dislocation of hip|Closed posterior dislocation of hip
C0159963|T037|AB|835.01|ICD9CM|Posterior disloc hip-cl|Posterior disloc hip-cl
C0159964|T037|PT|835.02|ICD9CM|Closed obturator dislocation of hip|Closed obturator dislocation of hip
C0159964|T037|AB|835.02|ICD9CM|Obturator disloc hip-cl|Obturator disloc hip-cl
C0159965|T037|AB|835.03|ICD9CM|Ant disloc hip NEC-clos|Ant disloc hip NEC-clos
C0159965|T037|PT|835.03|ICD9CM|Other closed anterior dislocation of hip|Other closed anterior dislocation of hip
C0434666|T037|HT|835.1|ICD9CM|Open dislocation of hip|Open dislocation of hip
C0375633|T037|AB|835.10|ICD9CM|Dislocation hip NOS-open|Dislocation hip NOS-open
C0375633|T037|PT|835.10|ICD9CM|Open dislocation of hip, unspecified site|Open dislocation of hip, unspecified site
C0434663|T037|PT|835.11|ICD9CM|Open posterior dislocation of hip|Open posterior dislocation of hip
C0434663|T037|AB|835.11|ICD9CM|Posterior disloc hip-opn|Posterior disloc hip-opn
C0159968|T037|AB|835.12|ICD9CM|Obturator disloc hip-opn|Obturator disloc hip-opn
C0159968|T037|PT|835.12|ICD9CM|Open obturator dislocation of hip|Open obturator dislocation of hip
C0159969|T037|AB|835.13|ICD9CM|Ant disloc hip NEC-open|Ant disloc hip NEC-open
C0159969|T037|PT|835.13|ICD9CM|Other open anterior dislocation of hip|Other open anterior dislocation of hip
C0159970|T037|HT|836|ICD9CM|Dislocation of knee|Dislocation of knee
C1281729|T037|AB|836.0|ICD9CM|Tear med menisc knee-cur|Tear med menisc knee-cur
C1281729|T037|PT|836.0|ICD9CM|Tear of medial cartilage or meniscus of knee, current|Tear of medial cartilage or meniscus of knee, current
C1281794|T037|AB|836.1|ICD9CM|Tear lat menisc knee-cur|Tear lat menisc knee-cur
C1281794|T037|PT|836.1|ICD9CM|Tear of lateral cartilage or meniscus of knee, current|Tear of lateral cartilage or meniscus of knee, current
C0159973|T037|PT|836.2|ICD9CM|Other tear of cartilage or meniscus of knee, current|Other tear of cartilage or meniscus of knee, current
C0159973|T037|AB|836.2|ICD9CM|Tear meniscus NEC-curren|Tear meniscus NEC-curren
C0434685|T037|AB|836.3|ICD9CM|Dislocat patella-closed|Dislocat patella-closed
C0434685|T037|PT|836.3|ICD9CM|Dislocation of patella, closed|Dislocation of patella, closed
C0159975|T037|PT|836.4|ICD9CM|Dislocation of patella, open|Dislocation of patella, open
C0159975|T037|AB|836.4|ICD9CM|Dislocation patella-open|Dislocation patella-open
C0159976|T037|HT|836.5|ICD9CM|Other dislocation of knee, closed|Other dislocation of knee, closed
C0375634|T037|AB|836.50|ICD9CM|Dislocat knee NOS-closed|Dislocat knee NOS-closed
C0375634|T037|PT|836.50|ICD9CM|Dislocation of knee, unspecified, closed|Dislocation of knee, unspecified, closed
C0159978|T037|AB|836.51|ICD9CM|Ant disloc prox tibia-cl|Ant disloc prox tibia-cl
C0159978|T037|PT|836.51|ICD9CM|Anterior dislocation of tibia, proximal end, closed|Anterior dislocation of tibia, proximal end, closed
C0159979|T037|AB|836.52|ICD9CM|Post disl prox tibia-cl|Post disl prox tibia-cl
C0159979|T037|PT|836.52|ICD9CM|Posterior dislocation of tibia, proximal end, closed|Posterior dislocation of tibia, proximal end, closed
C0159980|T037|AB|836.53|ICD9CM|Med disloc prox tibia-cl|Med disloc prox tibia-cl
C0159980|T037|PT|836.53|ICD9CM|Medial dislocation of tibia, proximal end, closed|Medial dislocation of tibia, proximal end, closed
C0159981|T037|AB|836.54|ICD9CM|Lat disloc prox tibia-cl|Lat disloc prox tibia-cl
C0159981|T037|PT|836.54|ICD9CM|Lateral dislocation of tibia, proximal end, closed|Lateral dislocation of tibia, proximal end, closed
C0159976|T037|AB|836.59|ICD9CM|Dislocat knee NEC-closed|Dislocat knee NEC-closed
C0159976|T037|PT|836.59|ICD9CM|Other dislocation of knee, closed|Other dislocation of knee, closed
C0159982|T037|HT|836.6|ICD9CM|Other dislocation of knee, open|Other dislocation of knee, open
C0272842|T037|AB|836.60|ICD9CM|Dislocat knee NOS-open|Dislocat knee NOS-open
C0272842|T037|PT|836.60|ICD9CM|Dislocation of knee, unspecified, open|Dislocation of knee, unspecified, open
C0159984|T037|AB|836.61|ICD9CM|Ant disl prox tibia-open|Ant disl prox tibia-open
C0159984|T037|PT|836.61|ICD9CM|Anterior dislocation of tibia, proximal end, open|Anterior dislocation of tibia, proximal end, open
C0159985|T037|AB|836.62|ICD9CM|Post disl prox tibia-opn|Post disl prox tibia-opn
C0159985|T037|PT|836.62|ICD9CM|Posterior dislocation of tibia, proximal end, open|Posterior dislocation of tibia, proximal end, open
C0159986|T037|AB|836.63|ICD9CM|Med disl prox tibia-open|Med disl prox tibia-open
C0159986|T037|PT|836.63|ICD9CM|Medial dislocation of tibia, proximal end, open|Medial dislocation of tibia, proximal end, open
C0159987|T037|AB|836.64|ICD9CM|Lat disl prox tibia-open|Lat disl prox tibia-open
C0159987|T037|PT|836.64|ICD9CM|Lateral dislocation of tibia, proximal end, open|Lateral dislocation of tibia, proximal end, open
C0159982|T037|AB|836.69|ICD9CM|Dislocat knee NEC-open|Dislocat knee NEC-open
C0159982|T037|PT|836.69|ICD9CM|Other dislocation of knee, open|Other dislocation of knee, open
C0434691|T037|HT|837|ICD9CM|Dislocation of ankle|Dislocation of ankle
C0434692|T037|PT|837.0|ICD9CM|Closed dislocation of ankle|Closed dislocation of ankle
C0434692|T037|AB|837.0|ICD9CM|Dislocation ankle-closed|Dislocation ankle-closed
C0159990|T037|AB|837.1|ICD9CM|Dislocation ankle-open|Dislocation ankle-open
C0159990|T037|PT|837.1|ICD9CM|Open dislocation of ankle|Open dislocation of ankle
C0434694|T037|HT|838|ICD9CM|Dislocation of foot|Dislocation of foot
C0434696|T037|HT|838.0|ICD9CM|Closed dislocation of foot|Closed dislocation of foot
C0375635|T037|PT|838.00|ICD9CM|Closed dislocation of foot, unspecified|Closed dislocation of foot, unspecified
C0375635|T037|AB|838.00|ICD9CM|Dislocat foot NOS-closed|Dislocat foot NOS-closed
C0159993|T037|PT|838.01|ICD9CM|Closed dislocation of tarsal (bone), joint unspecified|Closed dislocation of tarsal (bone), joint unspecified
C0159993|T037|AB|838.01|ICD9CM|Disloc tarsal NOS-closed|Disloc tarsal NOS-closed
C0159994|T037|PT|838.02|ICD9CM|Closed dislocation of midtarsal (joint)|Closed dislocation of midtarsal (joint)
C0159994|T037|AB|838.02|ICD9CM|Disloc midtarsal-closed|Disloc midtarsal-closed
C0159995|T037|PT|838.03|ICD9CM|Closed dislocation of tarsometatarsal (joint)|Closed dislocation of tarsometatarsal (joint)
C0159995|T037|AB|838.03|ICD9CM|Disloc tarsometatars-cl|Disloc tarsometatars-cl
C0159996|T037|PT|838.04|ICD9CM|Closed dislocation of metatarsal (bone), joint unspecified|Closed dislocation of metatarsal (bone), joint unspecified
C0159996|T037|AB|838.04|ICD9CM|Disloc metatarsal NOS-cl|Disloc metatarsal NOS-cl
C0159997|T037|PT|838.05|ICD9CM|Closed dislocation of metatarsophalangeal (joint)|Closed dislocation of metatarsophalangeal (joint)
C0159997|T037|AB|838.05|ICD9CM|Disl metatarsophalang-cl|Disl metatarsophalang-cl
C0159998|T037|PT|838.06|ICD9CM|Closed dislocation of interphalangeal (joint), foot|Closed dislocation of interphalangeal (joint), foot
C0159998|T037|AB|838.06|ICD9CM|Disl interphalan foot-cl|Disl interphalan foot-cl
C0159999|T037|PT|838.09|ICD9CM|Closed dislocation of foot, other|Closed dislocation of foot, other
C0159999|T037|AB|838.09|ICD9CM|Dislocat foot NEC-closed|Dislocat foot NEC-closed
C0434707|T037|HT|838.1|ICD9CM|Open dislocation of foot|Open dislocation of foot
C0375636|T037|AB|838.10|ICD9CM|Dislocat foot NOS-open|Dislocat foot NOS-open
C0375636|T037|PT|838.10|ICD9CM|Open dislocation of foot, unspecified|Open dislocation of foot, unspecified
C0160001|T037|AB|838.11|ICD9CM|Disloc tarsal NOS-open|Disloc tarsal NOS-open
C0160001|T037|PT|838.11|ICD9CM|Open dislocation of tarsal (bone), joint unspecified|Open dislocation of tarsal (bone), joint unspecified
C0434715|T037|AB|838.12|ICD9CM|Disloc midtarsal-open|Disloc midtarsal-open
C0434715|T037|PT|838.12|ICD9CM|Open dislocation of midtarsal (joint)|Open dislocation of midtarsal (joint)
C0434714|T037|AB|838.13|ICD9CM|Disl tarsometatarsal-opn|Disl tarsometatarsal-opn
C0434714|T037|PT|838.13|ICD9CM|Open dislocation of tarsometatarsal (joint)|Open dislocation of tarsometatarsal (joint)
C0160004|T037|AB|838.14|ICD9CM|Disl metatarsal NOS-open|Disl metatarsal NOS-open
C0160004|T037|PT|838.14|ICD9CM|Open dislocation of metatarsal (bone), joint unspecified|Open dislocation of metatarsal (bone), joint unspecified
C0160005|T037|AB|838.15|ICD9CM|Disloc metatarsophal-opn|Disloc metatarsophal-opn
C0160005|T037|PT|838.15|ICD9CM|Open dislocation of metatarsophalangeal (joint)|Open dislocation of metatarsophalangeal (joint)
C0160006|T037|AB|838.16|ICD9CM|Dis interphalan foot-opn|Dis interphalan foot-opn
C0160006|T037|PT|838.16|ICD9CM|Open dislocation of interphalangeal (joint), foot|Open dislocation of interphalangeal (joint), foot
C0160007|T037|AB|838.19|ICD9CM|Dislocat foot NEC-open|Dislocat foot NEC-open
C0160007|T037|PT|838.19|ICD9CM|Open dislocation of foot, other|Open dislocation of foot, other
C0029876|T037|HT|839|ICD9CM|Other, multiple, and ill-defined dislocations|Other, multiple, and ill-defined dislocations
C0160008|T037|HT|839.0|ICD9CM|Closed dislocation, cervical vertebra|Closed dislocation, cervical vertebra
C0160008|T037|PT|839.00|ICD9CM|Closed dislocation, cervical vertebra, unspecified|Closed dislocation, cervical vertebra, unspecified
C0160008|T037|AB|839.00|ICD9CM|Disloc cerv vert NOS-cl|Disloc cerv vert NOS-cl
C0160009|T037|PT|839.01|ICD9CM|Closed dislocation, first cervical vertebra|Closed dislocation, first cervical vertebra
C0160009|T037|AB|839.01|ICD9CM|Disloc 1st cerv vert-cl|Disloc 1st cerv vert-cl
C0160010|T037|PT|839.02|ICD9CM|Closed dislocation, second cervical vertebra|Closed dislocation, second cervical vertebra
C0160010|T037|AB|839.02|ICD9CM|Disloc 2nd cerv vert-cl|Disloc 2nd cerv vert-cl
C0160011|T037|PT|839.03|ICD9CM|Closed dislocation, third cervical vertebra|Closed dislocation, third cervical vertebra
C0160011|T037|AB|839.03|ICD9CM|Disloc 3rd cerv vert-cl|Disloc 3rd cerv vert-cl
C0160012|T037|PT|839.04|ICD9CM|Closed dislocation, fourth cervical vertebra|Closed dislocation, fourth cervical vertebra
C0160012|T037|AB|839.04|ICD9CM|Disloc 4th cerv vert-cl|Disloc 4th cerv vert-cl
C0160013|T037|PT|839.05|ICD9CM|Closed dislocation, fifth cervical vertebra|Closed dislocation, fifth cervical vertebra
C0160013|T037|AB|839.05|ICD9CM|Disloc 5th cerv vert-cl|Disloc 5th cerv vert-cl
C0160014|T037|PT|839.06|ICD9CM|Closed dislocation, sixth cervical vertebra|Closed dislocation, sixth cervical vertebra
C0160014|T037|AB|839.06|ICD9CM|Disloc 6th cerv vert-cl|Disloc 6th cerv vert-cl
C0160015|T037|PT|839.07|ICD9CM|Closed dislocation, seventh cervical vertebra|Closed dislocation, seventh cervical vertebra
C0160015|T037|AB|839.07|ICD9CM|Disloc 7th cerv vert-cl|Disloc 7th cerv vert-cl
C0160016|T037|PT|839.08|ICD9CM|Closed dislocation, multiple cervical vertebrae|Closed dislocation, multiple cervical vertebrae
C0160016|T037|AB|839.08|ICD9CM|Disloc mult cerv vert-cl|Disloc mult cerv vert-cl
C0160017|T037|HT|839.1|ICD9CM|Open dislocation, cervical vertebra|Open dislocation, cervical vertebra
C0160017|T037|AB|839.10|ICD9CM|Disloc cerv vert NOS-opn|Disloc cerv vert NOS-opn
C0160017|T037|PT|839.10|ICD9CM|Open dislocation, cervical vertebra, unspecified|Open dislocation, cervical vertebra, unspecified
C0160018|T037|AB|839.11|ICD9CM|Disloc lst cerv vert-opn|Disloc lst cerv vert-opn
C0160018|T037|PT|839.11|ICD9CM|Open dislocation, first cervical vertebra|Open dislocation, first cervical vertebra
C0160019|T037|AB|839.12|ICD9CM|Disloc 2nd cerv vert-opn|Disloc 2nd cerv vert-opn
C0160019|T037|PT|839.12|ICD9CM|Open dislocation, second cervical vertebra|Open dislocation, second cervical vertebra
C0160020|T037|AB|839.13|ICD9CM|Disloc 3rd cerv vert-opn|Disloc 3rd cerv vert-opn
C0160020|T037|PT|839.13|ICD9CM|Open dislocation, third cervical vertebra|Open dislocation, third cervical vertebra
C0160021|T037|AB|839.14|ICD9CM|Disloc 4th cerv vert-opn|Disloc 4th cerv vert-opn
C0160021|T037|PT|839.14|ICD9CM|Open dislocation, fourth cervical vertebra|Open dislocation, fourth cervical vertebra
C0160022|T037|AB|839.15|ICD9CM|Disloc 5th cerv vert-opn|Disloc 5th cerv vert-opn
C0160022|T037|PT|839.15|ICD9CM|Open dislocation, fifth cervical vertebra|Open dislocation, fifth cervical vertebra
C0160023|T037|AB|839.16|ICD9CM|Disloc 6th cerv vert-opn|Disloc 6th cerv vert-opn
C0160023|T037|PT|839.16|ICD9CM|Open dislocation, sixth cervical vertebra|Open dislocation, sixth cervical vertebra
C0160024|T037|AB|839.17|ICD9CM|Disloc 7th cerv vert-opn|Disloc 7th cerv vert-opn
C0160024|T037|PT|839.17|ICD9CM|Open dislocation, seventh cervical vertebra|Open dislocation, seventh cervical vertebra
C0160025|T037|AB|839.18|ICD9CM|Disloc mlt cerv vert-opn|Disloc mlt cerv vert-opn
C0160025|T037|PT|839.18|ICD9CM|Open dislocation, multiple cervical vertebrae|Open dislocation, multiple cervical vertebrae
C0160026|T037|HT|839.2|ICD9CM|Closed dislocation, thoracic and lumbar vertebra|Closed dislocation, thoracic and lumbar vertebra
C0160027|T037|PT|839.20|ICD9CM|Closed dislocation, lumbar vertebra|Closed dislocation, lumbar vertebra
C0160027|T037|AB|839.20|ICD9CM|Dislocat lumbar vert-cl|Dislocat lumbar vert-cl
C0160028|T037|PT|839.21|ICD9CM|Closed dislocation, thoracic vertebra|Closed dislocation, thoracic vertebra
C0160028|T037|AB|839.21|ICD9CM|Disloc thoracic vert-cl|Disloc thoracic vert-cl
C0160029|T037|HT|839.3|ICD9CM|Open dislocation, thoracic and lumbar vertebra|Open dislocation, thoracic and lumbar vertebra
C0160030|T037|AB|839.30|ICD9CM|Dislocat lumbar vert-opn|Dislocat lumbar vert-opn
C0160030|T037|PT|839.30|ICD9CM|Open dislocation, lumbar vertebra|Open dislocation, lumbar vertebra
C0160031|T037|AB|839.31|ICD9CM|Disloc thoracic vert-opn|Disloc thoracic vert-opn
C0160031|T037|PT|839.31|ICD9CM|Open dislocation, thoracic vertebra|Open dislocation, thoracic vertebra
C0160032|T037|HT|839.4|ICD9CM|Closed dislocation, other vertebra|Closed dislocation, other vertebra
C0160033|T037|PT|839.40|ICD9CM|Closed dislocation, vertebra, unspecified site|Closed dislocation, vertebra, unspecified site
C0160033|T037|AB|839.40|ICD9CM|Dislocat vertebra NOS-cl|Dislocat vertebra NOS-cl
C0160034|T037|PT|839.41|ICD9CM|Closed dislocation, coccyx|Closed dislocation, coccyx
C0160034|T037|AB|839.41|ICD9CM|Dislocat coccyx-closed|Dislocat coccyx-closed
C0160035|T037|PT|839.42|ICD9CM|Closed dislocation, sacrum|Closed dislocation, sacrum
C0160035|T037|AB|839.42|ICD9CM|Dislocat sacrum-closed|Dislocat sacrum-closed
C0160032|T037|PT|839.49|ICD9CM|Closed dislocation, vertebra, other|Closed dislocation, vertebra, other
C0160032|T037|AB|839.49|ICD9CM|Dislocat vertebra NEC-cl|Dislocat vertebra NEC-cl
C0160036|T037|HT|839.5|ICD9CM|Open dislocation, other vertebra|Open dislocation, other vertebra
C0160037|T037|AB|839.50|ICD9CM|Disloc vertebra NOS-open|Disloc vertebra NOS-open
C0160037|T037|PT|839.50|ICD9CM|Open dislocation, vertebra, unspecified site|Open dislocation, vertebra, unspecified site
C0160038|T037|AB|839.51|ICD9CM|Dislocat coccyx-open|Dislocat coccyx-open
C0160038|T037|PT|839.51|ICD9CM|Open dislocation, coccyx|Open dislocation, coccyx
C0160039|T037|AB|839.52|ICD9CM|Dislocat sacrum-open|Dislocat sacrum-open
C0160039|T037|PT|839.52|ICD9CM|Open dislocation, sacrum|Open dislocation, sacrum
C0160036|T037|AB|839.59|ICD9CM|Disloc vertebra NEC-open|Disloc vertebra NEC-open
C0160036|T037|PT|839.59|ICD9CM|Open dislocation, vertebra,other|Open dislocation, vertebra,other
C0160040|T037|HT|839.6|ICD9CM|Closed dislocation, other location|Closed dislocation, other location
C0160041|T037|PT|839.61|ICD9CM|Closed dislocation, sternum|Closed dislocation, sternum
C0160041|T037|AB|839.61|ICD9CM|Dislocat sternum-closed|Dislocat sternum-closed
C0160040|T037|PT|839.69|ICD9CM|Closed dislocation, other location|Closed dislocation, other location
C0160040|T037|AB|839.69|ICD9CM|Dislocat site NEC-closed|Dislocat site NEC-closed
C0160042|T037|HT|839.7|ICD9CM|Open dislocation, other location|Open dislocation, other location
C0160043|T037|AB|839.71|ICD9CM|Dislocation sternum-open|Dislocation sternum-open
C0160043|T037|PT|839.71|ICD9CM|Open dislocation, sternum|Open dislocation, sternum
C0160042|T037|AB|839.79|ICD9CM|Dislocat site NEC-open|Dislocat site NEC-open
C0160042|T037|PT|839.79|ICD9CM|Open dislocation, other location|Open dislocation, other location
C0009043|T037|PT|839.8|ICD9CM|Closed dislocation, multiple and ill-defined sites|Closed dislocation, multiple and ill-defined sites
C0009043|T037|AB|839.8|ICD9CM|Dislocation NEC-closed|Dislocation NEC-closed
C0160044|T037|AB|839.9|ICD9CM|Dislocation NEC-open|Dislocation NEC-open
C0160044|T037|PT|839.9|ICD9CM|Open dislocation, multiple and ill-defined sites|Open dislocation, multiple and ill-defined sites
C0160045|T037|HT|840|ICD9CM|Sprains and strains of shoulder and upper arm|Sprains and strains of shoulder and upper arm
C0038048|T037|HT|840-848.99|ICD9CM|SPRAINS AND STRAINS OF JOINTS AND ADJACENT MUSCLES|SPRAINS AND STRAINS OF JOINTS AND ADJACENT MUSCLES
C0272870|T037|PT|840.0|ICD9CM|Acromioclavicular (joint) (ligament) sprain|Acromioclavicular (joint) (ligament) sprain
C0272870|T037|AB|840.0|ICD9CM|Sprain acromioclavicular|Sprain acromioclavicular
C0160047|T037|PT|840.1|ICD9CM|Coracoclavicular (ligament) sprain|Coracoclavicular (ligament) sprain
C0160047|T037|AB|840.1|ICD9CM|Sprain coracoclavicular|Sprain coracoclavicular
C0435003|T037|PT|840.2|ICD9CM|Coracohumeral (ligament) sprain|Coracohumeral (ligament) sprain
C0435003|T037|AB|840.2|ICD9CM|Sprain coracohumeral|Sprain coracohumeral
C1306110|T037|PT|840.3|ICD9CM|Infraspinatus (muscle) (tendon) sprain|Infraspinatus (muscle) (tendon) sprain
C1306110|T037|AB|840.3|ICD9CM|Sprain infraspinatus|Sprain infraspinatus
C0434322|T037|PT|840.4|ICD9CM|Rotator cuff (capsule) sprain|Rotator cuff (capsule) sprain
C0434322|T037|AB|840.4|ICD9CM|Sprain rotator cuff|Sprain rotator cuff
C0160051|T037|AB|840.5|ICD9CM|Sprain subscapularis|Sprain subscapularis
C0160051|T037|PT|840.5|ICD9CM|Subscapularis (muscle) sprain|Subscapularis (muscle) sprain
C0749173|T037|AB|840.6|ICD9CM|Sprain supraspinatus|Sprain supraspinatus
C0749173|T037|PT|840.6|ICD9CM|Supraspinatus (muscle) (tendon) sprain|Supraspinatus (muscle) (tendon) sprain
C0949149|T037|AB|840.7|ICD9CM|Sup glenoid labrm lesion|Sup glenoid labrm lesion
C0949149|T037|PT|840.7|ICD9CM|Superior glenoid labrum lesion|Superior glenoid labrum lesion
C0160053|T037|AB|840.8|ICD9CM|Sprain shoulder/arm NEC|Sprain shoulder/arm NEC
C0160053|T037|PT|840.8|ICD9CM|Sprains and strains of other specified sites of shoulder and upper arm|Sprains and strains of other specified sites of shoulder and upper arm
C0160054|T037|AB|840.9|ICD9CM|Sprain shoulder/arm NOS|Sprain shoulder/arm NOS
C0160054|T037|PT|840.9|ICD9CM|Sprains and strains of unspecified site of shoulder and upper arm|Sprains and strains of unspecified site of shoulder and upper arm
C0160055|T037|HT|841|ICD9CM|Sprains and strains of elbow and forearm|Sprains and strains of elbow and forearm
C0160056|T037|PT|841.0|ICD9CM|Radial collateral ligament sprain|Radial collateral ligament sprain
C0160056|T037|AB|841.0|ICD9CM|Sprain radial collat lig|Sprain radial collat lig
C0160057|T037|AB|841.1|ICD9CM|Sprain ulnar collat lig|Sprain ulnar collat lig
C0160057|T037|PT|841.1|ICD9CM|Ulnar collateral ligament sprain|Ulnar collateral ligament sprain
C0160058|T037|PT|841.2|ICD9CM|Radiohumeral (joint) sprain|Radiohumeral (joint) sprain
C0160058|T037|AB|841.2|ICD9CM|Sprain radiohumeral|Sprain radiohumeral
C0160059|T037|AB|841.3|ICD9CM|Sprain ulnohumeral|Sprain ulnohumeral
C0160059|T037|PT|841.3|ICD9CM|Ulnohumeral (joint) sprain|Ulnohumeral (joint) sprain
C0160060|T037|AB|841.8|ICD9CM|Sprain elbow/forearm NEC|Sprain elbow/forearm NEC
C0160060|T037|PT|841.8|ICD9CM|Sprains and strains of other specified sites of elbow and forearm|Sprains and strains of other specified sites of elbow and forearm
C0160061|T037|AB|841.9|ICD9CM|Sprain elbow/forearm NOS|Sprain elbow/forearm NOS
C0160061|T037|PT|841.9|ICD9CM|Sprains and strains of unspecified site of elbow and forearm|Sprains and strains of unspecified site of elbow and forearm
C0160062|T037|HT|842|ICD9CM|Sprains and strains of wrist and hand|Sprains and strains of wrist and hand
C0160063|T037|HT|842.0|ICD9CM|Wrist sprain|Wrist sprain
C0160063|T037|AB|842.00|ICD9CM|Sprain of wrist NOS|Sprain of wrist NOS
C0160063|T037|PT|842.00|ICD9CM|Sprain of wrist, unspecified site|Sprain of wrist, unspecified site
C0272880|T037|AB|842.01|ICD9CM|Sprain carpal|Sprain carpal
C0272880|T037|PT|842.01|ICD9CM|Sprain of carpal (joint) of wrist|Sprain of carpal (joint) of wrist
C0272881|T037|PT|842.02|ICD9CM|Sprain of radiocarpal (joint) (ligament) of wrist|Sprain of radiocarpal (joint) (ligament) of wrist
C0272881|T037|AB|842.02|ICD9CM|Sprain radiocarpal|Sprain radiocarpal
C0160067|T037|PT|842.09|ICD9CM|Other sprains and strains of wrist|Other sprains and strains of wrist
C0160067|T037|AB|842.09|ICD9CM|Sprain of wrist NEC|Sprain of wrist NEC
C0160068|T037|HT|842.1|ICD9CM|Hand sprain|Hand sprain
C0160068|T037|AB|842.10|ICD9CM|Sprain of hand NOS|Sprain of hand NOS
C0160068|T037|PT|842.10|ICD9CM|Sprain of hand, unspecified site|Sprain of hand, unspecified site
C0160070|T037|AB|842.11|ICD9CM|Sprain carpometacarpal|Sprain carpometacarpal
C0160070|T037|PT|842.11|ICD9CM|Sprain of carpometacarpal (joint) of hand|Sprain of carpometacarpal (joint) of hand
C0160071|T037|AB|842.12|ICD9CM|Sprain metacarpophalang|Sprain metacarpophalang
C0160071|T037|PT|842.12|ICD9CM|Sprain of metacarpophalangeal (joint) of hand|Sprain of metacarpophalangeal (joint) of hand
C0160072|T037|AB|842.13|ICD9CM|Sprain interphalangeal|Sprain interphalangeal
C0160072|T037|PT|842.13|ICD9CM|Sprain of interphalangeal (joint) of hand|Sprain of interphalangeal (joint) of hand
C0160073|T037|PT|842.19|ICD9CM|Other sprains and strains of hand|Other sprains and strains of hand
C0160073|T037|AB|842.19|ICD9CM|Sprain of hand NEC|Sprain of hand NEC
C0160074|T037|HT|843|ICD9CM|Sprains and strains of hip and thigh|Sprains and strains of hip and thigh
C0160075|T037|PT|843.0|ICD9CM|Iliofemoral (ligament) sprain|Iliofemoral (ligament) sprain
C0160075|T037|AB|843.0|ICD9CM|Sprain iliofemoral|Sprain iliofemoral
C0434483|T037|PT|843.1|ICD9CM|Ischiocapsular (ligament) sprain|Ischiocapsular (ligament) sprain
C0434483|T037|AB|843.1|ICD9CM|Sprain ischiocapsular|Sprain ischiocapsular
C0160077|T037|AB|843.8|ICD9CM|Sprain hip & thigh NEC|Sprain hip & thigh NEC
C0160077|T037|PT|843.8|ICD9CM|Sprains and strains of other specified sites of hip and thigh|Sprains and strains of other specified sites of hip and thigh
C0160078|T037|AB|843.9|ICD9CM|Sprain hip & thigh NOS|Sprain hip & thigh NOS
C0160078|T037|PT|843.9|ICD9CM|Sprains and strains of unspecified site of hip and thigh|Sprains and strains of unspecified site of hip and thigh
C0160079|T037|HT|844|ICD9CM|Sprains and strains of knee and leg|Sprains and strains of knee and leg
C0160080|T037|AB|844.0|ICD9CM|Sprain lateral coll lig|Sprain lateral coll lig
C0160080|T037|PT|844.0|ICD9CM|Sprain of lateral collateral ligament of knee|Sprain of lateral collateral ligament of knee
C0160081|T037|AB|844.1|ICD9CM|Sprain medial collat lig|Sprain medial collat lig
C0160081|T037|PT|844.1|ICD9CM|Sprain of medial collateral ligament of knee|Sprain of medial collateral ligament of knee
C0160082|T037|AB|844.2|ICD9CM|Sprain cruciate lig knee|Sprain cruciate lig knee
C0160082|T037|PT|844.2|ICD9CM|Sprain of cruciate ligament of knee|Sprain of cruciate ligament of knee
C0435018|T037|PT|844.3|ICD9CM|Sprain of tibiofibular (joint) (ligament) superior, of knee|Sprain of tibiofibular (joint) (ligament) superior, of knee
C0435018|T037|AB|844.3|ICD9CM|Sprain super tibiofibula|Sprain super tibiofibula
C0160084|T037|AB|844.8|ICD9CM|Sprain of knee & leg NEC|Sprain of knee & leg NEC
C0160084|T037|PT|844.8|ICD9CM|Sprains and strains of other specified sites of knee and leg|Sprains and strains of other specified sites of knee and leg
C0160085|T037|AB|844.9|ICD9CM|Sprain of knee & leg NOS|Sprain of knee & leg NOS
C0160085|T037|PT|844.9|ICD9CM|Sprains and strains of unspecified site of knee and leg|Sprains and strains of unspecified site of knee and leg
C0160086|T037|HT|845|ICD9CM|Sprains and strains of ankle and foot|Sprains and strains of ankle and foot
C0160087|T037|HT|845.0|ICD9CM|Ankle sprain|Ankle sprain
C0160087|T037|AB|845.00|ICD9CM|Sprain of ankle NOS|Sprain of ankle NOS
C0160087|T037|PT|845.00|ICD9CM|Sprain of ankle, unspecified site|Sprain of ankle, unspecified site
C0160089|T037|AB|845.01|ICD9CM|Sprain of ankle deltoid|Sprain of ankle deltoid
C0160089|T037|PT|845.01|ICD9CM|Sprain of deltoid (ligament), ankle|Sprain of deltoid (ligament), ankle
C0160090|T037|AB|845.02|ICD9CM|Sprain calcaneofibular|Sprain calcaneofibular
C0160090|T037|PT|845.02|ICD9CM|Sprain of calcaneofibular (ligament) of ankle|Sprain of calcaneofibular (ligament) of ankle
C0160091|T037|AB|845.03|ICD9CM|Sprain distal tibiofibul|Sprain distal tibiofibul
C0160091|T037|PT|845.03|ICD9CM|Sprain of tibiofibular (ligament), distal of ankle|Sprain of tibiofibular (ligament), distal of ankle
C0160092|T037|PT|845.09|ICD9CM|Other sprains and strains of ankle|Other sprains and strains of ankle
C0160092|T037|AB|845.09|ICD9CM|Sprain of ankle NEC|Sprain of ankle NEC
C0160093|T037|HT|845.1|ICD9CM|Foot sprain|Foot sprain
C0160094|T037|AB|845.10|ICD9CM|Sprain of foot NOS|Sprain of foot NOS
C0160094|T037|PT|845.10|ICD9CM|Sprain of foot, unspecified site|Sprain of foot, unspecified site
C0272905|T037|PT|845.11|ICD9CM|Sprain of tarsometatarsal (joint) (ligament) of foot|Sprain of tarsometatarsal (joint) (ligament) of foot
C0272905|T037|AB|845.11|ICD9CM|Sprain tarsometatarsal|Sprain tarsometatarsal
C0160096|T037|AB|845.12|ICD9CM|Sprain metatarsophalang|Sprain metatarsophalang
C0160096|T037|PT|845.12|ICD9CM|Sprain of metatarsophalangeal (joint) of foot|Sprain of metatarsophalangeal (joint) of foot
C0160097|T037|AB|845.13|ICD9CM|Sprain interphalang toe|Sprain interphalang toe
C0160097|T037|PT|845.13|ICD9CM|Sprain of interphalangeal (joint), toe|Sprain of interphalangeal (joint), toe
C0160098|T037|PT|845.19|ICD9CM|Other sprain of foot|Other sprain of foot
C0160098|T037|AB|845.19|ICD9CM|Sprain of foot NEC|Sprain of foot NEC
C0160099|T037|HT|846|ICD9CM|Sprains and strains of sacroiliac region|Sprains and strains of sacroiliac region
C0272914|T037|AB|846.0|ICD9CM|Sprain lumbosacral|Sprain lumbosacral
C0272914|T037|PT|846.0|ICD9CM|Sprain of lumbosacral (joint) (ligament)|Sprain of lumbosacral (joint) (ligament)
C0434473|T037|PT|846.1|ICD9CM|Sprain of sacroiliac ligament|Sprain of sacroiliac ligament
C0434473|T037|AB|846.1|ICD9CM|Sprain sacroiliac|Sprain sacroiliac
C0160102|T037|PT|846.2|ICD9CM|Sprain of sacrospinatus (ligament)|Sprain of sacrospinatus (ligament)
C0160102|T037|AB|846.2|ICD9CM|Sprain sacrospinatus|Sprain sacrospinatus
C0160103|T037|PT|846.3|ICD9CM|Sprain of sacrotuberous (ligament)|Sprain of sacrotuberous (ligament)
C0160103|T037|AB|846.3|ICD9CM|Sprain sacrotuberous|Sprain sacrotuberous
C0160104|T037|PT|846.8|ICD9CM|Sprain of other specified sites of sacroiliac region|Sprain of other specified sites of sacroiliac region
C0160104|T037|AB|846.8|ICD9CM|Sprain sacroiliac NEC|Sprain sacroiliac NEC
C0160105|T037|PT|846.9|ICD9CM|Sprain of unspecified site of sacroiliac region|Sprain of unspecified site of sacroiliac region
C0160105|T037|AB|846.9|ICD9CM|Sprain sacroiliac NOS|Sprain sacroiliac NOS
C0160106|T037|HT|847|ICD9CM|Sprains and strains of other and unspecified parts of back|Sprains and strains of other and unspecified parts of back
C0027535|T037|AB|847.0|ICD9CM|Sprain of neck|Sprain of neck
C0027535|T037|PT|847.0|ICD9CM|Sprain of neck|Sprain of neck
C0160107|T037|PT|847.1|ICD9CM|Sprain of thoracic|Sprain of thoracic
C0160107|T037|AB|847.1|ICD9CM|Sprain thoracic region|Sprain thoracic region
C0160108|T037|AB|847.2|ICD9CM|Sprain lumbar region|Sprain lumbar region
C0160108|T037|PT|847.2|ICD9CM|Sprain of lumbar|Sprain of lumbar
C0160109|T037|AB|847.3|ICD9CM|Sprain of sacrum|Sprain of sacrum
C0160109|T037|PT|847.3|ICD9CM|Sprain of sacrum|Sprain of sacrum
C0160110|T037|AB|847.4|ICD9CM|Sprain of coccyx|Sprain of coccyx
C0160110|T037|PT|847.4|ICD9CM|Sprain of coccyx|Sprain of coccyx
C0160111|T037|AB|847.9|ICD9CM|Sprain of back NOS|Sprain of back NOS
C0160111|T037|PT|847.9|ICD9CM|Sprain of unspecified site of back|Sprain of unspecified site of back
C0029490|T037|HT|848|ICD9CM|Other and ill-defined sprains and strains|Other and ill-defined sprains and strains
C0160112|T037|AB|848.0|ICD9CM|Sprain of nasal septum|Sprain of nasal septum
C0160112|T037|PT|848.0|ICD9CM|Sprain of septal cartilage of nose|Sprain of septal cartilage of nose
C0160113|T037|AB|848.1|ICD9CM|Sprain of jaw|Sprain of jaw
C0160113|T037|PT|848.1|ICD9CM|Sprain of jaw|Sprain of jaw
C0160114|T037|AB|848.2|ICD9CM|Sprain of thyroid region|Sprain of thyroid region
C0160114|T037|PT|848.2|ICD9CM|Sprain of thyroid region|Sprain of thyroid region
C0160115|T037|AB|848.3|ICD9CM|Sprain of ribs|Sprain of ribs
C0160115|T037|PT|848.3|ICD9CM|Sprain of ribs|Sprain of ribs
C0434411|T037|HT|848.4|ICD9CM|Sternum sprain|Sternum sprain
C0434411|T037|AB|848.40|ICD9CM|Sprain of sternum NOS|Sprain of sternum NOS
C0434411|T037|PT|848.40|ICD9CM|Sprain of sternum, unspecified site|Sprain of sternum, unspecified site
C0272920|T037|PT|848.41|ICD9CM|Sprain of sternoclavicular (joint) (ligament)|Sprain of sternoclavicular (joint) (ligament)
C0272920|T037|AB|848.41|ICD9CM|Sprain sternoclavicular|Sprain sternoclavicular
C0160118|T037|AB|848.42|ICD9CM|Sprain chondrosternal|Sprain chondrosternal
C0160118|T037|PT|848.42|ICD9CM|Sprain of chondrosternal (joint)|Sprain of chondrosternal (joint)
C0160119|T037|AB|848.49|ICD9CM|Sprain of sternum NEC|Sprain of sternum NEC
C0160119|T037|PT|848.49|ICD9CM|Sprain of sternum, other|Sprain of sternum, other
C0435019|T037|PT|848.5|ICD9CM|Sprain of pelvic|Sprain of pelvic
C0435019|T037|AB|848.5|ICD9CM|Sprain of pelvis|Sprain of pelvis
C0029829|T037|PT|848.8|ICD9CM|Other specified sites of sprains and strains|Other specified sites of sprains and strains
C0029829|T037|AB|848.8|ICD9CM|Sprain NEC|Sprain NEC
C0041887|T037|AB|848.9|ICD9CM|Sprain NOS|Sprain NOS
C0041887|T037|PT|848.9|ICD9CM|Unspecified site of sprain and strain|Unspecified site of sprain and strain
C0006107|T037|HT|850|ICD9CM|Concussion|Concussion
C0178319|T037|HT|850-854.99|ICD9CM|INTRACRANIAL INJURY, EXCLUDING THOSE WITH SKULL FRACTURE|INTRACRANIAL INJURY, EXCLUDING THOSE WITH SKULL FRACTURE
C0160121|T037|AB|850.0|ICD9CM|Concussion w/o coma|Concussion w/o coma
C0160121|T037|PT|850.0|ICD9CM|Concussion with no loss of consciousness|Concussion with no loss of consciousness
C0160122|T037|HT|850.1|ICD9CM|Concussion with brief loss of consciousness|Concussion with brief loss of consciousness
C1260444|T037|AB|850.11|ICD9CM|Concus-brief coma <31 mn|Concus-brief coma <31 mn
C1260444|T037|PT|850.11|ICD9CM|Concussion, with loss of consciousness of 30 minutes or less|Concussion, with loss of consciousness of 30 minutes or less
C1260445|T037|AB|850.12|ICD9CM|Concus-brf coma 31-59 mn|Concus-brf coma 31-59 mn
C1260445|T037|PT|850.12|ICD9CM|Concussion, with loss of consciousness from 31 to 59 minutes|Concussion, with loss of consciousness from 31 to 59 minutes
C0160123|T037|PT|850.2|ICD9CM|Concussion with moderate loss of consciousness|Concussion with moderate loss of consciousness
C0160123|T037|AB|850.2|ICD9CM|Concussion-moderate coma|Concussion-moderate coma
C0160124|T037|PT|850.3|ICD9CM|Concussion with prolonged loss of consciousness and return to pre-existing conscious level|Concussion with prolonged loss of consciousness and return to pre-existing conscious level
C0160124|T037|AB|850.3|ICD9CM|Concussion-prolong coma|Concussion-prolong coma
C0160125|T037|PT|850.4|ICD9CM|Concussion with prolonged loss of consciousness, without return to pre-existing conscious level|Concussion with prolonged loss of consciousness, without return to pre-existing conscious level
C0160125|T037|AB|850.4|ICD9CM|Concussion-deep coma|Concussion-deep coma
C0160126|T037|AB|850.5|ICD9CM|Concussion w coma NOS|Concussion w coma NOS
C0160126|T037|PT|850.5|ICD9CM|Concussion with loss of consciousness of unspecified duration|Concussion with loss of consciousness of unspecified duration
C0006107|T037|AB|850.9|ICD9CM|Concussion NOS|Concussion NOS
C0006107|T037|PT|850.9|ICD9CM|Concussion, unspecified|Concussion, unspecified
C0160127|T037|HT|851|ICD9CM|Cerebral laceration and contusion|Cerebral laceration and contusion
C0160128|T037|HT|851.0|ICD9CM|Cortex (cerebral) contusion without mention of open intracranial wound|Cortex (cerebral) contusion without mention of open intracranial wound
C0433815|T037|AB|851.00|ICD9CM|Cerebral cortx contusion|Cerebral cortx contusion
C0433816|T037|AB|851.01|ICD9CM|Cortex contusion-no coma|Cortex contusion-no coma
C0160131|T037|AB|851.02|ICD9CM|Cortex contus-brief coma|Cortex contus-brief coma
C0272955|T037|AB|851.03|ICD9CM|Cortex contus-mod coma|Cortex contus-mod coma
C0160133|T037|AB|851.04|ICD9CM|Cortx contus-prolng coma|Cortx contus-prolng coma
C0160134|T037|AB|851.05|ICD9CM|Cortex contus-deep coma|Cortex contus-deep coma
C0433821|T037|AB|851.06|ICD9CM|Cortex contus-coma NOS|Cortex contus-coma NOS
C0695217|T037|PT|851.09|ICD9CM|Cortex (cerebral) contusion without mention of open intracranial wound, with concussion, unspecified|Cortex (cerebral) contusion without mention of open intracranial wound, with concussion, unspecified
C0695217|T037|AB|851.09|ICD9CM|Cortex contus-concus NOS|Cortex contus-concus NOS
C0160137|T037|HT|851.1|ICD9CM|Cortex (cerebral) contusion with open intracranial wound|Cortex (cerebral) contusion with open intracranial wound
C0160138|T037|PT|851.10|ICD9CM|Cortex (cerebral) contusion with open intracranial wound, unspecified state of consciousness|Cortex (cerebral) contusion with open intracranial wound, unspecified state of consciousness
C0160138|T037|AB|851.10|ICD9CM|Cortex contusion/opn wnd|Cortex contusion/opn wnd
C0272961|T037|PT|851.11|ICD9CM|Cortex (cerebral) contusion with open intracranial wound, with no loss of consciousness|Cortex (cerebral) contusion with open intracranial wound, with no loss of consciousness
C0272961|T037|AB|851.11|ICD9CM|Opn cortx contus-no coma|Opn cortx contus-no coma
C0160140|T037|AB|851.12|ICD9CM|Opn cort contus-brf coma|Opn cort contus-brf coma
C0160141|T037|AB|851.13|ICD9CM|Opn cort contus-mod coma|Opn cort contus-mod coma
C0160142|T037|AB|851.14|ICD9CM|Opn cort contu-prol coma|Opn cort contu-prol coma
C0160143|T037|AB|851.15|ICD9CM|Opn cort contu-deep coma|Opn cort contu-deep coma
C0272966|T037|AB|851.16|ICD9CM|Opn cort contus-coma NOS|Opn cort contus-coma NOS
C0272967|T037|PT|851.19|ICD9CM|Cortex (cerebral) contusion with open intracranial wound, with concussion, unspecified|Cortex (cerebral) contusion with open intracranial wound, with concussion, unspecified
C0272967|T037|AB|851.19|ICD9CM|Opn cortx contus-concuss|Opn cortx contus-concuss
C0433846|T037|HT|851.2|ICD9CM|Cortex (cerebral) laceration without mention of open intracranial wound|Cortex (cerebral) laceration without mention of open intracranial wound
C0433847|T037|AB|851.20|ICD9CM|Cerebral cortex lacerat|Cerebral cortex lacerat
C0433848|T037|AB|851.21|ICD9CM|Cortex lacerat w/o coma|Cortex lacerat w/o coma
C0160149|T037|AB|851.22|ICD9CM|Cortex lacera-brief coma|Cortex lacera-brief coma
C0160150|T037|AB|851.23|ICD9CM|Cortex lacerat-mod coma|Cortex lacerat-mod coma
C0160151|T037|AB|851.24|ICD9CM|Cortex lacerat-prol coma|Cortex lacerat-prol coma
C0160152|T037|AB|851.25|ICD9CM|Cortex lacerat-deep coma|Cortex lacerat-deep coma
C0433853|T037|AB|851.26|ICD9CM|Cortex lacerat-coma NOS|Cortex lacerat-coma NOS
C0433854|T037|AB|851.29|ICD9CM|Cortex lacerat-concuss|Cortex lacerat-concuss
C0272977|T037|HT|851.3|ICD9CM|Cortex (cerebral) laceration with open intracranial wound|Cortex (cerebral) laceration with open intracranial wound
C0272978|T037|PT|851.30|ICD9CM|Cortex (cerebral) laceration with open intracranial wound, unspecified state of consciousness|Cortex (cerebral) laceration with open intracranial wound, unspecified state of consciousness
C0272978|T037|AB|851.30|ICD9CM|Cortex lacer w opn wound|Cortex lacer w opn wound
C0272979|T037|PT|851.31|ICD9CM|Cortex (cerebral) laceration with open intracranial wound, with no loss of consciousness|Cortex (cerebral) laceration with open intracranial wound, with no loss of consciousness
C0272979|T037|AB|851.31|ICD9CM|Opn cortex lacer-no coma|Opn cortex lacer-no coma
C0160158|T037|AB|851.32|ICD9CM|Opn cortx lac-brief coma|Opn cortx lac-brief coma
C0160159|T037|AB|851.33|ICD9CM|Opn cortx lacer-mod coma|Opn cortx lacer-mod coma
C0160160|T037|AB|851.34|ICD9CM|Opn cortx lac-proln coma|Opn cortx lac-proln coma
C0433845|T037|AB|851.35|ICD9CM|Opn cortex lac-deep coma|Opn cortex lac-deep coma
C0272984|T037|AB|851.36|ICD9CM|Opn cortx lacer-coma NOS|Opn cortx lacer-coma NOS
C0272985|T037|PT|851.39|ICD9CM|Cortex (cerebral) laceration with open intracranial wound, with concussion, unspecified|Cortex (cerebral) laceration with open intracranial wound, with concussion, unspecified
C0272985|T037|AB|851.39|ICD9CM|Opn cortx lacer-concuss|Opn cortx lacer-concuss
C0160164|T037|HT|851.4|ICD9CM|Cerebellar or brain stem contusion without mention of open intracranial wound|Cerebellar or brain stem contusion without mention of open intracranial wound
C0160165|T037|AB|851.40|ICD9CM|Cerebel/brain stm contus|Cerebel/brain stm contus
C0160166|T037|AB|851.41|ICD9CM|Cerebell contus w/o coma|Cerebell contus w/o coma
C0160167|T037|AB|851.42|ICD9CM|Cerebell contus-brf coma|Cerebell contus-brf coma
C0160168|T037|AB|851.43|ICD9CM|Cerebell contus-mod coma|Cerebell contus-mod coma
C0160169|T037|AB|851.44|ICD9CM|Cerebel contus-prol coma|Cerebel contus-prol coma
C0160170|T037|AB|851.45|ICD9CM|Cerebel contus-deep coma|Cerebel contus-deep coma
C0160171|T037|AB|851.46|ICD9CM|Cerebell contus-coma NOS|Cerebell contus-coma NOS
C0695221|T037|AB|851.49|ICD9CM|Cerebell contus-concuss|Cerebell contus-concuss
C0160173|T037|HT|851.5|ICD9CM|Cerebellar or brain stem contusion with open intracranial wound|Cerebellar or brain stem contusion with open intracranial wound
C0160174|T037|AB|851.50|ICD9CM|Cerebel contus w opn wnd|Cerebel contus w opn wnd
C0160174|T037|PT|851.50|ICD9CM|Cerebellar or brain stem contusion with open intracranial wound, unspecified state of consciousness|Cerebellar or brain stem contusion with open intracranial wound, unspecified state of consciousness
C0160175|T037|PT|851.51|ICD9CM|Cerebellar or brain stem contusion with open intracranial wound, with no loss of consciousness|Cerebellar or brain stem contusion with open intracranial wound, with no loss of consciousness
C0160175|T037|AB|851.51|ICD9CM|Opn cerebe cont w/o coma|Opn cerebe cont w/o coma
C0160176|T037|AB|851.52|ICD9CM|Opn cerebe cont-brf coma|Opn cerebe cont-brf coma
C0160177|T037|AB|851.53|ICD9CM|Opn cerebe cont-mod coma|Opn cerebe cont-mod coma
C0160178|T037|AB|851.54|ICD9CM|Opn cerebe cont-prol com|Opn cerebe cont-prol com
C0160179|T037|AB|851.55|ICD9CM|Opn cerebe cont-deep com|Opn cerebe cont-deep com
C0160180|T037|AB|851.56|ICD9CM|Opn cerebe cont-coma NOS|Opn cerebe cont-coma NOS
C0695222|T037|PT|851.59|ICD9CM|Cerebellar or brain stem contusion with open intracranial wound, with concussion, unspecified|Cerebellar or brain stem contusion with open intracranial wound, with concussion, unspecified
C0695222|T037|AB|851.59|ICD9CM|Opn cerebel cont-concuss|Opn cerebel cont-concuss
C0160182|T037|HT|851.6|ICD9CM|Cerebellar or brain stem laceration without mention of open intracranial wound|Cerebellar or brain stem laceration without mention of open intracranial wound
C0160183|T037|AB|851.60|ICD9CM|Cerebel/brain stem lacer|Cerebel/brain stem lacer
C0160184|T037|AB|851.61|ICD9CM|Cerebel lacerat w/o coma|Cerebel lacerat w/o coma
C0160185|T037|AB|851.62|ICD9CM|Cerebel lacer-brief coma|Cerebel lacer-brief coma
C0160186|T037|AB|851.63|ICD9CM|Cerebel lacerat-mod coma|Cerebel lacerat-mod coma
C0160187|T037|AB|851.64|ICD9CM|Cerebel lacer-proln coma|Cerebel lacer-proln coma
C0160188|T037|AB|851.65|ICD9CM|Cerebell lacer-deep coma|Cerebell lacer-deep coma
C0160189|T037|AB|851.66|ICD9CM|Cerebel lacerat-coma NOS|Cerebel lacerat-coma NOS
C0695223|T037|AB|851.69|ICD9CM|Cerebel lacer-concussion|Cerebel lacer-concussion
C0160191|T037|HT|851.7|ICD9CM|Cerebellar or brain stem laceration with open intracranial wound|Cerebellar or brain stem laceration with open intracranial wound
C0160192|T037|AB|851.70|ICD9CM|Cerebel lacer w open wnd|Cerebel lacer w open wnd
C0160192|T037|PT|851.70|ICD9CM|Cerebellar or brain stem laceration with open intracranial wound, unspecified state of consciousness|Cerebellar or brain stem laceration with open intracranial wound, unspecified state of consciousness
C0160193|T037|PT|851.71|ICD9CM|Cerebellar or brain stem laceration with open intracranial wound, with no loss of consciousness|Cerebellar or brain stem laceration with open intracranial wound, with no loss of consciousness
C0160193|T037|AB|851.71|ICD9CM|Opn cerebel lac w/o coma|Opn cerebel lac w/o coma
C0160194|T037|AB|851.72|ICD9CM|Opn cerebel lac-brf coma|Opn cerebel lac-brf coma
C0160195|T037|AB|851.73|ICD9CM|Opn cerebel lac-mod coma|Opn cerebel lac-mod coma
C0160196|T037|AB|851.74|ICD9CM|Opn cerebe lac-prol coma|Opn cerebe lac-prol coma
C0160197|T037|AB|851.75|ICD9CM|Opn cerebe lac-deep coma|Opn cerebe lac-deep coma
C0160198|T037|AB|851.76|ICD9CM|Opn cerebel lac-coma NOS|Opn cerebel lac-coma NOS
C0695224|T037|PT|851.79|ICD9CM|Cerebellar or brain stem laceration with open intracranial wound, with concussion, unspecified|Cerebellar or brain stem laceration with open intracranial wound, with concussion, unspecified
C0695224|T037|AB|851.79|ICD9CM|Opn cerebell lac-concuss|Opn cerebell lac-concuss
C0160200|T037|HT|851.8|ICD9CM|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound
C0160201|T037|AB|851.80|ICD9CM|Brain laceration NEC|Brain laceration NEC
C0160202|T037|AB|851.81|ICD9CM|Brain lacer NEC w/o coma|Brain lacer NEC w/o coma
C0160203|T037|AB|851.82|ICD9CM|Brain lac NEC-brief coma|Brain lac NEC-brief coma
C0160204|T037|AB|851.83|ICD9CM|Brain lacer NEC-mod coma|Brain lacer NEC-mod coma
C0160205|T037|AB|851.84|ICD9CM|Brain lac NEC-proln coma|Brain lac NEC-proln coma
C0160206|T037|AB|851.85|ICD9CM|Brain lac NEC-deep coma|Brain lac NEC-deep coma
C0160207|T037|AB|851.86|ICD9CM|Brain lacer NEC-coma NOS|Brain lacer NEC-coma NOS
C0695225|T037|AB|851.89|ICD9CM|Brain lacer NEC-concuss|Brain lacer NEC-concuss
C0160209|T037|HT|851.9|ICD9CM|Other and unspecified cerebral laceration and contusion, with open intracranial wound|Other and unspecified cerebral laceration and contusion, with open intracranial wound
C0160210|T037|AB|851.90|ICD9CM|Brain lac NEC w open wnd|Brain lac NEC w open wnd
C0160211|T037|AB|851.91|ICD9CM|Opn brain lacer w/o coma|Opn brain lacer w/o coma
C0160212|T037|AB|851.92|ICD9CM|Opn brain lac-brief coma|Opn brain lac-brief coma
C0160213|T037|AB|851.93|ICD9CM|Opn brain lacer-mod coma|Opn brain lacer-mod coma
C0160214|T037|AB|851.94|ICD9CM|Opn brain lac-proln coma|Opn brain lac-proln coma
C0160215|T037|AB|851.95|ICD9CM|Open brain lac-deep coma|Open brain lac-deep coma
C0160216|T037|AB|851.96|ICD9CM|Opn brain lacer-coma NOS|Opn brain lacer-coma NOS
C0695226|T037|AB|851.99|ICD9CM|Open brain lacer-concuss|Open brain lacer-concuss
C0160218|T046|HT|852|ICD9CM|Subarachnoid, subdural, and extradural hemorrhage, following injury|Subarachnoid, subdural, and extradural hemorrhage, following injury
C0160219|T046|HT|852.0|ICD9CM|Subarachnoid hemorrhage following injury without mention of open intracranial wound|Subarachnoid hemorrhage following injury without mention of open intracranial wound
C0160220|T037|AB|852.00|ICD9CM|Traum subarachnoid hem|Traum subarachnoid hem
C0160221|T037|AB|852.01|ICD9CM|Subarachnoid hem-no coma|Subarachnoid hem-no coma
C0160222|T037|AB|852.02|ICD9CM|Subarach hem-brief coma|Subarach hem-brief coma
C0160223|T037|AB|852.03|ICD9CM|Subarach hem-mod coma|Subarach hem-mod coma
C0160224|T037|AB|852.04|ICD9CM|Subarach hem-prolng coma|Subarach hem-prolng coma
C0160225|T037|AB|852.05|ICD9CM|Subarach hem-deep coma|Subarach hem-deep coma
C0160226|T037|AB|852.06|ICD9CM|Subarach hem-coma NOS|Subarach hem-coma NOS
C0160227|T037|AB|852.09|ICD9CM|Subarach hem-concussion|Subarach hem-concussion
C0160228|T037|HT|852.1|ICD9CM|Subarachnoid hemorrhage following injury with open intracranial wound|Subarachnoid hemorrhage following injury with open intracranial wound
C0160229|T037|AB|852.10|ICD9CM|Subarach hem w opn wound|Subarach hem w opn wound
C0160230|T037|AB|852.11|ICD9CM|Opn subarach hem-no coma|Opn subarach hem-no coma
C0160230|T037|PT|852.11|ICD9CM|Subarachnoid hemorrhage following injury with open intracranial wound, with no loss of consciousness|Subarachnoid hemorrhage following injury with open intracranial wound, with no loss of consciousness
C0160231|T037|AB|852.12|ICD9CM|Op subarach hem-brf coma|Op subarach hem-brf coma
C0160232|T037|AB|852.13|ICD9CM|Op subarach hem-mod coma|Op subarach hem-mod coma
C0160233|T037|AB|852.14|ICD9CM|Op subarach hem-prol com|Op subarach hem-prol com
C0160234|T037|AB|852.15|ICD9CM|Op subarach hem-deep com|Op subarach hem-deep com
C0160235|T037|AB|852.16|ICD9CM|Op subarach hem-coma NOS|Op subarach hem-coma NOS
C0273088|T037|AB|852.19|ICD9CM|Opn subarach hem-concuss|Opn subarach hem-concuss
C0273088|T037|PT|852.19|ICD9CM|Subarachnoid hemorrhage following injury with open intracranial wound, with concussion, unspecified|Subarachnoid hemorrhage following injury with open intracranial wound, with concussion, unspecified
C0160237|T046|HT|852.2|ICD9CM|Subdural hemorrhage following injury without mention of open intracranial wound|Subdural hemorrhage following injury without mention of open intracranial wound
C0160238|T037|AB|852.20|ICD9CM|Traumatic subdural hem|Traumatic subdural hem
C0160239|T037|AB|852.21|ICD9CM|Subdural hem w/o coma|Subdural hem w/o coma
C0160240|T037|AB|852.22|ICD9CM|Subdural hem-brief coma|Subdural hem-brief coma
C0160241|T037|AB|852.23|ICD9CM|Subdural hemorr-mod coma|Subdural hemorr-mod coma
C0160242|T037|AB|852.24|ICD9CM|Subdural hem-prolng coma|Subdural hem-prolng coma
C0160243|T037|AB|852.25|ICD9CM|Subdural hem-deep coma|Subdural hem-deep coma
C0160244|T037|AB|852.26|ICD9CM|Subdural hemorr-coma NOS|Subdural hemorr-coma NOS
C0160245|T037|AB|852.29|ICD9CM|Subdural hem-concussion|Subdural hem-concussion
C0160246|T037|HT|852.3|ICD9CM|Subdural hemorrhage following injury, with open intracranial wound|Subdural hemorrhage following injury, with open intracranial wound
C0160247|T037|AB|852.30|ICD9CM|Subdural hem w opn wound|Subdural hem w opn wound
C0160248|T046|AB|852.31|ICD9CM|Open subdur hem w/o coma|Open subdur hem w/o coma
C0160248|T046|PT|852.31|ICD9CM|Subdural hemorrhage following injury with open intracranial wound, with no loss of consciousness|Subdural hemorrhage following injury with open intracranial wound, with no loss of consciousness
C0160249|T037|AB|852.32|ICD9CM|Opn subdur hem-brf coma|Opn subdur hem-brf coma
C0160250|T037|AB|852.33|ICD9CM|Opn subdur hem-mod coma|Opn subdur hem-mod coma
C0160251|T037|AB|852.34|ICD9CM|Opn subdur hem-prol coma|Opn subdur hem-prol coma
C0160252|T037|AB|852.35|ICD9CM|Opn subdur hem-deep coma|Opn subdur hem-deep coma
C0160253|T037|AB|852.36|ICD9CM|Opn subdur hem-coma NOS|Opn subdur hem-coma NOS
C0273097|T037|AB|852.39|ICD9CM|Opn subdur hem-concuss|Opn subdur hem-concuss
C0273097|T037|PT|852.39|ICD9CM|Subdural hemorrhage following injury with open intracranial wound, with concussion, unspecified|Subdural hemorrhage following injury with open intracranial wound, with concussion, unspecified
C0160255|T037|HT|852.4|ICD9CM|Extradural hemorrhage following injury without mention of open intracranial wound|Extradural hemorrhage following injury without mention of open intracranial wound
C0273099|T037|AB|852.40|ICD9CM|Traumatic extradural hem|Traumatic extradural hem
C0273100|T037|AB|852.41|ICD9CM|Extradural hem w/o coma|Extradural hem w/o coma
C0160258|T037|AB|852.42|ICD9CM|Extradur hem-brief coma|Extradur hem-brief coma
C0160259|T037|AB|852.43|ICD9CM|Extradural hem-mod coma|Extradural hem-mod coma
C0160260|T037|AB|852.44|ICD9CM|Extradur hem-proln coma|Extradur hem-proln coma
C0273104|T037|AB|852.45|ICD9CM|Extradural hem-deep coma|Extradural hem-deep coma
C0273104|T037|AB|852.46|ICD9CM|Extradural hem-coma NOS|Extradural hem-coma NOS
C0160263|T037|AB|852.49|ICD9CM|Extadural hem-concuss|Extadural hem-concuss
C0160264|T037|HT|852.5|ICD9CM|Extradural hemorrhage following injury with open intracranial wound|Extradural hemorrhage following injury with open intracranial wound
C0160265|T037|AB|852.50|ICD9CM|Extradural hem w opn wnd|Extradural hem w opn wnd
C0160266|T037|AB|852.51|ICD9CM|Extradural hemor-no coma|Extradural hemor-no coma
C0160266|T037|PT|852.51|ICD9CM|Extradural hemorrhage following injury with open intracranial wound, with no loss of consciousness|Extradural hemorrhage following injury with open intracranial wound, with no loss of consciousness
C0160267|T037|AB|852.52|ICD9CM|Extradur hem-brief coma|Extradur hem-brief coma
C0160268|T037|AB|852.53|ICD9CM|Extradural hem-mod coma|Extradural hem-mod coma
C0160269|T037|AB|852.54|ICD9CM|Extradur hem-proln coma|Extradur hem-proln coma
C0160270|T037|AB|852.55|ICD9CM|Extradur hem-deep coma|Extradur hem-deep coma
C0160271|T037|AB|852.56|ICD9CM|Extradural hem-coma NOS|Extradural hem-coma NOS
C0273106|T037|AB|852.59|ICD9CM|Extradural hem-concuss|Extradural hem-concuss
C0273106|T037|PT|852.59|ICD9CM|Extradural hemorrhage following injury with open intracranial wound, with concussion, unspecified|Extradural hemorrhage following injury with open intracranial wound, with concussion, unspecified
C0160273|T046|HT|853|ICD9CM|Other and unspecified intracranial hemorrhage following injury|Other and unspecified intracranial hemorrhage following injury
C0160275|T037|AB|853.00|ICD9CM|Traumatic brain hem NEC|Traumatic brain hem NEC
C0160276|T037|AB|853.01|ICD9CM|Brain hem NEC w/o coma|Brain hem NEC w/o coma
C0160277|T037|AB|853.02|ICD9CM|Brain hem NEC-brief coma|Brain hem NEC-brief coma
C0160278|T037|AB|853.03|ICD9CM|Brain hem NEC-mod coma|Brain hem NEC-mod coma
C0160279|T037|AB|853.04|ICD9CM|Brain hem NEC-proln coma|Brain hem NEC-proln coma
C0160280|T037|AB|853.05|ICD9CM|Brain hem NEC-deep coma|Brain hem NEC-deep coma
C0160281|T037|AB|853.06|ICD9CM|Brain hem NEC-coma NOS|Brain hem NEC-coma NOS
C0475036|T047|AB|853.09|ICD9CM|Brain hem NEC-concussion|Brain hem NEC-concussion
C0160283|T046|HT|853.1|ICD9CM|Other and unspecified intracranial hemorrhage following injury with open intracranial wound|Other and unspecified intracranial hemorrhage following injury with open intracranial wound
C0160284|T037|AB|853.10|ICD9CM|Brain hem NEC w opn wnd|Brain hem NEC w opn wnd
C0160285|T037|AB|853.11|ICD9CM|Brain hem opn w/o coma|Brain hem opn w/o coma
C0160286|T037|AB|853.12|ICD9CM|Brain hem opn-brf coma|Brain hem opn-brf coma
C0160287|T037|AB|853.13|ICD9CM|Brain hem open-mod coma|Brain hem open-mod coma
C0160288|T037|AB|853.14|ICD9CM|Brain hem opn-proln coma|Brain hem opn-proln coma
C0160289|T037|AB|853.15|ICD9CM|Brain hem open-deep coma|Brain hem open-deep coma
C0160290|T037|AB|853.16|ICD9CM|Brain hem open-coma NOS|Brain hem open-coma NOS
C0475045|T037|AB|853.19|ICD9CM|Brain hem opn-concussion|Brain hem opn-concussion
C0160292|T037|HT|854|ICD9CM|Intracranial injury of other and unspecified nature|Intracranial injury of other and unspecified nature
C0021878|T037|HT|854.0|ICD9CM|Intracranial injury of other and unspecified nature without mention of open intracranial wound|Intracranial injury of other and unspecified nature without mention of open intracranial wound
C0021879|T037|AB|854.00|ICD9CM|Brain injury NEC|Brain injury NEC
C0160293|T037|AB|854.01|ICD9CM|Brain injury NEC-no coma|Brain injury NEC-no coma
C0160294|T037|AB|854.02|ICD9CM|Brain inj NEC-brief coma|Brain inj NEC-brief coma
C0160295|T037|AB|854.03|ICD9CM|Brain inj NEC-mod coma|Brain inj NEC-mod coma
C0160296|T037|AB|854.04|ICD9CM|Brain inj NEC-proln coma|Brain inj NEC-proln coma
C0160297|T037|AB|854.05|ICD9CM|Brain inj NEC-deep coma|Brain inj NEC-deep coma
C0160298|T037|AB|854.06|ICD9CM|Brain inj NEC-coma NOS|Brain inj NEC-coma NOS
C0160299|T037|AB|854.09|ICD9CM|Brain inj NEC-concussion|Brain inj NEC-concussion
C0160300|T037|HT|854.1|ICD9CM|Intracranial injury of other and unspecified nature with open intracranial wound|Intracranial injury of other and unspecified nature with open intracranial wound
C0160301|T037|AB|854.10|ICD9CM|Brain injury w opn wnd|Brain injury w opn wnd
C0160302|T037|AB|854.11|ICD9CM|Opn brain inj w/o coma|Opn brain inj w/o coma
C0160303|T037|AB|854.12|ICD9CM|Opn brain inj-brief coma|Opn brain inj-brief coma
C0160304|T037|AB|854.13|ICD9CM|Opn brain inj-mod coma|Opn brain inj-mod coma
C0160305|T037|AB|854.14|ICD9CM|Opn brain inj-proln coma|Opn brain inj-proln coma
C0160306|T037|AB|854.15|ICD9CM|Opn brain inj-deep coma|Opn brain inj-deep coma
C0160307|T037|AB|854.16|ICD9CM|Open brain inj-coma NOS|Open brain inj-coma NOS
C0160308|T037|AB|854.19|ICD9CM|Opn brain inj-concussion|Opn brain inj-concussion
C0340008|T037|HT|860|ICD9CM|Traumatic pneumothorax and hemothorax|Traumatic pneumothorax and hemothorax
C0376106|T037|HT|860-869.99|ICD9CM|INTERNAL INJURY OF THORAX, ABDOMEN, AND PELVIS|INTERNAL INJURY OF THORAX, ABDOMEN, AND PELVIS
C0347620|T037|AB|860.0|ICD9CM|Traum pneumothorax-close|Traum pneumothorax-close
C0347620|T037|PT|860.0|ICD9CM|Traumatic pneumothorax without mention of open wound into thorax|Traumatic pneumothorax without mention of open wound into thorax
C0347619|T037|AB|860.1|ICD9CM|Traum pneumothorax-open|Traum pneumothorax-open
C0347619|T037|PT|860.1|ICD9CM|Traumatic pneumothorax with open wound into thorax|Traumatic pneumothorax with open wound into thorax
C0160312|T037|AB|860.2|ICD9CM|Traum hemothorax-closed|Traum hemothorax-closed
C0160312|T037|PT|860.2|ICD9CM|Traumatic hemothorax without mention of open wound into thorax|Traumatic hemothorax without mention of open wound into thorax
C0347621|T037|AB|860.3|ICD9CM|Traum hemothorax-open|Traum hemothorax-open
C0347621|T037|PT|860.3|ICD9CM|Traumatic hemothorax with open wound into thorax|Traumatic hemothorax with open wound into thorax
C0347624|T047|AB|860.4|ICD9CM|Traum pneumohemothor-cl|Traum pneumohemothor-cl
C0347624|T047|PT|860.4|ICD9CM|Traumatic pneumohemothorax without mention of open wound into thorax|Traumatic pneumohemothorax without mention of open wound into thorax
C0347623|T047|AB|860.5|ICD9CM|Traum pneumohemothor-opn|Traum pneumohemothor-opn
C0347623|T047|PT|860.5|ICD9CM|Traumatic pneumohemothorax with open wound into thorax|Traumatic pneumohemothorax with open wound into thorax
C0160316|T037|HT|861|ICD9CM|Injury to heart and lung|Injury to heart and lung
C0160318|T037|HT|861.0|ICD9CM|Heart injury, without mention of open wound into thorax|Heart injury, without mention of open wound into thorax
C0160318|T037|AB|861.00|ICD9CM|Heart injury NOS-closed|Heart injury NOS-closed
C0160318|T037|PT|861.00|ICD9CM|Unspecified injury of heart without mention of open wound into thorax|Unspecified injury of heart without mention of open wound into thorax
C0160319|T037|PT|861.01|ICD9CM|Contusion of heart without mention of open wound into thorax|Contusion of heart without mention of open wound into thorax
C0160319|T037|AB|861.01|ICD9CM|Heart contusion-closed|Heart contusion-closed
C0160320|T037|AB|861.02|ICD9CM|Heart laceration-closed|Heart laceration-closed
C0160321|T037|AB|861.03|ICD9CM|Heart chamber lacerat-cl|Heart chamber lacerat-cl
C0160321|T037|PT|861.03|ICD9CM|Laceration of heart with penetration of heart chambers without mention of open wound into thorax|Laceration of heart with penetration of heart chambers without mention of open wound into thorax
C0160323|T037|HT|861.1|ICD9CM|Heart injury, with open wound into thorax|Heart injury, with open wound into thorax
C0160323|T037|AB|861.10|ICD9CM|Heart injury NOS-open|Heart injury NOS-open
C0160323|T037|PT|861.10|ICD9CM|Unspecified injury of heart with open wound into thorax|Unspecified injury of heart with open wound into thorax
C0160324|T037|PT|861.11|ICD9CM|Contusion of heart with open wound into thorax|Contusion of heart with open wound into thorax
C0160324|T037|AB|861.11|ICD9CM|Heart contusion-open|Heart contusion-open
C0160325|T037|AB|861.12|ICD9CM|Heart laceration-open|Heart laceration-open
C0160325|T037|PT|861.12|ICD9CM|Laceration of heart without penetration of heart chambers, with open wound into thorax|Laceration of heart without penetration of heart chambers, with open wound into thorax
C0160326|T037|AB|861.13|ICD9CM|Heart chamber lacer-opn|Heart chamber lacer-opn
C0160326|T037|PT|861.13|ICD9CM|Laceration of heart with penetration of heart chambers with open wound into thorax|Laceration of heart with penetration of heart chambers with open wound into thorax
C0160328|T037|HT|861.2|ICD9CM|Lung injury, without mention of open wound into thorax|Lung injury, without mention of open wound into thorax
C0160328|T037|AB|861.20|ICD9CM|Lung injury NOS-closed|Lung injury NOS-closed
C0160328|T037|PT|861.20|ICD9CM|Unspecified injury of lung without mention of open wound into thorax|Unspecified injury of lung without mention of open wound into thorax
C0160329|T037|PT|861.21|ICD9CM|Contusion of lung without mention of open wound into thorax|Contusion of lung without mention of open wound into thorax
C0160329|T037|AB|861.21|ICD9CM|Lung contusion-closed|Lung contusion-closed
C0160330|T037|PT|861.22|ICD9CM|Laceration of lung without mention of open wound into thorax|Laceration of lung without mention of open wound into thorax
C0160330|T037|AB|861.22|ICD9CM|Lung laceration-closed|Lung laceration-closed
C0160332|T037|HT|861.3|ICD9CM|Lung injury, with open wound into thorax|Lung injury, with open wound into thorax
C0160332|T037|AB|861.30|ICD9CM|Lung injury NOS-open|Lung injury NOS-open
C0160332|T037|PT|861.30|ICD9CM|Unspecified injury of lung with open wound into thorax|Unspecified injury of lung with open wound into thorax
C0160333|T037|PT|861.31|ICD9CM|Contusion of lung with open wound into thorax|Contusion of lung with open wound into thorax
C0160333|T037|AB|861.31|ICD9CM|Lung contusion-open|Lung contusion-open
C0160334|T037|PT|861.32|ICD9CM|Laceration of lung with open wound into thorax|Laceration of lung with open wound into thorax
C0160334|T037|AB|861.32|ICD9CM|Lung laceration-open|Lung laceration-open
C0160335|T037|HT|862|ICD9CM|Injury to other and unspecified intrathoracic organs|Injury to other and unspecified intrathoracic organs
C0021505|T037|AB|862.0|ICD9CM|Diaphragm injury-closed|Diaphragm injury-closed
C0021505|T037|PT|862.0|ICD9CM|Injury to diaphragm, without mention of open wound into cavity|Injury to diaphragm, without mention of open wound into cavity
C0160336|T037|AB|862.1|ICD9CM|Diaphragm injury-open|Diaphragm injury-open
C0160336|T037|PT|862.1|ICD9CM|Injury to diaphragm, with open wound into cavity|Injury to diaphragm, with open wound into cavity
C0160337|T037|HT|862.2|ICD9CM|Injury to other specified intrathoracic organs without mention of open wound into cavity|Injury to other specified intrathoracic organs without mention of open wound into cavity
C0160338|T037|AB|862.21|ICD9CM|Bronchus injury-closed|Bronchus injury-closed
C0160338|T037|PT|862.21|ICD9CM|Injury to bronchus without mention of open wound into cavity|Injury to bronchus without mention of open wound into cavity
C1318512|T037|AB|862.22|ICD9CM|Esophagus injury-closed|Esophagus injury-closed
C1318512|T037|PT|862.22|ICD9CM|Injury to esophagus without mention of open wound into cavity|Injury to esophagus without mention of open wound into cavity
C0160337|T037|PT|862.29|ICD9CM|Injury to other specified intrathoracic organs without mention of open wound into cavity|Injury to other specified intrathoracic organs without mention of open wound into cavity
C0160337|T037|AB|862.29|ICD9CM|Intrathoracic inj NEC-cl|Intrathoracic inj NEC-cl
C0160340|T037|HT|862.3|ICD9CM|Injury to other specified intrathoracic organs with open wound into cavity|Injury to other specified intrathoracic organs with open wound into cavity
C0160341|T037|AB|862.31|ICD9CM|Bronchus injury-open|Bronchus injury-open
C0160341|T037|PT|862.31|ICD9CM|Injury to bronchus with open wound into cavity|Injury to bronchus with open wound into cavity
C0160342|T037|AB|862.32|ICD9CM|Esophagus injury-open|Esophagus injury-open
C0160342|T037|PT|862.32|ICD9CM|Injury to esophagus with open wound into cavity|Injury to esophagus with open wound into cavity
C0160340|T037|PT|862.39|ICD9CM|Injury to other specified intrathoracic organs with open wound into cavity|Injury to other specified intrathoracic organs with open wound into cavity
C0160340|T037|AB|862.39|ICD9CM|Intrathorac inj NEC-open|Intrathorac inj NEC-open
C0160343|T037|PT|862.8|ICD9CM|Injury to multiple and unspecified intrathoracic organs, without mention of open wound into cavity|Injury to multiple and unspecified intrathoracic organs, without mention of open wound into cavity
C0160343|T037|AB|862.8|ICD9CM|Intrathoracic inj NOS-cl|Intrathoracic inj NOS-cl
C0273127|T037|PT|862.9|ICD9CM|Injury to multiple and unspecified intrathoracic organs, with open wound into cavity|Injury to multiple and unspecified intrathoracic organs, with open wound into cavity
C0273127|T037|AB|862.9|ICD9CM|Intrathorac inj NOS-open|Intrathorac inj NOS-open
C0160345|T037|HT|863|ICD9CM|Injury to gastrointestinal tract|Injury to gastrointestinal tract
C0160346|T037|PT|863.0|ICD9CM|Injury to stomach, without mention of open wound into cavity|Injury to stomach, without mention of open wound into cavity
C0160346|T037|AB|863.0|ICD9CM|Stomach injury-closed|Stomach injury-closed
C0160347|T037|PT|863.1|ICD9CM|Injury to stomach, with open wound into cavity|Injury to stomach, with open wound into cavity
C0160347|T037|AB|863.1|ICD9CM|Stomach injury-open|Stomach injury-open
C0160348|T037|HT|863.2|ICD9CM|Injury to small intestine without mention of open wound into cavity|Injury to small intestine without mention of open wound into cavity
C0160349|T037|PT|863.20|ICD9CM|Injury to small intestine, unspecified site, without open wound into cavity|Injury to small intestine, unspecified site, without open wound into cavity
C0160349|T037|AB|863.20|ICD9CM|Small intest inj NOS-cl|Small intest inj NOS-cl
C0160350|T037|AB|863.21|ICD9CM|Duodenum injury-closed|Duodenum injury-closed
C0160350|T037|PT|863.21|ICD9CM|Injury to duodenum, without open wound into cavity|Injury to duodenum, without open wound into cavity
C0160351|T037|PT|863.29|ICD9CM|Other injury to small intestine, without mention of open wound into cavity|Other injury to small intestine, without mention of open wound into cavity
C0160351|T037|AB|863.29|ICD9CM|Small intest inj NEC-cl|Small intest inj NEC-cl
C0160352|T037|HT|863.3|ICD9CM|Injury to small intestine with open wound into cavity|Injury to small intestine with open wound into cavity
C0160353|T037|PT|863.30|ICD9CM|Injury to small intestine, unspecified site, with open wound into cavity|Injury to small intestine, unspecified site, with open wound into cavity
C0160353|T037|AB|863.30|ICD9CM|Small intest inj NOS-opn|Small intest inj NOS-opn
C0160354|T037|AB|863.31|ICD9CM|Duodenum injury-open|Duodenum injury-open
C0160354|T037|PT|863.31|ICD9CM|Injury to duodenum, with open wound into cavity|Injury to duodenum, with open wound into cavity
C0160355|T037|PT|863.39|ICD9CM|Other injury to small intestine, with open wound into cavity|Other injury to small intestine, with open wound into cavity
C0160355|T037|AB|863.39|ICD9CM|Small intest inj NEC-opn|Small intest inj NEC-opn
C0160356|T037|HT|863.4|ICD9CM|Injury to colon or rectum without mention of open wound into cavity|Injury to colon or rectum without mention of open wound into cavity
C0160357|T037|AB|863.40|ICD9CM|Colon injury NOS-closed|Colon injury NOS-closed
C0160357|T037|PT|863.40|ICD9CM|Injury to colon, unspecified site, without mention of open wound into cavity|Injury to colon, unspecified site, without mention of open wound into cavity
C0160358|T037|AB|863.41|ICD9CM|Ascending colon inj-clos|Ascending colon inj-clos
C0160358|T037|PT|863.41|ICD9CM|Injury to ascending [right] colon, without mention of open wound into cavity|Injury to ascending [right] colon, without mention of open wound into cavity
C0160359|T037|PT|863.42|ICD9CM|Injury to transverse colon, without mention of open wound into cavity|Injury to transverse colon, without mention of open wound into cavity
C0160359|T037|AB|863.42|ICD9CM|Transverse colon inj-cl|Transverse colon inj-cl
C0160360|T037|AB|863.43|ICD9CM|Descending colon inj-cl|Descending colon inj-cl
C0160360|T037|PT|863.43|ICD9CM|Injury to descending [left] colon, without mention of open wound into cavity|Injury to descending [left] colon, without mention of open wound into cavity
C0160361|T037|PT|863.44|ICD9CM|Injury to sigmoid colon, without mention of open wound into cavity|Injury to sigmoid colon, without mention of open wound into cavity
C0160361|T037|AB|863.44|ICD9CM|Sigmoid colon inj-closed|Sigmoid colon inj-closed
C0160362|T037|PT|863.45|ICD9CM|Injury to rectum, without mention of open wound into cavity|Injury to rectum, without mention of open wound into cavity
C0160362|T037|AB|863.45|ICD9CM|Rectum injury-closed|Rectum injury-closed
C0160363|T037|AB|863.46|ICD9CM|Colon inj mult site-clos|Colon inj mult site-clos
C0160363|T037|PT|863.46|ICD9CM|Injury to multiple sites in colon and rectum, without mention of open wound into cavity|Injury to multiple sites in colon and rectum, without mention of open wound into cavity
C0434062|T037|AB|863.49|ICD9CM|Colon injury NEC-closed|Colon injury NEC-closed
C0434062|T037|PT|863.49|ICD9CM|Other injury to colon or rectum, without mention of open wound into cavity|Other injury to colon or rectum, without mention of open wound into cavity
C0160365|T037|HT|863.5|ICD9CM|Injury to colon or rectum with open wound into cavity|Injury to colon or rectum with open wound into cavity
C0160366|T037|AB|863.50|ICD9CM|Colon injury NOS-open|Colon injury NOS-open
C0160366|T037|PT|863.50|ICD9CM|Injury to colon, unspecified site, with open wound into cavity|Injury to colon, unspecified site, with open wound into cavity
C0160367|T037|AB|863.51|ICD9CM|Ascending colon inj-open|Ascending colon inj-open
C0160367|T037|PT|863.51|ICD9CM|Injury to ascending [right] colon, with open wound into cavity|Injury to ascending [right] colon, with open wound into cavity
C0160368|T037|PT|863.52|ICD9CM|Injury to transverse colon, with open wound into cavity|Injury to transverse colon, with open wound into cavity
C0160368|T037|AB|863.52|ICD9CM|Transverse colon inj-opn|Transverse colon inj-opn
C0160369|T037|AB|863.53|ICD9CM|Descending colon inj-opn|Descending colon inj-opn
C0160369|T037|PT|863.53|ICD9CM|Injury to descending [left] colon, with open wound into cavity|Injury to descending [left] colon, with open wound into cavity
C0160370|T037|PT|863.54|ICD9CM|Injury to sigmoid colon, with open wound into cavity|Injury to sigmoid colon, with open wound into cavity
C0160370|T037|AB|863.54|ICD9CM|Sigmoid colon inj-open|Sigmoid colon inj-open
C0160371|T037|PT|863.55|ICD9CM|Injury to rectum, with open wound into cavity|Injury to rectum, with open wound into cavity
C0160371|T037|AB|863.55|ICD9CM|Rectum injury-open|Rectum injury-open
C0160372|T037|AB|863.56|ICD9CM|Colon inj mult site-open|Colon inj mult site-open
C0160372|T037|PT|863.56|ICD9CM|Injury to multiple sites in colon and rectum, with open wound into cavity|Injury to multiple sites in colon and rectum, with open wound into cavity
C0434058|T037|AB|863.59|ICD9CM|Colon injury NEC-open|Colon injury NEC-open
C0434058|T037|PT|863.59|ICD9CM|Other injury to colon or rectum, with open wound into cavity|Other injury to colon or rectum, with open wound into cavity
C0160374|T037|HT|863.8|ICD9CM|Injury to other and unspecified gastrointestinal sites without mention of open wound into cavity|Injury to other and unspecified gastrointestinal sites without mention of open wound into cavity
C0160375|T037|AB|863.80|ICD9CM|GI injury NOS-closed|GI injury NOS-closed
C0160375|T037|PT|863.80|ICD9CM|Injury to gastrointestinal tract, unspecified site, without mention of open wound into cavity|Injury to gastrointestinal tract, unspecified site, without mention of open wound into cavity
C0273164|T037|PT|863.81|ICD9CM|Injury to pancreas, head, without mention of open wound into cavity|Injury to pancreas, head, without mention of open wound into cavity
C0273164|T037|AB|863.81|ICD9CM|Pancreas, head inj-close|Pancreas, head inj-close
C0160377|T037|PT|863.82|ICD9CM|Injury to pancreas, body, without mention of open wound into cavity|Injury to pancreas, body, without mention of open wound into cavity
C0160377|T037|AB|863.82|ICD9CM|Pancreas, body inj-close|Pancreas, body inj-close
C0160378|T037|PT|863.83|ICD9CM|Injury to pancreas, tail, without mention of open wound into cavity|Injury to pancreas, tail, without mention of open wound into cavity
C0160378|T037|AB|863.83|ICD9CM|Pancreas, tail inj-close|Pancreas, tail inj-close
C0160379|T037|PT|863.84|ICD9CM|Injury to pancreas, multiple and unspecified sites, without mention of open wound into cavity|Injury to pancreas, multiple and unspecified sites, without mention of open wound into cavity
C0160379|T037|AB|863.84|ICD9CM|Pancreas injury NOS-clos|Pancreas injury NOS-clos
C0160380|T037|AB|863.85|ICD9CM|Appendix injury-closed|Appendix injury-closed
C0160380|T037|PT|863.85|ICD9CM|Injury to appendix, without mention of open wound into cavity|Injury to appendix, without mention of open wound into cavity
C0160381|T037|AB|863.89|ICD9CM|GI injury NEC-closed|GI injury NEC-closed
C0160381|T037|PT|863.89|ICD9CM|Injury to other gastrointestinal sites, without mention of open wound into cavity|Injury to other gastrointestinal sites, without mention of open wound into cavity
C0160389|T037|HT|863.9|ICD9CM|Injury to other and unspecified gastrointestinal sites, with open wound into cavity|Injury to other and unspecified gastrointestinal sites, with open wound into cavity
C0160383|T037|AB|863.90|ICD9CM|GI injury NOS-open|GI injury NOS-open
C0160383|T037|PT|863.90|ICD9CM|Injury to gastrointestinal tract, unspecified site, with open wound into cavity|Injury to gastrointestinal tract, unspecified site, with open wound into cavity
C0160384|T037|PT|863.91|ICD9CM|Injury to pancreas, head, with open wound into cavity|Injury to pancreas, head, with open wound into cavity
C0160384|T037|AB|863.91|ICD9CM|Pancreas, head inj-open|Pancreas, head inj-open
C0160385|T037|PT|863.92|ICD9CM|Injury to pancreas, body, with open wound into cavity|Injury to pancreas, body, with open wound into cavity
C0160385|T037|AB|863.92|ICD9CM|Pancreas, body inj-open|Pancreas, body inj-open
C0160386|T037|PT|863.93|ICD9CM|Injury to pancreas, tail, with open wound into cavity|Injury to pancreas, tail, with open wound into cavity
C0160386|T037|AB|863.93|ICD9CM|Pancreas, tail inj-open|Pancreas, tail inj-open
C0160387|T037|PT|863.94|ICD9CM|Injury to pancreas, multiple and unspecified sites, with open wound into cavity|Injury to pancreas, multiple and unspecified sites, with open wound into cavity
C0160387|T037|AB|863.94|ICD9CM|Pancreas injury NOS-open|Pancreas injury NOS-open
C0160388|T037|AB|863.95|ICD9CM|Appendix injury-open|Appendix injury-open
C0160388|T037|PT|863.95|ICD9CM|Injury to appendix, with open wound into cavity|Injury to appendix, with open wound into cavity
C0160389|T037|AB|863.99|ICD9CM|GI injury NEC-open|GI injury NEC-open
C0160389|T037|PT|863.99|ICD9CM|Injury to other gastrointestinal sites, with open wound into cavity|Injury to other gastrointestinal sites, with open wound into cavity
C0160390|T037|HT|864|ICD9CM|Injury to liver|Injury to liver
C0160392|T037|HT|864.0|ICD9CM|Injury to liver without mention of open wound into cavity|Injury to liver without mention of open wound into cavity
C0160392|T037|PT|864.00|ICD9CM|Injury to liver without mention of open wound into cavity, unspecified injury|Injury to liver without mention of open wound into cavity, unspecified injury
C0160392|T037|AB|864.00|ICD9CM|Liver injury NOS-closed|Liver injury NOS-closed
C0160393|T037|PT|864.01|ICD9CM|Injury to liver without mention of open wound into cavity, hematoma and contusion|Injury to liver without mention of open wound into cavity, hematoma and contusion
C0160393|T037|AB|864.01|ICD9CM|Liver hematoma/contusion|Liver hematoma/contusion
C0160394|T037|PT|864.02|ICD9CM|Injury to liver without mention of open wound into cavity, laceration, minor|Injury to liver without mention of open wound into cavity, laceration, minor
C0160394|T037|AB|864.02|ICD9CM|Liver laceration, minor|Liver laceration, minor
C0273175|T037|PT|864.03|ICD9CM|Injury to liver without mention of open wound into cavity, laceration, moderate|Injury to liver without mention of open wound into cavity, laceration, moderate
C0273175|T037|AB|864.03|ICD9CM|Liver laceration, mod|Liver laceration, mod
C0160396|T037|PT|864.04|ICD9CM|Injury to liver without mention of open wound into cavity, laceration, major|Injury to liver without mention of open wound into cavity, laceration, major
C0160396|T037|AB|864.04|ICD9CM|Liver laceration, major|Liver laceration, major
C0375639|T037|PT|864.05|ICD9CM|Injury to liver without mention of open wound into cavity laceration, unspecified|Injury to liver without mention of open wound into cavity laceration, unspecified
C0375639|T037|AB|864.05|ICD9CM|Liver lacerat unspcf cls|Liver lacerat unspcf cls
C0160397|T037|AB|864.09|ICD9CM|Liver injury NEC-closed|Liver injury NEC-closed
C0160397|T037|PT|864.09|ICD9CM|Other injury to liver without mention of open wound into cavity|Other injury to liver without mention of open wound into cavity
C0160399|T037|HT|864.1|ICD9CM|Injury to liver with open wound into cavity|Injury to liver with open wound into cavity
C0160399|T037|PT|864.10|ICD9CM|Injury to liver with open wound into cavity, unspecified injury|Injury to liver with open wound into cavity, unspecified injury
C0160399|T037|AB|864.10|ICD9CM|Liver injury NOS-open|Liver injury NOS-open
C0160400|T037|PT|864.11|ICD9CM|Injury to liver with open wound into cavity, hematoma and contusion|Injury to liver with open wound into cavity, hematoma and contusion
C0160400|T037|AB|864.11|ICD9CM|Liver hematom/contus-opn|Liver hematom/contus-opn
C0160401|T037|PT|864.12|ICD9CM|Injury to liver with open wound into cavity, laceration, minor|Injury to liver with open wound into cavity, laceration, minor
C0160401|T037|AB|864.12|ICD9CM|Liver lacerat, minor-opn|Liver lacerat, minor-opn
C0160402|T037|PT|864.13|ICD9CM|Injury to liver with open wound into cavity, laceration, moderate|Injury to liver with open wound into cavity, laceration, moderate
C0160402|T037|AB|864.13|ICD9CM|Liver lacerat, mod-open|Liver lacerat, mod-open
C0273182|T037|PT|864.14|ICD9CM|Injury to liver with open wound into cavity, laceration, major|Injury to liver with open wound into cavity, laceration, major
C0273182|T037|AB|864.14|ICD9CM|Liver lacerat, major-opn|Liver lacerat, major-opn
C0859268|T037|PT|864.15|ICD9CM|Injury to liver with open wound into cavity, laceration, unspecified|Injury to liver with open wound into cavity, laceration, unspecified
C0859268|T037|AB|864.15|ICD9CM|Liver lacerat unspcf opn|Liver lacerat unspcf opn
C0160404|T037|AB|864.19|ICD9CM|Liver injury NEC-open|Liver injury NEC-open
C0160404|T037|PT|864.19|ICD9CM|Other injury to liver with open wound into cavity|Other injury to liver with open wound into cavity
C0160405|T037|HT|865|ICD9CM|Injury to spleen|Injury to spleen
C0160407|T037|HT|865.0|ICD9CM|Injury to spleen without mention of open wound into cavity|Injury to spleen without mention of open wound into cavity
C0160407|T037|PT|865.00|ICD9CM|Injury to spleen without mention of open wound into cavity, unspecified injury|Injury to spleen without mention of open wound into cavity, unspecified injury
C0160407|T037|AB|865.00|ICD9CM|Spleen injury NOS-closed|Spleen injury NOS-closed
C0160408|T046|PT|865.01|ICD9CM|Injury to spleen without mention of open wound into cavity, hematoma without rupture of capsule|Injury to spleen without mention of open wound into cavity, hematoma without rupture of capsule
C0160408|T046|AB|865.01|ICD9CM|Spleen hematoma-closed|Spleen hematoma-closed
C0160409|T037|AB|865.02|ICD9CM|Spleen capsular tear|Spleen capsular tear
C0160410|T037|PT|865.03|ICD9CM|Injury to spleen without mention of open wound into cavity, laceration extending into parenchyma|Injury to spleen without mention of open wound into cavity, laceration extending into parenchyma
C0160410|T037|AB|865.03|ICD9CM|Spleen parenchyma lacer|Spleen parenchyma lacer
C0160411|T037|PT|865.04|ICD9CM|Injury to spleen without mention of open wound into cavity, massive parenchymal disruption|Injury to spleen without mention of open wound into cavity, massive parenchymal disruption
C0160411|T037|AB|865.04|ICD9CM|Spleen disruption-clos|Spleen disruption-clos
C0160412|T037|PT|865.09|ICD9CM|Other injury into spleen without mention of open wound into cavity|Other injury into spleen without mention of open wound into cavity
C0160412|T037|AB|865.09|ICD9CM|Spleen injury NEC-closed|Spleen injury NEC-closed
C0160414|T037|HT|865.1|ICD9CM|Injury to spleen with open wound into cavity|Injury to spleen with open wound into cavity
C0160414|T037|PT|865.10|ICD9CM|Injury to spleen with open wound into cavity, unspecified injury|Injury to spleen with open wound into cavity, unspecified injury
C0160414|T037|AB|865.10|ICD9CM|Spleen injury NOS-open|Spleen injury NOS-open
C0160415|T037|PT|865.11|ICD9CM|Injury to spleen with open wound into cavity, hematoma without rupture of capsule|Injury to spleen with open wound into cavity, hematoma without rupture of capsule
C0160415|T037|AB|865.11|ICD9CM|Spleen hematoma-open|Spleen hematoma-open
C0160416|T037|PT|865.12|ICD9CM|Injury to spleen with open wound into cavity, capsular tears, without major disruption of parenchyma|Injury to spleen with open wound into cavity, capsular tears, without major disruption of parenchyma
C0160416|T037|AB|865.12|ICD9CM|Spleen capsular tear-opn|Spleen capsular tear-opn
C0160417|T037|PT|865.13|ICD9CM|Injury to spleen with open wound into cavity, laceration extending into parenchyma|Injury to spleen with open wound into cavity, laceration extending into parenchyma
C0160417|T037|AB|865.13|ICD9CM|Spleen parnchym lac-opn|Spleen parnchym lac-opn
C0160418|T037|PT|865.14|ICD9CM|Injury to spleen with open wound into cavity, massive parenchyma disruption|Injury to spleen with open wound into cavity, massive parenchyma disruption
C0160418|T037|AB|865.14|ICD9CM|Spleen disruption-open|Spleen disruption-open
C0160419|T037|PT|865.19|ICD9CM|Other injury to spleen with open wound into cavity|Other injury to spleen with open wound into cavity
C0160419|T037|AB|865.19|ICD9CM|Spleen injury NEC-open|Spleen injury NEC-open
C0160420|T037|HT|866|ICD9CM|Injury to kidney|Injury to kidney
C0160422|T037|HT|866.0|ICD9CM|Injury to kidney without mention of open wound into cavity|Injury to kidney without mention of open wound into cavity
C0160422|T037|PT|866.00|ICD9CM|Injury to kidney without mention of open wound into cavity, unspecified injury|Injury to kidney without mention of open wound into cavity, unspecified injury
C0160422|T037|AB|866.00|ICD9CM|Kidney injury NOS-closed|Kidney injury NOS-closed
C0160423|T037|PT|866.01|ICD9CM|Injury to kidney without mention of open wound into cavity, hematoma without rupture of capsule|Injury to kidney without mention of open wound into cavity, hematoma without rupture of capsule
C0160423|T037|AB|866.01|ICD9CM|Kidney hematoma-closed|Kidney hematoma-closed
C0160424|T037|PT|866.02|ICD9CM|Injury to kidney without mention of open wound into cavity, laceration|Injury to kidney without mention of open wound into cavity, laceration
C0160424|T037|AB|866.02|ICD9CM|Kidney laceration-closed|Kidney laceration-closed
C0273197|T037|PT|866.03|ICD9CM|Injury to kidney without mention of open wound into cavity, complete disruption of kidney parenchyma|Injury to kidney without mention of open wound into cavity, complete disruption of kidney parenchyma
C0273197|T037|AB|866.03|ICD9CM|Kidney disruption-closed|Kidney disruption-closed
C0160427|T037|HT|866.1|ICD9CM|Injury to kidney with open wound into cavity|Injury to kidney with open wound into cavity
C0160427|T037|PT|866.10|ICD9CM|Injury to kidney with open wound into cavity, unspecified injury|Injury to kidney with open wound into cavity, unspecified injury
C0160427|T037|AB|866.10|ICD9CM|Kidney injury NOS-open|Kidney injury NOS-open
C0160428|T037|PT|866.11|ICD9CM|Injury to kidney with open wound into cavity, hematoma without rupture of capsule|Injury to kidney with open wound into cavity, hematoma without rupture of capsule
C0160428|T037|AB|866.11|ICD9CM|Kidney hematoma-open|Kidney hematoma-open
C0160429|T037|PT|866.12|ICD9CM|Injury to kidney with open wound into cavity, laceration|Injury to kidney with open wound into cavity, laceration
C0160429|T037|AB|866.12|ICD9CM|Kidney laceration-open|Kidney laceration-open
C0160430|T037|PT|866.13|ICD9CM|Injury to kidney with open wound into cavity, complete disruption of kidney parenchyma|Injury to kidney with open wound into cavity, complete disruption of kidney parenchyma
C0160430|T037|AB|866.13|ICD9CM|Kidney disruption-open|Kidney disruption-open
C0478263|T037|HT|867|ICD9CM|Injury to pelvic organs|Injury to pelvic organs
C0160432|T037|AB|867.0|ICD9CM|Bladder/urethra inj-clos|Bladder/urethra inj-clos
C0160432|T037|PT|867.0|ICD9CM|Injury to bladder and urethra, without mention of open wound into cavity|Injury to bladder and urethra, without mention of open wound into cavity
C0160433|T037|AB|867.1|ICD9CM|Bladder/urethra inj-open|Bladder/urethra inj-open
C0160433|T037|PT|867.1|ICD9CM|Injury to bladder and urethra, with open wound into cavity|Injury to bladder and urethra, with open wound into cavity
C0160434|T037|PT|867.2|ICD9CM|Injury to ureter, without mention of open wound into cavity|Injury to ureter, without mention of open wound into cavity
C0160434|T037|AB|867.2|ICD9CM|Ureter injury-closed|Ureter injury-closed
C0160435|T037|PT|867.3|ICD9CM|Injury to ureter, with open wound into cavity|Injury to ureter, with open wound into cavity
C0160435|T037|AB|867.3|ICD9CM|Ureter injury-open|Ureter injury-open
C0160436|T037|PT|867.4|ICD9CM|Injury to uterus, without mention of open wound into cavity|Injury to uterus, without mention of open wound into cavity
C0160436|T037|AB|867.4|ICD9CM|Uterus injury-closed|Uterus injury-closed
C0160437|T037|PT|867.5|ICD9CM|Injury to uterus, with open wound into cavity|Injury to uterus, with open wound into cavity
C0160437|T037|AB|867.5|ICD9CM|Uterus injury-open|Uterus injury-open
C0160438|T037|PT|867.6|ICD9CM|Injury to other specified pelvic organs, without mention of open wound into cavity|Injury to other specified pelvic organs, without mention of open wound into cavity
C0160438|T037|AB|867.6|ICD9CM|Pelvic organ inj NEC-cl|Pelvic organ inj NEC-cl
C0160439|T037|PT|867.7|ICD9CM|Injury to other specified pelvic organs, with open wound into cavity|Injury to other specified pelvic organs, with open wound into cavity
C0160439|T037|AB|867.7|ICD9CM|Pelvic organ inj NEC-opn|Pelvic organ inj NEC-opn
C0160440|T037|PT|867.8|ICD9CM|Injury to unspecified pelvic organ, without mention of open wound into cavity|Injury to unspecified pelvic organ, without mention of open wound into cavity
C0160440|T037|AB|867.8|ICD9CM|Pelvic organ inj NOS-cl|Pelvic organ inj NOS-cl
C0160441|T037|PT|867.9|ICD9CM|Injury to unspecified pelvic organ, with open wound into cavity|Injury to unspecified pelvic organ, with open wound into cavity
C0160441|T037|AB|867.9|ICD9CM|Pelvic organ inj NOS-opn|Pelvic organ inj NOS-opn
C3495413|T037|HT|868|ICD9CM|Injury to other intra-abdominal organs|Injury to other intra-abdominal organs
C0160443|T037|HT|868.0|ICD9CM|Injury to other intra-abdominal organs without mention of open wound into cavity|Injury to other intra-abdominal organs without mention of open wound into cavity
C0160444|T037|AB|868.00|ICD9CM|Intra-abdom inj NOS-clos|Intra-abdom inj NOS-clos
C0160445|T037|AB|868.01|ICD9CM|Adrenal gland injury-cl|Adrenal gland injury-cl
C0160445|T037|PT|868.01|ICD9CM|Injury to other intra-abdominal organs without mention of open wound into cavity, adrenal gland|Injury to other intra-abdominal organs without mention of open wound into cavity, adrenal gland
C0160446|T037|AB|868.02|ICD9CM|Biliary tract injury-cl|Biliary tract injury-cl
C0160447|T037|PT|868.03|ICD9CM|Injury to other intra-abdominal organs without mention of open wound into cavity, peritoneum|Injury to other intra-abdominal organs without mention of open wound into cavity, peritoneum
C0160447|T037|AB|868.03|ICD9CM|Peritoneum injury-closed|Peritoneum injury-closed
C0160448|T037|PT|868.04|ICD9CM|Injury to other intra-abdominal organs without mention of open wound into cavity, retroperitoneum|Injury to other intra-abdominal organs without mention of open wound into cavity, retroperitoneum
C0160448|T037|AB|868.04|ICD9CM|Retroperitoneum inj-cl|Retroperitoneum inj-cl
C0160449|T037|PT|868.09|ICD9CM|Injury to other and multiple intra-abdominal organs without mention of open wound into cavity|Injury to other and multiple intra-abdominal organs without mention of open wound into cavity
C0160449|T037|AB|868.09|ICD9CM|Intra-abdom inj NEC-clos|Intra-abdom inj NEC-clos
C0160450|T037|HT|868.1|ICD9CM|Injury to other intra-abdominal organs with open wound into cavity|Injury to other intra-abdominal organs with open wound into cavity
C0160451|T037|AB|868.10|ICD9CM|Intra-abdom inj NOS-open|Intra-abdom inj NOS-open
C0160452|T037|AB|868.11|ICD9CM|Adrenal gland injury-opn|Adrenal gland injury-opn
C0160452|T037|PT|868.11|ICD9CM|Injury to other intra-abdominal organs with open wound into cavity, adrenal gland|Injury to other intra-abdominal organs with open wound into cavity, adrenal gland
C0160453|T037|AB|868.12|ICD9CM|Biliary tract injury-opn|Biliary tract injury-opn
C0160453|T037|PT|868.12|ICD9CM|Injury to other intra-abdominal organs with open wound into cavity, bile duct and gallbladder|Injury to other intra-abdominal organs with open wound into cavity, bile duct and gallbladder
C0160454|T037|PT|868.13|ICD9CM|Injury to other intra-abdominal organs with open wound into cavity, peritoneum|Injury to other intra-abdominal organs with open wound into cavity, peritoneum
C0160454|T037|AB|868.13|ICD9CM|Peritoneum injury-open|Peritoneum injury-open
C0160455|T037|PT|868.14|ICD9CM|Injury to other intra-abdominal organs with open wound into cavity, retroperitoneum|Injury to other intra-abdominal organs with open wound into cavity, retroperitoneum
C0160455|T037|AB|868.14|ICD9CM|Retroperitoneum inj-open|Retroperitoneum inj-open
C0160456|T037|PT|868.19|ICD9CM|Injury to other and multiple intra-abdominal organs, with open wound into cavity|Injury to other and multiple intra-abdominal organs, with open wound into cavity
C0160456|T037|AB|868.19|ICD9CM|Intra-abdom inj NEC-open|Intra-abdom inj NEC-open
C0160457|T037|HT|869|ICD9CM|Internal injury to unspecified or ill-defined organs|Internal injury to unspecified or ill-defined organs
C0021779|T037|AB|869.0|ICD9CM|Internal inj NOS-closed|Internal inj NOS-closed
C0021779|T037|PT|869.0|ICD9CM|Internal injury to unspecified or ill-defined organs without mention of open wound into cavity|Internal injury to unspecified or ill-defined organs without mention of open wound into cavity
C0160458|T037|AB|869.1|ICD9CM|Internal injury NOS-open|Internal injury NOS-open
C0160458|T037|PT|869.1|ICD9CM|Internal injury to unspecified or ill-defined organs with open wound into cavity|Internal injury to unspecified or ill-defined organs with open wound into cavity
C0160459|T037|HT|870|ICD9CM|Open wound of ocular adnexa|Open wound of ocular adnexa
C0178321|T037|HT|870-879.99|ICD9CM|OPEN WOUND OF HEAD, NECK, AND TRUNK|OPEN WOUND OF HEAD, NECK, AND TRUNK
C0332798|T037|HT|870-897.99|ICD9CM|OPEN WOUNDS|OPEN WOUNDS
C0160460|T037|AB|870.0|ICD9CM|Lac eyelid skn/perioculr|Lac eyelid skn/perioculr
C0160460|T037|PT|870.0|ICD9CM|Laceration of skin of eyelid and periocular area|Laceration of skin of eyelid and periocular area
C0433980|T037|AB|870.1|ICD9CM|Full-thicknes lac eyelid|Full-thicknes lac eyelid
C0433980|T037|PT|870.1|ICD9CM|Laceration of eyelid, full-thickness, not involving lacrimal passages|Laceration of eyelid, full-thickness, not involving lacrimal passages
C0433981|T037|AB|870.2|ICD9CM|Lac eyelid inv lacrm pas|Lac eyelid inv lacrm pas
C0433981|T037|PT|870.2|ICD9CM|Laceration of eyelid involving lacrimal passages|Laceration of eyelid involving lacrimal passages
C0273244|T037|AB|870.3|ICD9CM|Penetr wnd orbit w/o FB|Penetr wnd orbit w/o FB
C0273244|T037|PT|870.3|ICD9CM|Penetrating wound of orbit, without mention of foreign body|Penetrating wound of orbit, without mention of foreign body
C0160464|T037|AB|870.4|ICD9CM|Penetrat wnd orbit w FB|Penetrat wnd orbit w FB
C0160464|T037|PT|870.4|ICD9CM|Penetrating wound of orbit with foreign body|Penetrating wound of orbit with foreign body
C0160465|T037|AB|870.8|ICD9CM|Opn wnd ocular adnex NEC|Opn wnd ocular adnex NEC
C0160465|T037|PT|870.8|ICD9CM|Other specified open wounds of ocular adnexa|Other specified open wounds of ocular adnexa
C0160466|T037|AB|870.9|ICD9CM|Opn wnd ocular adnex NOS|Opn wnd ocular adnex NOS
C0160466|T037|PT|870.9|ICD9CM|Unspecified open wound of ocular adnexa|Unspecified open wound of ocular adnexa
C0160474|T037|HT|871|ICD9CM|Open wound of eyeball|Open wound of eyeball
C0433976|T037|AB|871.0|ICD9CM|Ocular lac w/o prolapse|Ocular lac w/o prolapse
C0433976|T037|PT|871.0|ICD9CM|Ocular laceration without prolapse of intraocular tissue|Ocular laceration without prolapse of intraocular tissue
C0160468|T037|AB|871.1|ICD9CM|Ocular lacera w prolapse|Ocular lacera w prolapse
C0160468|T037|PT|871.1|ICD9CM|Ocular laceration with prolapse or exposure of intraocular tissue|Ocular laceration with prolapse or exposure of intraocular tissue
C0160469|T037|AB|871.2|ICD9CM|Rupture eye w tissu loss|Rupture eye w tissu loss
C0160469|T037|PT|871.2|ICD9CM|Rupture of eye with partial loss of intraocular tissue|Rupture of eye with partial loss of intraocular tissue
C0004445|T037|AB|871.3|ICD9CM|Avulsion of eye|Avulsion of eye
C0004445|T037|PT|871.3|ICD9CM|Avulsion of eye|Avulsion of eye
C0160470|T037|AB|871.4|ICD9CM|Laceration of eye NOS|Laceration of eye NOS
C0160470|T037|PT|871.4|ICD9CM|Unspecified laceration of eye|Unspecified laceration of eye
C0160471|T037|AB|871.5|ICD9CM|Penetrat magnet FB eye|Penetrat magnet FB eye
C0160471|T037|PT|871.5|ICD9CM|Penetration of eyeball with magnetic foreign body|Penetration of eyeball with magnetic foreign body
C0160472|T037|AB|871.6|ICD9CM|Penetrat FB NEC eye|Penetrat FB NEC eye
C0160472|T037|PT|871.6|ICD9CM|Penetration of eyeball with (nonmagnetic) foreign body|Penetration of eyeball with (nonmagnetic) foreign body
C0015409|T037|AB|871.7|ICD9CM|Ocular penetration NOS|Ocular penetration NOS
C0015409|T037|PT|871.7|ICD9CM|Unspecified ocular penetration|Unspecified ocular penetration
C0160474|T037|AB|871.9|ICD9CM|Opn wound of eyeball NOS|Opn wound of eyeball NOS
C0160474|T037|PT|871.9|ICD9CM|Unspecified open wound of eyeball|Unspecified open wound of eyeball
C0160475|T037|HT|872|ICD9CM|Open wound of ear|Open wound of ear
C0160476|T037|HT|872.0|ICD9CM|Open wound of external ear, without mention of complication|Open wound of external ear, without mention of complication
C0375641|T037|PT|872.00|ICD9CM|Open wound of external ear, unspecified site, without mention of complication|Open wound of external ear, unspecified site, without mention of complication
C0375641|T037|AB|872.00|ICD9CM|Opn wound extern ear NOS|Opn wound extern ear NOS
C0273248|T037|AB|872.01|ICD9CM|Open wound of auricle|Open wound of auricle
C0273248|T037|PT|872.01|ICD9CM|Open wound of auricle, ear, without mention of complication|Open wound of auricle, ear, without mention of complication
C0375643|T037|PT|872.02|ICD9CM|Open wound of auditory canal, without mention of complication|Open wound of auditory canal, without mention of complication
C0375643|T037|AB|872.02|ICD9CM|Opn wound auditory canal|Opn wound auditory canal
C0273251|T037|HT|872.1|ICD9CM|Open wound of external ear, complicated|Open wound of external ear, complicated
C0160481|T037|PT|872.10|ICD9CM|Open wound of external ear, unspecified site, complicated|Open wound of external ear, unspecified site, complicated
C0160481|T037|AB|872.10|ICD9CM|Opn wnd ex ear NOS-compl|Opn wnd ex ear NOS-compl
C0160482|T037|AB|872.11|ICD9CM|Open wound auricle-compl|Open wound auricle-compl
C0160482|T037|PT|872.11|ICD9CM|Open wound of auricle, ear, complicated|Open wound of auricle, ear, complicated
C0160483|T037|AB|872.12|ICD9CM|Open wnd aud canal-compl|Open wnd aud canal-compl
C0160483|T037|PT|872.12|ICD9CM|Open wound of auditory canal, complicated|Open wound of auditory canal, complicated
C0160484|T037|HT|872.6|ICD9CM|Open wound of other specified parts of ear, without mention of complication|Open wound of other specified parts of ear, without mention of complication
C0273253|T037|AB|872.61|ICD9CM|Open wound of ear drum|Open wound of ear drum
C0273253|T037|PT|872.61|ICD9CM|Open wound of ear drum, without mention of complication|Open wound of ear drum, without mention of complication
C0273254|T037|AB|872.62|ICD9CM|Open wound of ossicles|Open wound of ossicles
C0273254|T037|PT|872.62|ICD9CM|Open wound of ossicles, without mention of complication|Open wound of ossicles, without mention of complication
C0375646|T037|AB|872.63|ICD9CM|Open wnd eustachian tube|Open wnd eustachian tube
C0375646|T037|PT|872.63|ICD9CM|Open wound of eustachian tube, without mention of complication|Open wound of eustachian tube, without mention of complication
C0273256|T037|AB|872.64|ICD9CM|Open wound of cochlea|Open wound of cochlea
C0273256|T037|PT|872.64|ICD9CM|Open wound of cochlea, without mention of complication|Open wound of cochlea, without mention of complication
C0490055|T037|AB|872.69|ICD9CM|Open wound of ear NEC|Open wound of ear NEC
C0490055|T037|PT|872.69|ICD9CM|Open wound of other and multiple sites of ear, without mention of complication|Open wound of other and multiple sites of ear, without mention of complication
C0160489|T037|HT|872.7|ICD9CM|Open wound of other specified parts of ear, complicated|Open wound of other specified parts of ear, complicated
C0160490|T037|AB|872.71|ICD9CM|Open wnd ear drum-compl|Open wnd ear drum-compl
C0160490|T037|PT|872.71|ICD9CM|Open wound of ear drum, complicated|Open wound of ear drum, complicated
C0160491|T037|AB|872.72|ICD9CM|Open wnd ossicles-compl|Open wnd ossicles-compl
C0160491|T037|PT|872.72|ICD9CM|Open wound of ossicles, complicated|Open wound of ossicles, complicated
C0160492|T037|PT|872.73|ICD9CM|Open wound of eustachian tube, complicated|Open wound of eustachian tube, complicated
C0160492|T037|AB|872.73|ICD9CM|Opn wnd eustach tb-compl|Opn wnd eustach tb-compl
C0160493|T037|AB|872.74|ICD9CM|Open wound cochlea-compl|Open wound cochlea-compl
C0160493|T037|PT|872.74|ICD9CM|Open wound of cochlea, complicated|Open wound of cochlea, complicated
C0490056|T037|AB|872.79|ICD9CM|Open wound ear NEC-compl|Open wound ear NEC-compl
C0490056|T037|PT|872.79|ICD9CM|Open wound of other and multiple sites of ear, complicated|Open wound of other and multiple sites of ear, complicated
C0160475|T037|AB|872.8|ICD9CM|Open wound of ear NOS|Open wound of ear NOS
C0160475|T037|PT|872.8|ICD9CM|Open wound of ear, part unspecified, without mention of complication|Open wound of ear, part unspecified, without mention of complication
C0273250|T037|AB|872.9|ICD9CM|Open wound ear NOS-compl|Open wound ear NOS-compl
C0273250|T037|PT|872.9|ICD9CM|Open wound of ear, part unspecified, complicated|Open wound of ear, part unspecified, complicated
C0160496|T037|HT|873|ICD9CM|Other open wound of head|Other open wound of head
C0273259|T037|AB|873.0|ICD9CM|Open wound of scalp|Open wound of scalp
C0273259|T037|PT|873.0|ICD9CM|Open wound of scalp, without mention of complication|Open wound of scalp, without mention of complication
C0160498|T037|PT|873.1|ICD9CM|Open wound of scalp, complicated|Open wound of scalp, complicated
C0160498|T037|AB|873.1|ICD9CM|Open wound scalp-compl|Open wound scalp-compl
C0273260|T037|HT|873.2|ICD9CM|Open wound of nose, without mention of complication|Open wound of nose, without mention of complication
C0273260|T037|AB|873.20|ICD9CM|Open wound of nose NOS|Open wound of nose NOS
C0273260|T037|PT|873.20|ICD9CM|Open wound of nose, unspecified site, without mention of complication|Open wound of nose, unspecified site, without mention of complication
C0375650|T037|AB|873.21|ICD9CM|Open wound nasal septum|Open wound nasal septum
C0375650|T037|PT|873.21|ICD9CM|Open wound of nasal septum, without mention of complication|Open wound of nasal septum, without mention of complication
C0160502|T037|AB|873.22|ICD9CM|Open wound nasal cavity|Open wound nasal cavity
C0160502|T037|PT|873.22|ICD9CM|Open wound of nasal cavity, without mention of complication|Open wound of nasal cavity, without mention of complication
C0160503|T037|AB|873.23|ICD9CM|Open wound nasal sinus|Open wound nasal sinus
C0160503|T037|PT|873.23|ICD9CM|Open wound of nasal sinus, without mention of complication|Open wound of nasal sinus, without mention of complication
C0375653|T037|AB|873.29|ICD9CM|Mult open wound nose|Mult open wound nose
C0375653|T037|PT|873.29|ICD9CM|Open wound of multiple sites of nose, without mention of complication|Open wound of multiple sites of nose, without mention of complication
C0160505|T037|HT|873.3|ICD9CM|Open wound of nose, complicated|Open wound of nose, complicated
C0160505|T037|AB|873.30|ICD9CM|Open wnd nose NOS-compl|Open wnd nose NOS-compl
C0160505|T037|PT|873.30|ICD9CM|Open wound of nose, unspecified site, complicated|Open wound of nose, unspecified site, complicated
C0160507|T037|PT|873.31|ICD9CM|Open wound of nasal septum, complicated|Open wound of nasal septum, complicated
C0160507|T037|AB|873.31|ICD9CM|Opn wnd nas septum-compl|Opn wnd nas septum-compl
C0160508|T037|AB|873.32|ICD9CM|Open wnd nasal cav-compl|Open wnd nasal cav-compl
C0160508|T037|PT|873.32|ICD9CM|Open wound of nasal cavity, complicated|Open wound of nasal cavity, complicated
C0160509|T037|AB|873.33|ICD9CM|Open wnd nas sinus-compl|Open wnd nas sinus-compl
C0160509|T037|PT|873.33|ICD9CM|Open wound of nasal sinus, complicated|Open wound of nasal sinus, complicated
C0273237|T037|AB|873.39|ICD9CM|Mult open wnd nose-compl|Mult open wnd nose-compl
C0273237|T037|PT|873.39|ICD9CM|Open wound of multiple sites of nose, complicated|Open wound of multiple sites of nose, complicated
C0160511|T037|HT|873.4|ICD9CM|Open wound of face, without mention of complication|Open wound of face, without mention of complication
C0375654|T037|AB|873.40|ICD9CM|Open wound of face NOS|Open wound of face NOS
C0375654|T037|PT|873.40|ICD9CM|Open wound of face, unspecified site, without mention of complication|Open wound of face, unspecified site, without mention of complication
C0273267|T037|AB|873.41|ICD9CM|Open wound of cheek|Open wound of cheek
C0273267|T037|PT|873.41|ICD9CM|Open wound of cheek, without mention of complication|Open wound of cheek, without mention of complication
C0273268|T037|AB|873.42|ICD9CM|Open wound of forehead|Open wound of forehead
C0273268|T037|PT|873.42|ICD9CM|Open wound of forehead, without mention of complication|Open wound of forehead, without mention of complication
C0273270|T037|AB|873.43|ICD9CM|Open wound of lip|Open wound of lip
C0273270|T037|PT|873.43|ICD9CM|Open wound of lip, without mention of complication|Open wound of lip, without mention of complication
C0273271|T037|AB|873.44|ICD9CM|Open wound of jaw|Open wound of jaw
C0273271|T037|PT|873.44|ICD9CM|Open wound of jaw, without mention of complication|Open wound of jaw, without mention of complication
C0490057|T037|AB|873.49|ICD9CM|Open wound of face NEC|Open wound of face NEC
C0490057|T037|PT|873.49|ICD9CM|Open wound of other and multiple sites of face, without mention of complication|Open wound of other and multiple sites of face, without mention of complication
C0160517|T037|HT|873.5|ICD9CM|Open wound of face, complicated|Open wound of face, complicated
C0160517|T037|AB|873.50|ICD9CM|Open wnd face NOS-compl|Open wnd face NOS-compl
C0160517|T037|PT|873.50|ICD9CM|Open wound of face, unspecified site, complicated|Open wound of face, unspecified site, complicated
C0160519|T037|AB|873.51|ICD9CM|Open wound cheek-compl|Open wound cheek-compl
C0160519|T037|PT|873.51|ICD9CM|Open wound of cheek, complicated|Open wound of cheek, complicated
C0160520|T037|AB|873.52|ICD9CM|Open wnd forehead-compl|Open wnd forehead-compl
C0160520|T037|PT|873.52|ICD9CM|Open wound of forehead, complicated|Open wound of forehead, complicated
C0160521|T037|AB|873.53|ICD9CM|Open wound lip-complicat|Open wound lip-complicat
C0160521|T037|PT|873.53|ICD9CM|Open wound of lip, complicated|Open wound of lip, complicated
C0160522|T037|AB|873.54|ICD9CM|Open wound jaw-complicat|Open wound jaw-complicat
C0160522|T037|PT|873.54|ICD9CM|Open wound of jaw, complicated|Open wound of jaw, complicated
C0490058|T037|AB|873.59|ICD9CM|Open wnd face NEC-compl|Open wnd face NEC-compl
C0490058|T037|PT|873.59|ICD9CM|Open wound of other and multiple sites of face, complicated|Open wound of other and multiple sites of face, complicated
C0160523|T037|HT|873.6|ICD9CM|Open wound of internal structures of mouth, without mention of complication|Open wound of internal structures of mouth, without mention of complication
C0375659|T037|AB|873.60|ICD9CM|Open wound of mouth NOS|Open wound of mouth NOS
C0375659|T037|PT|873.60|ICD9CM|Open wound of mouth, unspecified site, without mention of complication|Open wound of mouth, unspecified site, without mention of complication
C0273276|T037|AB|873.61|ICD9CM|Open wound buccal mucosa|Open wound buccal mucosa
C0273276|T037|PT|873.61|ICD9CM|Open wound of buccal mucosa, without mention of complication|Open wound of buccal mucosa, without mention of complication
C0273277|T037|AB|873.62|ICD9CM|Open wound of gum|Open wound of gum
C0273277|T037|PT|873.62|ICD9CM|Open wound of gum (alveolar process), without mention of complication|Open wound of gum (alveolar process), without mention of complication
C0375662|T037|AB|873.63|ICD9CM|Broken tooth-uncomplic|Broken tooth-uncomplic
C0375662|T037|PT|873.63|ICD9CM|Open wound of tooth (broken) (fractured) (due to trauma), without mention of complication|Open wound of tooth (broken) (fractured) (due to trauma), without mention of complication
C0375663|T037|PT|873.64|ICD9CM|Open wound of tongue and floor of mouth, without mention of complication|Open wound of tongue and floor of mouth, without mention of complication
C0375663|T037|AB|873.64|ICD9CM|Opn wnd tongue/mouth flr|Opn wnd tongue/mouth flr
C0273282|T037|AB|873.65|ICD9CM|Open wound of palate|Open wound of palate
C0273282|T037|PT|873.65|ICD9CM|Open wound of palate, without mention of complication|Open wound of palate, without mention of complication
C0490059|T037|AB|873.69|ICD9CM|Open wound mouth NEC|Open wound mouth NEC
C0490059|T037|PT|873.69|ICD9CM|Open wound of other and multiple sites of mouth, without mention of complication|Open wound of other and multiple sites of mouth, without mention of complication
C0160529|T037|HT|873.7|ICD9CM|Open wound of internal structure of mouth, complicated|Open wound of internal structure of mouth, complicated
C0273284|T037|AB|873.70|ICD9CM|Open wnd mouth NOS-compl|Open wnd mouth NOS-compl
C0273284|T037|PT|873.70|ICD9CM|Open wound of mouth, unspecified site, complicated|Open wound of mouth, unspecified site, complicated
C0160531|T037|PT|873.71|ICD9CM|Open wound of buccal mucosa, complicated|Open wound of buccal mucosa, complicated
C0160531|T037|AB|873.71|ICD9CM|Opn wnd buc mucosa-compl|Opn wnd buc mucosa-compl
C0273286|T037|AB|873.72|ICD9CM|Open wound gum-compl|Open wound gum-compl
C0273286|T037|PT|873.72|ICD9CM|Open wound of gum (alveolar process), complicated|Open wound of gum (alveolar process), complicated
C0160533|T037|AB|873.73|ICD9CM|Broken tooth-complicated|Broken tooth-complicated
C0160533|T037|PT|873.73|ICD9CM|Open wound of tooth (broken) (fractured) (due to trauma), complicated|Open wound of tooth (broken) (fractured) (due to trauma), complicated
C0160534|T037|PT|873.74|ICD9CM|Open wound of tongue and floor of mouth, complicated|Open wound of tongue and floor of mouth, complicated
C0160534|T037|AB|873.74|ICD9CM|Open wound tongue-compl|Open wound tongue-compl
C0160535|T037|PT|873.75|ICD9CM|Open wound of palate, complicated|Open wound of palate, complicated
C0160535|T037|AB|873.75|ICD9CM|Open wound palate-compl|Open wound palate-compl
C0490060|T037|AB|873.79|ICD9CM|Open wnd mouth NOS-compl|Open wnd mouth NOS-compl
C0490060|T037|PT|873.79|ICD9CM|Open wound of other and multiple sites of mouth, complicated|Open wound of other and multiple sites of mouth, complicated
C0160536|T037|AB|873.8|ICD9CM|Open wound of head NEC|Open wound of head NEC
C0160536|T037|PT|873.8|ICD9CM|Other and unspecified open wound of head without mention of complication|Other and unspecified open wound of head without mention of complication
C0160537|T037|AB|873.9|ICD9CM|Open wnd head NEC-compl|Open wnd head NEC-compl
C0160537|T037|PT|873.9|ICD9CM|Other and unspecified open wound of head, complicated|Other and unspecified open wound of head, complicated
C0160538|T037|HT|874|ICD9CM|Open wound of neck|Open wound of neck
C0160539|T037|HT|874.0|ICD9CM|Open wound of larynx and trachea, without mention of complication|Open wound of larynx and trachea, without mention of complication
C0160539|T037|PT|874.00|ICD9CM|Open wound of larynx with trachea, without mention of complication|Open wound of larynx with trachea, without mention of complication
C0160539|T037|AB|874.00|ICD9CM|Opn wnd larynx w trachea|Opn wnd larynx w trachea
C0273300|T037|AB|874.01|ICD9CM|Open wound of larynx|Open wound of larynx
C0273300|T037|PT|874.01|ICD9CM|Open wound of larynx, without mention of complication|Open wound of larynx, without mention of complication
C0273301|T037|AB|874.02|ICD9CM|Open wound of trachea|Open wound of trachea
C0273301|T037|PT|874.02|ICD9CM|Open wound of trachea, without mention of complication|Open wound of trachea, without mention of complication
C0160543|T037|HT|874.1|ICD9CM|Open wound of larynx and trachea, complicated|Open wound of larynx and trachea, complicated
C0160543|T037|PT|874.10|ICD9CM|Open wound of larynx with trachea, complicated|Open wound of larynx with trachea, complicated
C0160543|T037|AB|874.10|ICD9CM|Opn wnd lary w trac-comp|Opn wnd lary w trac-comp
C0160544|T037|AB|874.11|ICD9CM|Open wound larynx-compl|Open wound larynx-compl
C0160544|T037|PT|874.11|ICD9CM|Open wound of larynx, complicated|Open wound of larynx, complicated
C0160545|T037|PT|874.12|ICD9CM|Open wound of trachea, complicated|Open wound of trachea, complicated
C0160545|T037|AB|874.12|ICD9CM|Open wound trachea-compl|Open wound trachea-compl
C0273302|T037|PT|874.2|ICD9CM|Open wound of thyroid gland, without mention of complication|Open wound of thyroid gland, without mention of complication
C0273302|T037|AB|874.2|ICD9CM|Open wound thyroid gland|Open wound thyroid gland
C0160547|T037|PT|874.3|ICD9CM|Open wound of thyroid gland, complicated|Open wound of thyroid gland, complicated
C0160547|T037|AB|874.3|ICD9CM|Open wound thyroid-compl|Open wound thyroid-compl
C0273292|T037|AB|874.4|ICD9CM|Open wound of pharynx|Open wound of pharynx
C0273292|T037|PT|874.4|ICD9CM|Open wound of pharynx, without mention of complication|Open wound of pharynx, without mention of complication
C0160549|T037|PT|874.5|ICD9CM|Open wound of pharynx, complicated|Open wound of pharynx, complicated
C0160549|T037|AB|874.5|ICD9CM|Open wound pharynx-compl|Open wound pharynx-compl
C0160550|T037|AB|874.8|ICD9CM|Open wound of neck NEC|Open wound of neck NEC
C0160550|T037|PT|874.8|ICD9CM|Open wound of other and unspecified parts of neck, without mention of complication|Open wound of other and unspecified parts of neck, without mention of complication
C0160551|T037|PT|874.9|ICD9CM|Open wound of other and unspecified parts of neck, complicated|Open wound of other and unspecified parts of neck, complicated
C0160551|T037|AB|874.9|ICD9CM|Opn wound neck NEC-compl|Opn wound neck NEC-compl
C0160552|T037|HT|875|ICD9CM|Open wound of chest (wall)|Open wound of chest (wall)
C0273313|T037|AB|875.0|ICD9CM|Open wound of chest|Open wound of chest
C0273313|T037|PT|875.0|ICD9CM|Open wound of chest (wall), without mention of complication|Open wound of chest (wall), without mention of complication
C0273314|T037|AB|875.1|ICD9CM|Open wound chest-compl|Open wound chest-compl
C0273314|T037|PT|875.1|ICD9CM|Open wound of chest (wall), complicated|Open wound of chest (wall), complicated
C0160555|T037|HT|876|ICD9CM|Open wound of back|Open wound of back
C0273315|T037|AB|876.0|ICD9CM|Open wound of back|Open wound of back
C0273315|T037|PT|876.0|ICD9CM|Open wound of back, without mention of complication|Open wound of back, without mention of complication
C0160557|T037|AB|876.1|ICD9CM|Open wound back-compl|Open wound back-compl
C0160557|T037|PT|876.1|ICD9CM|Open wound of back, complicated|Open wound of back, complicated
C0160558|T037|HT|877|ICD9CM|Open wound of buttock|Open wound of buttock
C0273318|T037|AB|877.0|ICD9CM|Open wound of buttock|Open wound of buttock
C0273318|T037|PT|877.0|ICD9CM|Open wound of buttock, without mention of complication|Open wound of buttock, without mention of complication
C0160560|T037|AB|877.1|ICD9CM|Open wound buttock-compl|Open wound buttock-compl
C0160560|T037|PT|877.1|ICD9CM|Open wound of buttock, complicated|Open wound of buttock, complicated
C0160561|T037|HT|878|ICD9CM|Open wound of genital organs (external), including traumatic amputation|Open wound of genital organs (external), including traumatic amputation
C0160562|T037|AB|878.0|ICD9CM|Open wound of penis|Open wound of penis
C0160562|T037|PT|878.0|ICD9CM|Open wound of penis, without mention of complication|Open wound of penis, without mention of complication
C0160563|T037|PT|878.1|ICD9CM|Open wound of penis, complicated|Open wound of penis, complicated
C0160563|T037|AB|878.1|ICD9CM|Open wound penis-compl|Open wound penis-compl
C0434143|T037|PT|878.2|ICD9CM|Open wound of scrotum and testes, without mention of complication|Open wound of scrotum and testes, without mention of complication
C0434143|T037|AB|878.2|ICD9CM|Opn wound scrotum/testes|Opn wound scrotum/testes
C0160565|T037|PT|878.3|ICD9CM|Open wound of scrotum and testes, complicated|Open wound of scrotum and testes, complicated
C0160565|T037|AB|878.3|ICD9CM|Opn wnd scrot/test-compl|Opn wnd scrot/test-compl
C0273329|T037|AB|878.4|ICD9CM|Open wound of vulva|Open wound of vulva
C0273329|T037|PT|878.4|ICD9CM|Open wound of vulva, without mention of complication|Open wound of vulva, without mention of complication
C0160567|T037|PT|878.5|ICD9CM|Open wound of vulva, complicated|Open wound of vulva, complicated
C0160567|T037|AB|878.5|ICD9CM|Open wound vulva-compl|Open wound vulva-compl
C0273330|T037|AB|878.6|ICD9CM|Open wound of vagina|Open wound of vagina
C0273330|T037|PT|878.6|ICD9CM|Open wound of vagina, without mention of complication|Open wound of vagina, without mention of complication
C0160569|T037|PT|878.7|ICD9CM|Open wound of vagina, complicated|Open wound of vagina, complicated
C0160569|T037|AB|878.7|ICD9CM|Open wound vagina-compl|Open wound vagina-compl
C0160570|T037|AB|878.8|ICD9CM|Open wound genital NEC|Open wound genital NEC
C0160571|T037|PT|878.9|ICD9CM|Open wound of other and unspecified parts of genital organs (external), complicated|Open wound of other and unspecified parts of genital organs (external), complicated
C0160571|T037|AB|878.9|ICD9CM|Opn wnd genital NEC-comp|Opn wnd genital NEC-comp
C0160572|T037|HT|879|ICD9CM|Open wound of other and unspecified sites, except limbs|Open wound of other and unspecified sites, except limbs
C0347564|T037|AB|879.0|ICD9CM|Open wound of breast|Open wound of breast
C0347564|T037|PT|879.0|ICD9CM|Open wound of breast, without mention of complication|Open wound of breast, without mention of complication
C0160574|T037|AB|879.1|ICD9CM|Open wound breast-compl|Open wound breast-compl
C0160574|T037|PT|879.1|ICD9CM|Open wound of breast, complicated|Open wound of breast, complicated
C0160575|T037|PT|879.2|ICD9CM|Open wound of abdominal wall, anterior, without mention of complication|Open wound of abdominal wall, anterior, without mention of complication
C0160575|T037|AB|879.2|ICD9CM|Opn wnd anterior abdomen|Opn wnd anterior abdomen
C0160576|T037|PT|879.3|ICD9CM|Open wound of abdominal wall, anterior, complicated|Open wound of abdominal wall, anterior, complicated
C0160576|T037|AB|879.3|ICD9CM|Opn wnd ant abdomen-comp|Opn wnd ant abdomen-comp
C0160577|T037|PT|879.4|ICD9CM|Open wound of abdominal wall, lateral, without mention of complication|Open wound of abdominal wall, lateral, without mention of complication
C0160577|T037|AB|879.4|ICD9CM|Opn wnd lateral abdomen|Opn wnd lateral abdomen
C0160578|T037|PT|879.5|ICD9CM|Open wound of abdominal wall, lateral, complicated|Open wound of abdominal wall, lateral, complicated
C0160578|T037|AB|879.5|ICD9CM|Opn wnd lat abdomen-comp|Opn wnd lat abdomen-comp
C0160579|T037|PT|879.6|ICD9CM|Open wound of other and unspecified parts of trunk, without mention of complication|Open wound of other and unspecified parts of trunk, without mention of complication
C0160579|T037|AB|879.6|ICD9CM|Open wound of trunk NEC|Open wound of trunk NEC
C0160580|T037|AB|879.7|ICD9CM|Open wnd trunk NEC-compl|Open wnd trunk NEC-compl
C0160580|T037|PT|879.7|ICD9CM|Open wound of other and unspecified parts of trunk, complicated|Open wound of other and unspecified parts of trunk, complicated
C0273236|T037|AB|879.8|ICD9CM|Open wound site NOS|Open wound site NOS
C0273236|T037|PT|879.8|ICD9CM|Open wound(s) (multiple) of unspecified site(s), without mention of complication|Open wound(s) (multiple) of unspecified site(s), without mention of complication
C0273237|T037|PT|879.9|ICD9CM|Open wound(s) (multiple) of unspecified site(s), complicated|Open wound(s) (multiple) of unspecified site(s), complicated
C0273237|T037|AB|879.9|ICD9CM|Opn wound site NOS-compl|Opn wound site NOS-compl
C0432959|T037|HT|880|ICD9CM|Open wound of shoulder and upper arm|Open wound of shoulder and upper arm
C0178322|T037|HT|880-887.99|ICD9CM|OPEN WOUND OF UPPER LIMB|OPEN WOUND OF UPPER LIMB
C0160584|T037|HT|880.0|ICD9CM|Open wound of shoulder and upper arm, without mention of complication|Open wound of shoulder and upper arm, without mention of complication
C0273354|T037|AB|880.00|ICD9CM|Open wound of shoulder|Open wound of shoulder
C0273354|T037|PT|880.00|ICD9CM|Open wound of shoulder region, without mention of complication|Open wound of shoulder region, without mention of complication
C0160586|T037|AB|880.01|ICD9CM|Open wound of scapula|Open wound of scapula
C0160586|T037|PT|880.01|ICD9CM|Open wound of scapular region, without mention of complication|Open wound of scapular region, without mention of complication
C0160587|T037|AB|880.02|ICD9CM|Open wound of axilla|Open wound of axilla
C0160587|T037|PT|880.02|ICD9CM|Open wound of axillary region, without mention of complication|Open wound of axillary region, without mention of complication
C0160588|T037|AB|880.03|ICD9CM|Open wound of upper arm|Open wound of upper arm
C0160588|T037|PT|880.03|ICD9CM|Open wound of upper arm, without mention of complication|Open wound of upper arm, without mention of complication
C0495858|T037|AB|880.09|ICD9CM|Mult open wound shoulder|Mult open wound shoulder
C0495858|T037|PT|880.09|ICD9CM|Open wound of multiple sites of shoulder and upper arm, without mention of complication|Open wound of multiple sites of shoulder and upper arm, without mention of complication
C0160590|T037|HT|880.1|ICD9CM|Open wound of shoulder and upper arm, complicated|Open wound of shoulder and upper arm, complicated
C0160591|T037|AB|880.10|ICD9CM|Open wnd shoulder-compl|Open wnd shoulder-compl
C0160591|T037|PT|880.10|ICD9CM|Open wound of shoulder region, complicated|Open wound of shoulder region, complicated
C0160592|T037|PT|880.11|ICD9CM|Open wound of scapular region, complicated|Open wound of scapular region, complicated
C0160592|T037|AB|880.11|ICD9CM|Open wound scapula-compl|Open wound scapula-compl
C0160593|T037|AB|880.12|ICD9CM|Open wound axilla-compl|Open wound axilla-compl
C0160593|T037|PT|880.12|ICD9CM|Open wound of axillary region, complicated|Open wound of axillary region, complicated
C0160594|T037|AB|880.13|ICD9CM|Open wnd upper arm-compl|Open wnd upper arm-compl
C0160594|T037|PT|880.13|ICD9CM|Open wound of upper arm, complicated|Open wound of upper arm, complicated
C0160595|T037|AB|880.19|ICD9CM|Mult opn wnd should-comp|Mult opn wnd should-comp
C0160595|T037|PT|880.19|ICD9CM|Open wound of multiple sites of shoulder and upper arm, complicated|Open wound of multiple sites of shoulder and upper arm, complicated
C0160596|T037|HT|880.2|ICD9CM|Open wound of shoulder and upper arm, with tendon involvement|Open wound of shoulder and upper arm, with tendon involvement
C0160597|T037|PT|880.20|ICD9CM|Open wound of shoulder region, with tendon involvement|Open wound of shoulder region, with tendon involvement
C0160597|T037|AB|880.20|ICD9CM|Opn wnd shouldr w tendon|Opn wnd shouldr w tendon
C0160598|T037|PT|880.21|ICD9CM|Open wound of scapular region, with tendon involvement|Open wound of scapular region, with tendon involvement
C0160598|T037|AB|880.21|ICD9CM|Opn wnd scapula w tendon|Opn wnd scapula w tendon
C0160599|T037|AB|880.22|ICD9CM|Open wnd axilla w tendon|Open wnd axilla w tendon
C0160599|T037|PT|880.22|ICD9CM|Open wound of axillary region, with tendon involvement|Open wound of axillary region, with tendon involvement
C0160600|T037|AB|880.23|ICD9CM|Open wnd up arm w tendon|Open wnd up arm w tendon
C0160600|T037|PT|880.23|ICD9CM|Open wound of upper arm, with tendon involvement|Open wound of upper arm, with tendon involvement
C0160601|T037|AB|880.29|ICD9CM|Mlt opn wnd shldr w tend|Mlt opn wnd shldr w tend
C0160601|T037|PT|880.29|ICD9CM|Open wound of multiple sites of shoulder and upper arm, with tendon involvement|Open wound of multiple sites of shoulder and upper arm, with tendon involvement
C0160602|T037|HT|881|ICD9CM|Open wound of elbow, forearm, and wrist|Open wound of elbow, forearm, and wrist
C0160603|T037|HT|881.0|ICD9CM|Open wound of elbow, forearm, and wrist, without mention of complication|Open wound of elbow, forearm, and wrist, without mention of complication
C0160604|T037|AB|881.00|ICD9CM|Open wound of forearm|Open wound of forearm
C0160604|T037|PT|881.00|ICD9CM|Open wound of forearm, without mention of complication|Open wound of forearm, without mention of complication
C0160605|T037|AB|881.01|ICD9CM|Open wound of elbow|Open wound of elbow
C0160605|T037|PT|881.01|ICD9CM|Open wound of elbow, without mention of complication|Open wound of elbow, without mention of complication
C0160606|T037|AB|881.02|ICD9CM|Open wound of wrist|Open wound of wrist
C0160606|T037|PT|881.02|ICD9CM|Open wound of wrist, without mention of complication|Open wound of wrist, without mention of complication
C0160607|T037|HT|881.1|ICD9CM|Open wound of elbow, forearm, and wrist, complicated|Open wound of elbow, forearm, and wrist, complicated
C0160608|T037|AB|881.10|ICD9CM|Open wound forearm-compl|Open wound forearm-compl
C0160608|T037|PT|881.10|ICD9CM|Open wound of forearm, complicated|Open wound of forearm, complicated
C0160609|T037|AB|881.11|ICD9CM|Open wound elbow-complic|Open wound elbow-complic
C0160609|T037|PT|881.11|ICD9CM|Open wound of elbow, complicated|Open wound of elbow, complicated
C0160610|T037|PT|881.12|ICD9CM|Open wound of wrist, complicated|Open wound of wrist, complicated
C0160610|T037|AB|881.12|ICD9CM|Open wound wrist-complic|Open wound wrist-complic
C0160611|T037|HT|881.2|ICD9CM|Open wound of elbow, forearm, and wrist, with tendon involvement|Open wound of elbow, forearm, and wrist, with tendon involvement
C0160612|T037|AB|881.20|ICD9CM|Open wnd forearm w tendn|Open wnd forearm w tendn
C0160612|T037|PT|881.20|ICD9CM|Open wound of forearm, with tendon involvement|Open wound of forearm, with tendon involvement
C0160613|T037|PT|881.21|ICD9CM|Open wound of elbow, with tendon involvement|Open wound of elbow, with tendon involvement
C0160613|T037|AB|881.21|ICD9CM|Opn wound elbow w tendon|Opn wound elbow w tendon
C0160614|T037|PT|881.22|ICD9CM|Open wound of wrist, with tendon involvement|Open wound of wrist, with tendon involvement
C0160614|T037|AB|881.22|ICD9CM|Opn wound wrist w tendon|Opn wound wrist w tendon
C0160615|T037|HT|882|ICD9CM|Open wound of hand except finger(s) alone|Open wound of hand except finger(s) alone
C0160616|T037|AB|882.0|ICD9CM|Open wound of hand|Open wound of hand
C0160616|T037|PT|882.0|ICD9CM|Open wound of hand except finger(s) alone, without mention of complication|Open wound of hand except finger(s) alone, without mention of complication
C0160617|T037|PT|882.1|ICD9CM|Open wound of hand except finger(s) alone, complicated|Open wound of hand except finger(s) alone, complicated
C0160617|T037|AB|882.1|ICD9CM|Opn wound hand-complicat|Opn wound hand-complicat
C0160618|T037|AB|882.2|ICD9CM|Open wound hand w tendon|Open wound hand w tendon
C0160618|T037|PT|882.2|ICD9CM|Open wound of hand except finger(s) alone, with tendon involvement|Open wound of hand except finger(s) alone, with tendon involvement
C0555295|T037|HT|883|ICD9CM|Open wound of finger(s)|Open wound of finger(s)
C0273365|T037|AB|883.0|ICD9CM|Open wound of finger|Open wound of finger
C0273365|T037|PT|883.0|ICD9CM|Open wound of finger(s), without mention of complication|Open wound of finger(s), without mention of complication
C0160621|T037|AB|883.1|ICD9CM|Open wound finger-compl|Open wound finger-compl
C0160621|T037|PT|883.1|ICD9CM|Open wound of finger(s), complicated|Open wound of finger(s), complicated
C0160622|T037|AB|883.2|ICD9CM|Open wnd finger w tendon|Open wnd finger w tendon
C0160622|T037|PT|883.2|ICD9CM|Open wound of finger(s), with tendon involvement|Open wound of finger(s), with tendon involvement
C1744615|T037|HT|884|ICD9CM|Multiple and unspecified open wound of upper limb|Multiple and unspecified open wound of upper limb
C0160623|T037|PT|884.0|ICD9CM|Multiple and unspecified open wound of upper limb, without mention of complication|Multiple and unspecified open wound of upper limb, without mention of complication
C0160623|T037|AB|884.0|ICD9CM|Open wound arm mult/NOS|Open wound arm mult/NOS
C0160625|T037|PT|884.1|ICD9CM|Multiple and unspecified open wound of upper limb, complicated|Multiple and unspecified open wound of upper limb, complicated
C0160625|T037|AB|884.1|ICD9CM|Open wound arm NOS-compl|Open wound arm NOS-compl
C0160626|T037|PT|884.2|ICD9CM|Multiple and unspecified open wound of upper limb, with tendon involvement|Multiple and unspecified open wound of upper limb, with tendon involvement
C0160626|T037|AB|884.2|ICD9CM|Opn wnd arm NOS w tendon|Opn wnd arm NOS w tendon
C0160627|T037|HT|885|ICD9CM|Traumatic amputation of thumb (complete) (partial)|Traumatic amputation of thumb (complete) (partial)
C0433638|T037|AB|885.0|ICD9CM|Amputation thumb|Amputation thumb
C0433638|T037|PT|885.0|ICD9CM|Traumatic amputation of thumb (complete)(partial), without mention of complication|Traumatic amputation of thumb (complete)(partial), without mention of complication
C0160629|T037|AB|885.1|ICD9CM|Amputation thumb-compl|Amputation thumb-compl
C0160629|T037|PT|885.1|ICD9CM|Traumatic amputation of thumb (complete)(partial), complicated|Traumatic amputation of thumb (complete)(partial), complicated
C0160630|T037|HT|886|ICD9CM|Traumatic amputation of other finger(s) (complete) (partial)|Traumatic amputation of other finger(s) (complete) (partial)
C0160631|T037|AB|886.0|ICD9CM|Amputation finger|Amputation finger
C0160631|T037|PT|886.0|ICD9CM|Traumatic amputation of other finger(s) (complete) (partial), without mention of complication|Traumatic amputation of other finger(s) (complete) (partial), without mention of complication
C0160632|T037|AB|886.1|ICD9CM|Amputation finger-compl|Amputation finger-compl
C0160632|T037|PT|886.1|ICD9CM|Traumatic amputation of other finger(s) (complete) (partial), complicated|Traumatic amputation of other finger(s) (complete) (partial), complicated
C0160633|T037|HT|887|ICD9CM|Traumatic amputation of arm and hand (complete) (partial)|Traumatic amputation of arm and hand (complete) (partial)
C0160634|T037|AB|887.0|ICD9CM|Amput below elb, unilat|Amput below elb, unilat
C0273389|T037|AB|887.1|ICD9CM|Amp below elb, unil-comp|Amp below elb, unil-comp
C0273389|T037|PT|887.1|ICD9CM|Traumatic amputation of arm and hand (complete) (partial), unilateral, below elbow, complicated|Traumatic amputation of arm and hand (complete) (partial), unilateral, below elbow, complicated
C0160636|T037|AB|887.2|ICD9CM|Amput abv elbow, unilat|Amput abv elbow, unilat
C0273387|T037|AB|887.3|ICD9CM|Amput abv elb, unil-comp|Amput abv elb, unil-comp
C0160638|T037|AB|887.4|ICD9CM|Amputat arm, unilat NOS|Amputat arm, unilat NOS
C0160639|T037|AB|887.5|ICD9CM|Amput arm, unil NOS-comp|Amput arm, unil NOS-comp
C0160640|T037|AB|887.6|ICD9CM|Amputation arm, bilat|Amputation arm, bilat
C0160641|T037|AB|887.7|ICD9CM|Amputat arm, bilat-compl|Amputat arm, bilat-compl
C0160641|T037|PT|887.7|ICD9CM|Traumatic amputation of arm and hand (complete) (partial), bilateral [any level], complicated|Traumatic amputation of arm and hand (complete) (partial), bilateral [any level], complicated
C0160643|T037|HT|890|ICD9CM|Open wound of hip and thigh|Open wound of hip and thigh
C0178323|T037|HT|890-897.99|ICD9CM|OPEN WOUND OF LOWER LIMB|OPEN WOUND OF LOWER LIMB
C1279573|T037|PT|890.0|ICD9CM|Open wound of hip and thigh, without mention of complication|Open wound of hip and thigh, without mention of complication
C1279573|T037|AB|890.0|ICD9CM|Open wound of hip/thigh|Open wound of hip/thigh
C0160644|T037|AB|890.1|ICD9CM|Open wnd hip/thigh-compl|Open wnd hip/thigh-compl
C0160644|T037|PT|890.1|ICD9CM|Open wound of hip and thigh, complicated|Open wound of hip and thigh, complicated
C0160645|T037|PT|890.2|ICD9CM|Open wound of hip and thigh, with tendon involvement|Open wound of hip and thigh, with tendon involvement
C0160645|T037|AB|890.2|ICD9CM|Opn wnd hip/thigh w tend|Opn wnd hip/thigh w tend
C1744616|T037|HT|891|ICD9CM|Open wound of knee, leg [except thigh], and ankle|Open wound of knee, leg [except thigh], and ankle
C0160647|T037|AB|891.0|ICD9CM|Open wnd knee/leg/ankle|Open wnd knee/leg/ankle
C0160647|T037|PT|891.0|ICD9CM|Open wound of knee, leg [except thigh], and ankle, without mention of complication|Open wound of knee, leg [except thigh], and ankle, without mention of complication
C0160648|T037|AB|891.1|ICD9CM|Open wnd knee/leg-compl|Open wnd knee/leg-compl
C0160648|T037|PT|891.1|ICD9CM|Open wound of knee, leg [except thigh], and ankle, complicated|Open wound of knee, leg [except thigh], and ankle, complicated
C0160649|T037|PT|891.2|ICD9CM|Open wound of knee, leg [except thigh], and ankle, with tendon involvement|Open wound of knee, leg [except thigh], and ankle, with tendon involvement
C0160649|T037|AB|891.2|ICD9CM|Opn wnd knee/leg w tendn|Opn wnd knee/leg w tendn
C0160650|T037|HT|892|ICD9CM|Open wound of foot except toe(s) alone|Open wound of foot except toe(s) alone
C0160651|T037|AB|892.0|ICD9CM|Open wound of foot|Open wound of foot
C0160651|T037|PT|892.0|ICD9CM|Open wound of foot except toe(s) alone, without mention of complication|Open wound of foot except toe(s) alone, without mention of complication
C0160652|T037|AB|892.1|ICD9CM|Open wound foot-compl|Open wound foot-compl
C0160652|T037|PT|892.1|ICD9CM|Open wound of foot except toe(s) alone, complicated|Open wound of foot except toe(s) alone, complicated
C0160653|T037|AB|892.2|ICD9CM|Open wound foot w tendon|Open wound foot w tendon
C0160653|T037|PT|892.2|ICD9CM|Open wound of foot except toe(s) alone, with tendon involvement|Open wound of foot except toe(s) alone, with tendon involvement
C0562512|T037|HT|893|ICD9CM|Open wound of toe(s)|Open wound of toe(s)
C0160655|T037|AB|893.0|ICD9CM|Open wound of toe|Open wound of toe
C0160655|T037|PT|893.0|ICD9CM|Open wound of toe(s), without mention of complication|Open wound of toe(s), without mention of complication
C0273412|T037|PT|893.1|ICD9CM|Open wound of toe(s), complicated|Open wound of toe(s), complicated
C0273412|T037|AB|893.1|ICD9CM|Open wound toe-compl|Open wound toe-compl
C0273413|T037|PT|893.2|ICD9CM|Open wound of toe(s), with tendon involvement|Open wound of toe(s), with tendon involvement
C0273413|T037|AB|893.2|ICD9CM|Open wound toe w tendon|Open wound toe w tendon
C0160658|T037|HT|894|ICD9CM|Multiple and unspecified open wound of lower limb|Multiple and unspecified open wound of lower limb
C1812613|T037|PT|894.0|ICD9CM|Multiple and unspecified open wound of lower limb, without mention of complication|Multiple and unspecified open wound of lower limb, without mention of complication
C1812613|T037|AB|894.0|ICD9CM|Open wound of leg NEC|Open wound of leg NEC
C0160660|T037|PT|894.1|ICD9CM|Multiple and unspecified open wound of lower limb, complicated|Multiple and unspecified open wound of lower limb, complicated
C0160660|T037|AB|894.1|ICD9CM|Open wound leg NEC-compl|Open wound leg NEC-compl
C0160661|T037|PT|894.2|ICD9CM|Multiple and unspecified open wound of lower limb, with tendon involvement|Multiple and unspecified open wound of lower limb, with tendon involvement
C0160661|T037|AB|894.2|ICD9CM|Opn wnd leg NEC w tendon|Opn wnd leg NEC w tendon
C1744632|T037|HT|895|ICD9CM|Traumatic amputation of toe(s) (complete) (partial)|Traumatic amputation of toe(s) (complete) (partial)
C0160662|T037|AB|895.0|ICD9CM|Amputation toe|Amputation toe
C0160662|T037|PT|895.0|ICD9CM|Traumatic amputation of toe(s) (complete) (partial), without mention of complication|Traumatic amputation of toe(s) (complete) (partial), without mention of complication
C0433625|T037|AB|895.1|ICD9CM|Amputation toe-complicat|Amputation toe-complicat
C0433625|T037|PT|895.1|ICD9CM|Traumatic amputation of toe(s) (complete) (partial), complicated|Traumatic amputation of toe(s) (complete) (partial), complicated
C0160665|T037|HT|896|ICD9CM|Traumatic amputation of foot (complete) (partial)|Traumatic amputation of foot (complete) (partial)
C1366330|T037|AB|896.0|ICD9CM|Amputation foot, unilat|Amputation foot, unilat
C1366330|T037|PT|896.0|ICD9CM|Traumatic amputation of foot (complete) (partial), unilateral, without mention of complication|Traumatic amputation of foot (complete) (partial), unilateral, without mention of complication
C0273417|T037|AB|896.1|ICD9CM|Amput foot, unilat-compl|Amput foot, unilat-compl
C0273417|T037|PT|896.1|ICD9CM|Traumatic amputation of foot (complete) (partial), unilateral, complicated|Traumatic amputation of foot (complete) (partial), unilateral, complicated
C0160668|T037|AB|896.2|ICD9CM|Amputation foot, bilat|Amputation foot, bilat
C0160668|T037|PT|896.2|ICD9CM|Traumatic amputation of foot (complete) (partial), bilateral, without mention of complication|Traumatic amputation of foot (complete) (partial), bilateral, without mention of complication
C0273419|T037|AB|896.3|ICD9CM|Amputat foot, bilat-comp|Amputat foot, bilat-comp
C0273419|T037|PT|896.3|ICD9CM|Traumatic amputation of foot (complete) (partial), bilateral, complicated|Traumatic amputation of foot (complete) (partial), bilateral, complicated
C0160675|T037|HT|897|ICD9CM|Traumatic amputation of leg(s) (complete) (partial)|Traumatic amputation of leg(s) (complete) (partial)
C0160671|T037|AB|897.0|ICD9CM|Amput below knee, unilat|Amput below knee, unilat
C0160672|T037|AB|897.1|ICD9CM|Amputat bk, unilat-compl|Amputat bk, unilat-compl
C0160672|T037|PT|897.1|ICD9CM|Traumatic amputation of leg(s) (complete) (partial), unilateral, below knee, complicated|Traumatic amputation of leg(s) (complete) (partial), unilateral, below knee, complicated
C0160673|T037|AB|897.2|ICD9CM|Amput above knee, unilat|Amput above knee, unilat
C0160674|T037|AB|897.3|ICD9CM|Amput abv kn, unil-compl|Amput abv kn, unil-compl
C0160674|T037|PT|897.3|ICD9CM|Traumatic amputation of leg(s) (complete) (partial), unilateral, at or above knee, complicated|Traumatic amputation of leg(s) (complete) (partial), unilateral, at or above knee, complicated
C0478347|T037|AB|897.4|ICD9CM|Amputat leg, unilat NOS|Amputat leg, unilat NOS
C0160676|T037|AB|897.5|ICD9CM|Amput leg, unil NOS-comp|Amput leg, unil NOS-comp
C0160676|T037|PT|897.5|ICD9CM|Traumatic amputation of leg(s) (complete) (partial), unilateral, level not specified, complicated|Traumatic amputation of leg(s) (complete) (partial), unilateral, level not specified, complicated
C0160677|T037|AB|897.6|ICD9CM|Amputation leg, bilat|Amputation leg, bilat
C0160678|T037|AB|897.7|ICD9CM|Amputat leg, bilat-compl|Amputat leg, bilat-compl
C0160678|T037|PT|897.7|ICD9CM|Traumatic amputation of leg(s) (complete) (partial), bilateral [any level], complicated|Traumatic amputation of leg(s) (complete) (partial), bilateral [any level], complicated
C0160679|T037|HT|900|ICD9CM|Injury to blood vessels of head and neck|Injury to blood vessels of head and neck
C0178324|T037|HT|900-904.99|ICD9CM|INJURY TO BLOOD VESSELS|INJURY TO BLOOD VESSELS
C0160680|T037|HT|900.0|ICD9CM|Injury to carotid artery|Injury to carotid artery
C0160680|T037|AB|900.00|ICD9CM|Injur carotid artery NOS|Injur carotid artery NOS
C0160680|T037|PT|900.00|ICD9CM|Injury to carotid artery, unspecified|Injury to carotid artery, unspecified
C0160681|T037|AB|900.01|ICD9CM|Inj common carotid arter|Inj common carotid arter
C0160681|T037|PT|900.01|ICD9CM|Injury to common carotid artery|Injury to common carotid artery
C0160682|T037|AB|900.02|ICD9CM|Inj external carotid art|Inj external carotid art
C0160682|T037|PT|900.02|ICD9CM|Injury to external carotid artery|Injury to external carotid artery
C0160683|T037|AB|900.03|ICD9CM|Inj internal carotid art|Inj internal carotid art
C0160683|T037|PT|900.03|ICD9CM|Injury to internal carotid artery|Injury to internal carotid artery
C0160684|T037|AB|900.1|ICD9CM|Inj internl jugular vein|Inj internl jugular vein
C0160684|T037|PT|900.1|ICD9CM|Injury to internal jugular vein|Injury to internal jugular vein
C0160685|T037|HT|900.8|ICD9CM|Injury to other specified blood vessels of head and neck|Injury to other specified blood vessels of head and neck
C0160686|T037|AB|900.81|ICD9CM|Inj extern jugular vein|Inj extern jugular vein
C0160686|T037|PT|900.81|ICD9CM|Injury to external jugular vein|Injury to external jugular vein
C0160687|T037|AB|900.82|ICD9CM|Inj mlt head/neck vessel|Inj mlt head/neck vessel
C0160687|T037|PT|900.82|ICD9CM|Injury to multiple blood vessels of head and neck|Injury to multiple blood vessels of head and neck
C0160685|T037|AB|900.89|ICD9CM|Inj head/neck vessel NEC|Inj head/neck vessel NEC
C0160685|T037|PT|900.89|ICD9CM|Injury to other specified blood vessels of head and neck|Injury to other specified blood vessels of head and neck
C0160679|T037|AB|900.9|ICD9CM|Inj head/neck vessel NOS|Inj head/neck vessel NOS
C0160679|T037|PT|900.9|ICD9CM|Injury to unspecified blood vessel of head and neck|Injury to unspecified blood vessel of head and neck
C0160689|T037|HT|901|ICD9CM|Injury to blood vessels of thorax|Injury to blood vessels of thorax
C0160690|T037|AB|901.0|ICD9CM|Injury thoracic aorta|Injury thoracic aorta
C0160690|T037|PT|901.0|ICD9CM|Injury to thoracic aorta|Injury to thoracic aorta
C0495833|T037|AB|901.1|ICD9CM|Inj innomin/subclav art|Inj innomin/subclav art
C0495833|T037|PT|901.1|ICD9CM|Injury to innominate and subclavian arteries|Injury to innominate and subclavian arteries
C0160692|T037|AB|901.2|ICD9CM|Inj superior vena cava|Inj superior vena cava
C0160692|T037|PT|901.2|ICD9CM|Injury to superior vena cava|Injury to superior vena cava
C0160693|T037|AB|901.3|ICD9CM|Inj innomin/subclav vein|Inj innomin/subclav vein
C0160693|T037|PT|901.3|ICD9CM|Injury to innominate and subclavian veins|Injury to innominate and subclavian veins
C0273454|T037|HT|901.4|ICD9CM|Injury to pulmonary blood vessels|Injury to pulmonary blood vessels
C0273454|T037|AB|901.40|ICD9CM|Inj pulmonary vessel NOS|Inj pulmonary vessel NOS
C0273454|T037|PT|901.40|ICD9CM|Injury to pulmonary vessel(s), unspecified|Injury to pulmonary vessel(s), unspecified
C0160696|T037|AB|901.41|ICD9CM|Injury pulmonary artery|Injury pulmonary artery
C0160696|T037|PT|901.41|ICD9CM|Injury to pulmonary artery|Injury to pulmonary artery
C0160697|T037|AB|901.42|ICD9CM|Injury pulmonary vein|Injury pulmonary vein
C0160697|T037|PT|901.42|ICD9CM|Injury to pulmonary vein|Injury to pulmonary vein
C0160698|T037|HT|901.8|ICD9CM|Injury to other specified blood vessels of thorax|Injury to other specified blood vessels of thorax
C0392044|T037|AB|901.81|ICD9CM|Inj intercostal art/vein|Inj intercostal art/vein
C0392044|T037|PT|901.81|ICD9CM|Injury to intercostal artery or vein|Injury to intercostal artery or vein
C0160700|T037|AB|901.82|ICD9CM|Inj int mammary art/vein|Inj int mammary art/vein
C0160700|T037|PT|901.82|ICD9CM|Injury to internal mammary artery or vein|Injury to internal mammary artery or vein
C0160701|T037|AB|901.83|ICD9CM|Inj mult thoracic vessel|Inj mult thoracic vessel
C0160701|T037|PT|901.83|ICD9CM|Injury to multiple blood vessels of thorax|Injury to multiple blood vessels of thorax
C0160698|T037|AB|901.89|ICD9CM|Inj thoracic vessel NEC|Inj thoracic vessel NEC
C0160698|T037|PT|901.89|ICD9CM|Injury to other specified blood vessels of thorax|Injury to other specified blood vessels of thorax
C0160689|T037|AB|901.9|ICD9CM|Inj thoracic vessel NOS|Inj thoracic vessel NOS
C0160689|T037|PT|901.9|ICD9CM|Injury to unspecified blood vessel of thorax|Injury to unspecified blood vessel of thorax
C0160703|T037|HT|902|ICD9CM|Injury to blood vessels of abdomen and pelvis|Injury to blood vessels of abdomen and pelvis
C0160704|T037|AB|902.0|ICD9CM|Injury abdominal aorta|Injury abdominal aorta
C0160704|T037|PT|902.0|ICD9CM|Injury to abdominal aorta|Injury to abdominal aorta
C0160705|T037|HT|902.1|ICD9CM|Injury to inferior vena cava|Injury to inferior vena cava
C0160705|T037|AB|902.10|ICD9CM|Inj infer vena cava NOS|Inj infer vena cava NOS
C0160705|T037|PT|902.10|ICD9CM|Injury to inferior vena cava, unspecified|Injury to inferior vena cava, unspecified
C0160706|T037|AB|902.11|ICD9CM|Injury hepatic veins|Injury hepatic veins
C0160706|T037|PT|902.11|ICD9CM|Injury to hepatic veins|Injury to hepatic veins
C0160707|T037|AB|902.19|ICD9CM|Inj infer vena cava NEC|Inj infer vena cava NEC
C0160707|T037|PT|902.19|ICD9CM|Injury to inferior vena cava, other|Injury to inferior vena cava, other
C0160708|T037|HT|902.2|ICD9CM|Injury to celiac and mesenteric arteries|Injury to celiac and mesenteric arteries
C0160708|T037|AB|902.20|ICD9CM|Inj celiac/mesen art NOS|Inj celiac/mesen art NOS
C0160708|T037|PT|902.20|ICD9CM|Injury to celiac and mesenteric arteries, unspecified|Injury to celiac and mesenteric arteries, unspecified
C0160709|T037|AB|902.21|ICD9CM|Injury gastric artery|Injury gastric artery
C0160709|T037|PT|902.21|ICD9CM|Injury to gastric artery|Injury to gastric artery
C0160710|T037|AB|902.22|ICD9CM|Injury hepatic artery|Injury hepatic artery
C0160710|T037|PT|902.22|ICD9CM|Injury to hepatic artery|Injury to hepatic artery
C0160711|T037|AB|902.23|ICD9CM|Injury splenic artery|Injury splenic artery
C0160711|T037|PT|902.23|ICD9CM|Injury to splenic artery|Injury to splenic artery
C0160712|T037|AB|902.24|ICD9CM|Injury celiac axis NEC|Injury celiac axis NEC
C0160712|T037|PT|902.24|ICD9CM|Injury to other specified branches of celiac axis|Injury to other specified branches of celiac axis
C0273463|T037|AB|902.25|ICD9CM|Inj super mesenteric art|Inj super mesenteric art
C0273463|T037|PT|902.25|ICD9CM|Injury to superior mesenteric artery (trunk)|Injury to superior mesenteric artery (trunk)
C0160714|T037|AB|902.26|ICD9CM|Inj brnch sup mesent art|Inj brnch sup mesent art
C0160714|T037|PT|902.26|ICD9CM|Injury to primary branches of superior mesenteric artery|Injury to primary branches of superior mesenteric artery
C0160715|T037|AB|902.27|ICD9CM|Inj infer mesenteric art|Inj infer mesenteric art
C0160715|T037|PT|902.27|ICD9CM|Injury to inferior mesenteric artery|Injury to inferior mesenteric artery
C0160716|T037|AB|902.29|ICD9CM|Inj mesenteric vess NEC|Inj mesenteric vess NEC
C0160716|T037|PT|902.29|ICD9CM|Injury to celiac and mesenteric arteries, other|Injury to celiac and mesenteric arteries, other
C0160717|T037|HT|902.3|ICD9CM|Injury to portal and splenic veins|Injury to portal and splenic veins
C0160718|T037|AB|902.31|ICD9CM|Inj superior mesent vein|Inj superior mesent vein
C0160718|T037|PT|902.31|ICD9CM|Injury to superior mesenteric vein and primary subdivisions|Injury to superior mesenteric vein and primary subdivisions
C0160719|T037|AB|902.32|ICD9CM|Inj inferior mesent vein|Inj inferior mesent vein
C0160719|T037|PT|902.32|ICD9CM|Injury to inferior mesenteric vein|Injury to inferior mesenteric vein
C0160720|T037|AB|902.33|ICD9CM|Injury portal vein|Injury portal vein
C0160720|T037|PT|902.33|ICD9CM|Injury to portal vein|Injury to portal vein
C0160721|T037|AB|902.34|ICD9CM|Injury splenic vein|Injury splenic vein
C0160721|T037|PT|902.34|ICD9CM|Injury to splenic vein|Injury to splenic vein
C0160722|T037|AB|902.39|ICD9CM|Inj port/splen vess NEC|Inj port/splen vess NEC
C0160722|T037|PT|902.39|ICD9CM|Injury to portal and splenic veins, other|Injury to portal and splenic veins, other
C0160723|T037|HT|902.4|ICD9CM|Injury to renal blood vessels|Injury to renal blood vessels
C0160723|T037|AB|902.40|ICD9CM|Injury renal vessel NOS|Injury renal vessel NOS
C0160723|T037|PT|902.40|ICD9CM|Injury to renal vessel(s), unspecified|Injury to renal vessel(s), unspecified
C0160725|T037|AB|902.41|ICD9CM|Injury renal artery|Injury renal artery
C0160725|T037|PT|902.41|ICD9CM|Injury to renal artery|Injury to renal artery
C0160726|T037|AB|902.42|ICD9CM|Injury renal vein|Injury renal vein
C0160726|T037|PT|902.42|ICD9CM|Injury to renal vein|Injury to renal vein
C0160727|T037|AB|902.49|ICD9CM|Injury renal vessel NEC|Injury renal vessel NEC
C0160727|T037|PT|902.49|ICD9CM|Injury to renal blood vessels, other|Injury to renal blood vessels, other
C0160728|T037|HT|902.5|ICD9CM|Injury to iliac blood vessels|Injury to iliac blood vessels
C0160728|T037|AB|902.50|ICD9CM|Injury iliac vessel NOS|Injury iliac vessel NOS
C0160728|T037|PT|902.50|ICD9CM|Injury to iliac vessel(s), unspecified|Injury to iliac vessel(s), unspecified
C0160730|T037|AB|902.51|ICD9CM|Inj hypogastric artery|Inj hypogastric artery
C0160730|T037|PT|902.51|ICD9CM|Injury to hypogastric artery|Injury to hypogastric artery
C0160731|T037|AB|902.52|ICD9CM|Injury hypogastric vein|Injury hypogastric vein
C0160731|T037|PT|902.52|ICD9CM|Injury to hypogastric vein|Injury to hypogastric vein
C0160732|T037|AB|902.53|ICD9CM|Injury iliac artery|Injury iliac artery
C0160732|T037|PT|902.53|ICD9CM|Injury to iliac artery|Injury to iliac artery
C0160733|T037|AB|902.54|ICD9CM|Injury iliac vein|Injury iliac vein
C0160733|T037|PT|902.54|ICD9CM|Injury to iliac vein|Injury to iliac vein
C0160734|T037|PT|902.55|ICD9CM|Injury to uterine artery|Injury to uterine artery
C0160734|T037|AB|902.55|ICD9CM|Injury uterine artery|Injury uterine artery
C0160735|T037|PT|902.56|ICD9CM|Injury to uterine vein|Injury to uterine vein
C0160735|T037|AB|902.56|ICD9CM|Injury uterine vein|Injury uterine vein
C0160736|T037|AB|902.59|ICD9CM|Injury iliac vessel NEC|Injury iliac vessel NEC
C0160736|T037|PT|902.59|ICD9CM|Injury to iliac blood vessels, other|Injury to iliac blood vessels, other
C0160737|T037|HT|902.8|ICD9CM|Injury to other specified blood vessels of abdomen and pelvis|Injury to other specified blood vessels of abdomen and pelvis
C0160738|T037|AB|902.81|ICD9CM|Injury ovarian artery|Injury ovarian artery
C0160738|T037|PT|902.81|ICD9CM|Injury to ovarian artery|Injury to ovarian artery
C0160739|T037|AB|902.82|ICD9CM|Injury ovarian vein|Injury ovarian vein
C0160739|T037|PT|902.82|ICD9CM|Injury to ovarian vein|Injury to ovarian vein
C0160740|T037|AB|902.87|ICD9CM|Inj mult abd/pelv vessel|Inj mult abd/pelv vessel
C0160740|T037|PT|902.87|ICD9CM|Injury to multiple blood vessels of abdomen and pelvis|Injury to multiple blood vessels of abdomen and pelvis
C0160737|T037|AB|902.89|ICD9CM|Inj abdominal vessel NEC|Inj abdominal vessel NEC
C0160737|T037|PT|902.89|ICD9CM|Injury to other specified blood vessels of abdomen and pelvis|Injury to other specified blood vessels of abdomen and pelvis
C0160703|T037|AB|902.9|ICD9CM|Inj abdominal vessel NOS|Inj abdominal vessel NOS
C0160703|T037|PT|902.9|ICD9CM|Injury to unspecified blood vessel of abdomen and pelvis|Injury to unspecified blood vessel of abdomen and pelvis
C0160742|T037|HT|903|ICD9CM|Injury to blood vessels of upper extremity|Injury to blood vessels of upper extremity
C0273471|T037|HT|903.0|ICD9CM|Injury to axillary blood vessels|Injury to axillary blood vessels
C0273471|T037|AB|903.00|ICD9CM|Inj axillary vessel NOS|Inj axillary vessel NOS
C0273471|T037|PT|903.00|ICD9CM|Injury to axillary vessel(s), unspecified|Injury to axillary vessel(s), unspecified
C0160745|T037|AB|903.01|ICD9CM|Injury axillary artery|Injury axillary artery
C0160745|T037|PT|903.01|ICD9CM|Injury to axillary artery|Injury to axillary artery
C0160746|T037|AB|903.02|ICD9CM|Injury axillary vein|Injury axillary vein
C0160746|T037|PT|903.02|ICD9CM|Injury to axillary vein|Injury to axillary vein
C0434195|T037|AB|903.1|ICD9CM|Injury brachial vessels|Injury brachial vessels
C0434195|T037|PT|903.1|ICD9CM|Injury to brachial blood vessels|Injury to brachial blood vessels
C0160748|T037|AB|903.2|ICD9CM|Injury radial vessels|Injury radial vessels
C0160748|T037|PT|903.2|ICD9CM|Injury to radial blood vessels|Injury to radial blood vessels
C0160749|T037|PT|903.3|ICD9CM|Injury to ulnar blood vessels|Injury to ulnar blood vessels
C0160749|T037|AB|903.3|ICD9CM|Injury ulnar vessels|Injury ulnar vessels
C0160750|T037|AB|903.4|ICD9CM|Injury palmar artery|Injury palmar artery
C0160750|T037|PT|903.4|ICD9CM|Injury to palmar artery|Injury to palmar artery
C0160751|T037|AB|903.5|ICD9CM|Injury finger vessels|Injury finger vessels
C0160751|T037|PT|903.5|ICD9CM|Injury to digital blood vessels|Injury to digital blood vessels
C0160752|T037|AB|903.8|ICD9CM|Injury arm vessels NEC|Injury arm vessels NEC
C0160752|T037|PT|903.8|ICD9CM|Injury to other specified blood vessels of upper extremity|Injury to other specified blood vessels of upper extremity
C0160742|T037|AB|903.9|ICD9CM|Injury arm vessel NOS|Injury arm vessel NOS
C0160742|T037|PT|903.9|ICD9CM|Injury to unspecified blood vessel of upper extremity|Injury to unspecified blood vessel of upper extremity
C0160754|T037|HT|904|ICD9CM|Injury to blood vessels of lower extremity and unspecified sites|Injury to blood vessels of lower extremity and unspecified sites
C0160755|T037|AB|904.0|ICD9CM|Inj common femoral arter|Inj common femoral arter
C0160755|T037|PT|904.0|ICD9CM|Injury to common femoral artery|Injury to common femoral artery
C0160756|T037|AB|904.1|ICD9CM|Inj superfic femoral art|Inj superfic femoral art
C0160756|T037|PT|904.1|ICD9CM|Injury to superficial femoral artery|Injury to superficial femoral artery
C0160757|T037|AB|904.2|ICD9CM|Injury femoral vein|Injury femoral vein
C0160757|T037|PT|904.2|ICD9CM|Injury to femoral veins|Injury to femoral veins
C0160758|T037|AB|904.3|ICD9CM|Injury saphenous vein|Injury saphenous vein
C0160758|T037|PT|904.3|ICD9CM|Injury to saphenous veins|Injury to saphenous veins
C0273480|T037|HT|904.4|ICD9CM|Injury to popliteal blood vessels|Injury to popliteal blood vessels
C0273480|T037|AB|904.40|ICD9CM|Inj popliteal vessel NOS|Inj popliteal vessel NOS
C0273480|T037|PT|904.40|ICD9CM|Injury to popliteal vessel(s), unspecified|Injury to popliteal vessel(s), unspecified
C0160761|T037|AB|904.41|ICD9CM|Injury popliteal artery|Injury popliteal artery
C0160761|T037|PT|904.41|ICD9CM|Injury to popliteal artery|Injury to popliteal artery
C0160762|T037|AB|904.42|ICD9CM|Injury popliteal vein|Injury popliteal vein
C0160762|T037|PT|904.42|ICD9CM|Injury to popliteal vein|Injury to popliteal vein
C0160763|T037|HT|904.5|ICD9CM|Injury to tibial blood vessels|Injury to tibial blood vessels
C0160763|T037|AB|904.50|ICD9CM|Injury tibial vessel NOS|Injury tibial vessel NOS
C0160763|T037|PT|904.50|ICD9CM|Injury to tibial vessel(s), unspecified|Injury to tibial vessel(s), unspecified
C0160765|T037|AB|904.51|ICD9CM|Inj anter tibial artery|Inj anter tibial artery
C0160765|T037|PT|904.51|ICD9CM|Injury to anterior tibial artery|Injury to anterior tibial artery
C0160766|T037|AB|904.52|ICD9CM|Inj anterior tibial vein|Inj anterior tibial vein
C0160766|T037|PT|904.52|ICD9CM|Injury to anterior tibial vein|Injury to anterior tibial vein
C0160767|T037|AB|904.53|ICD9CM|Inj post tibial artery|Inj post tibial artery
C0160767|T037|PT|904.53|ICD9CM|Injury to posterior tibial artery|Injury to posterior tibial artery
C0160768|T037|AB|904.54|ICD9CM|Inj post tibial vein|Inj post tibial vein
C0160768|T037|PT|904.54|ICD9CM|Injury to posterior tibial vein|Injury to posterior tibial vein
C0160769|T037|AB|904.6|ICD9CM|Inj deep plantar vessel|Inj deep plantar vessel
C0160769|T037|PT|904.6|ICD9CM|Injury to deep plantar blood vessels|Injury to deep plantar blood vessels
C0160770|T037|AB|904.7|ICD9CM|Injury leg vessels NEC|Injury leg vessels NEC
C0160770|T037|PT|904.7|ICD9CM|Injury to other specified blood vessels of lower extremity|Injury to other specified blood vessels of lower extremity
C0273478|T037|AB|904.8|ICD9CM|Injury leg vessel NOS|Injury leg vessel NOS
C0273478|T037|PT|904.8|ICD9CM|Injury to unspecified blood vessel of lower extremity|Injury to unspecified blood vessel of lower extremity
C0178324|T037|AB|904.9|ICD9CM|Blood vessel injury NOS|Blood vessel injury NOS
C0178324|T037|PT|904.9|ICD9CM|Injury to blood vessels of unspecified site|Injury to blood vessels of unspecified site
C0160773|T046|HT|905|ICD9CM|Late effects of musculoskeletal and connective tissue injuries|Late effects of musculoskeletal and connective tissue injuries
C0178325|T037|HT|905-909.99|ICD9CM|LATE EFFECTS OF INJURIES, POISONINGS, TOXIC EFFECTS, AND OTHER EXTERNAL CAUSES|LATE EFFECTS OF INJURIES, POISONINGS, TOXIC EFFECTS, AND OTHER EXTERNAL CAUSES
C0160774|T046|AB|905.0|ICD9CM|Late effec skull/face fx|Late effec skull/face fx
C0160774|T046|PT|905.0|ICD9CM|Late effect of fracture of skull and face bones|Late effect of fracture of skull and face bones
C1331611|T046|AB|905.1|ICD9CM|Late eff spine/trunk fx|Late eff spine/trunk fx
C1331611|T046|PT|905.1|ICD9CM|Late effect of fracture of spine and trunk without mention of spinal cord lesion|Late effect of fracture of spine and trunk without mention of spinal cord lesion
C0436099|T046|AB|905.2|ICD9CM|Late effect arm fx|Late effect arm fx
C0436099|T046|PT|905.2|ICD9CM|Late effect of fracture of upper extremities|Late effect of fracture of upper extremities
C0160777|T046|AB|905.3|ICD9CM|Late eff femoral neck fx|Late eff femoral neck fx
C0160777|T046|PT|905.3|ICD9CM|Late effect of fracture of neck of femur|Late effect of fracture of neck of femur
C0160778|T046|AB|905.4|ICD9CM|Late effect leg fx|Late effect leg fx
C0160778|T046|PT|905.4|ICD9CM|Late effect of fracture of lower extremities|Late effect of fracture of lower extremities
C0160779|T046|AB|905.5|ICD9CM|Late effect fracture NEC|Late effect fracture NEC
C0160779|T046|PT|905.5|ICD9CM|Late effect of fracture of multiple and unspecified bones|Late effect of fracture of multiple and unspecified bones
C0160780|T046|AB|905.6|ICD9CM|Late effect dislocation|Late effect dislocation
C0160780|T046|PT|905.6|ICD9CM|Late effect of dislocation|Late effect of dislocation
C0160781|T037|AB|905.7|ICD9CM|Late effec sprain/strain|Late effec sprain/strain
C0160781|T037|PT|905.7|ICD9CM|Late effect of sprain and strain without mention of tendon injury|Late effect of sprain and strain without mention of tendon injury
C0160782|T046|AB|905.8|ICD9CM|Late effec tendon injury|Late effec tendon injury
C0160782|T046|PT|905.8|ICD9CM|Late effect of tendon injury|Late effect of tendon injury
C0160783|T046|AB|905.9|ICD9CM|Late eff traumat amputat|Late eff traumat amputat
C0160783|T046|PT|905.9|ICD9CM|Late effect of traumatic amputation|Late effect of traumatic amputation
C0160784|T046|HT|906|ICD9CM|Late effects of injuries to skin and subcutaneous tissues|Late effects of injuries to skin and subcutaneous tissues
C0160785|T046|PT|906.0|ICD9CM|Late effect of open wound of head, neck, and trunk|Late effect of open wound of head, neck, and trunk
C0160785|T046|AB|906.0|ICD9CM|Lt eff opn wnd head/trnk|Lt eff opn wnd head/trnk
C0160786|T037|AB|906.1|ICD9CM|Late eff open wnd extrem|Late eff open wnd extrem
C0160786|T037|PT|906.1|ICD9CM|Late effect of open wound of extremities without mention of tendon injury|Late effect of open wound of extremities without mention of tendon injury
C0160787|T046|AB|906.2|ICD9CM|Late eff superficial inj|Late eff superficial inj
C0160787|T046|PT|906.2|ICD9CM|Late effect of superficial injury|Late effect of superficial injury
C0160788|T046|AB|906.3|ICD9CM|Late effect of contusion|Late effect of contusion
C0160788|T046|PT|906.3|ICD9CM|Late effect of contusion|Late effect of contusion
C0274276|T046|AB|906.4|ICD9CM|Late effect of crushing|Late effect of crushing
C0274276|T046|PT|906.4|ICD9CM|Late effect of crushing|Late effect of crushing
C0160790|T046|AB|906.5|ICD9CM|Late eff head/neck burn|Late eff head/neck burn
C0160790|T046|PT|906.5|ICD9CM|Late effect of burn of eye, face, head, and neck|Late effect of burn of eye, face, head, and neck
C0160791|T046|AB|906.6|ICD9CM|Late eff wrist/hand burn|Late eff wrist/hand burn
C0160791|T046|PT|906.6|ICD9CM|Late effect of burn of wrist and hand|Late effect of burn of wrist and hand
C0160792|T046|AB|906.7|ICD9CM|Late eff burn extrem NEC|Late eff burn extrem NEC
C0160792|T046|PT|906.7|ICD9CM|Late effect of burn of other extremities|Late effect of burn of other extremities
C0160793|T037|AB|906.8|ICD9CM|Late effect of burns NEC|Late effect of burns NEC
C0160793|T037|PT|906.8|ICD9CM|Late effect of burns of other specified sites|Late effect of burns of other specified sites
C0160794|T046|AB|906.9|ICD9CM|Late effect of burn NOS|Late effect of burn NOS
C0160794|T046|PT|906.9|ICD9CM|Late effect of burn of unspecified site|Late effect of burn of unspecified site
C0160795|T046|HT|907|ICD9CM|Late effects of injuries to the nervous system|Late effects of injuries to the nervous system
C0274278|T037|PT|907.0|ICD9CM|Late effect of intracranial injury without mention of skull fracture|Late effect of intracranial injury without mention of skull fracture
C0274278|T037|AB|907.0|ICD9CM|Lt eff intracranial inj|Lt eff intracranial inj
C0160796|T046|AB|907.1|ICD9CM|Late eff cran nerve inj|Late eff cran nerve inj
C0160796|T046|PT|907.1|ICD9CM|Late effect of injury to cranial nerve|Late effect of injury to cranial nerve
C0160797|T046|AB|907.2|ICD9CM|Late eff spinal cord inj|Late eff spinal cord inj
C0160797|T046|PT|907.2|ICD9CM|Late effect of spinal cord injury|Late effect of spinal cord injury
C0160798|T047|PT|907.3|ICD9CM|Late effect of injury to nerve root(s), spinal plexus(es), and other nerves of trunk|Late effect of injury to nerve root(s), spinal plexus(es), and other nerves of trunk
C0160798|T047|AB|907.3|ICD9CM|Lt eff nerv inj trnk NEC|Lt eff nerv inj trnk NEC
C0160799|T046|PT|907.4|ICD9CM|Late effect of injury to peripheral nerve of shoulder girdle and upper limb|Late effect of injury to peripheral nerve of shoulder girdle and upper limb
C0160799|T046|AB|907.4|ICD9CM|Lt eff nerv inj shld/arm|Lt eff nerv inj shld/arm
C0160800|T046|PT|907.5|ICD9CM|Late effect of injury to peripheral nerve of pelvic girdle and lower limb|Late effect of injury to peripheral nerve of pelvic girdle and lower limb
C0160800|T046|AB|907.5|ICD9CM|Lt eff nerv inj pelv/leg|Lt eff nerv inj pelv/leg
C0160801|T037|AB|907.9|ICD9CM|Late eff nerve inj NEC|Late eff nerve inj NEC
C0160801|T037|PT|907.9|ICD9CM|Late effect of injury to other and unspecified nerve|Late effect of injury to other and unspecified nerve
C0160802|T046|HT|908|ICD9CM|Late effects of other and unspecified injuries|Late effects of other and unspecified injuries
C0160803|T046|AB|908.0|ICD9CM|Late eff int injur chest|Late eff int injur chest
C0160803|T046|PT|908.0|ICD9CM|Late effect of internal injury to chest|Late effect of internal injury to chest
C0859827|T046|AB|908.1|ICD9CM|Late eff int inj abdomen|Late eff int inj abdomen
C0859827|T046|PT|908.1|ICD9CM|Late effect of internal injury to intra-abdominal organs|Late effect of internal injury to intra-abdominal organs
C0160805|T037|AB|908.2|ICD9CM|Late eff int injury NEC|Late eff int injury NEC
C0160805|T037|PT|908.2|ICD9CM|Late effect of internal injury to other internal organs|Late effect of internal injury to other internal organs
C0160806|T046|AB|908.3|ICD9CM|Late eff inj periph vess|Late eff inj periph vess
C0160806|T046|PT|908.3|ICD9CM|Late effect of injury to blood vessel of head, neck, and extremities|Late effect of injury to blood vessel of head, neck, and extremities
C0160807|T046|PT|908.4|ICD9CM|Late effect of injury to blood vessel of thorax, abdomen, and pelvis|Late effect of injury to blood vessel of thorax, abdomen, and pelvis
C0160807|T046|AB|908.4|ICD9CM|Lt eff inj thor/abd vess|Lt eff inj thor/abd vess
C0160808|T046|AB|908.5|ICD9CM|Late eff FB in orifice|Late eff FB in orifice
C0160808|T046|PT|908.5|ICD9CM|Late effect of foreign body in orifice|Late effect of foreign body in orifice
C0160809|T046|AB|908.6|ICD9CM|Late eff complic trauma|Late eff complic trauma
C0160809|T046|PT|908.6|ICD9CM|Late effect of certain complications of trauma|Late effect of certain complications of trauma
C1313863|T046|AB|908.9|ICD9CM|Late effect injury NOS|Late effect injury NOS
C1313863|T046|PT|908.9|ICD9CM|Late effect of unspecified injury|Late effect of unspecified injury
C0436115|T037|HT|909|ICD9CM|Late effects of other and unspecified external causes|Late effects of other and unspecified external causes
C0496180|T046|AB|909.0|ICD9CM|Late eff drug poisoning|Late eff drug poisoning
C0496180|T046|PT|909.0|ICD9CM|Late effect of poisoning due to drug, medicinal or biological substance|Late effect of poisoning due to drug, medicinal or biological substance
C0436114|T046|AB|909.1|ICD9CM|Late eff nonmed substanc|Late eff nonmed substanc
C0436114|T046|PT|909.1|ICD9CM|Late effect of toxic effects of nonmedical substances|Late effect of toxic effects of nonmedical substances
C0160814|T046|AB|909.2|ICD9CM|Late effect of radiation|Late effect of radiation
C0160814|T046|PT|909.2|ICD9CM|Late effect of radiation|Late effect of radiation
C3665468|T046|AB|909.3|ICD9CM|Late eff surg/med compl|Late eff surg/med compl
C3665468|T046|PT|909.3|ICD9CM|Late effect of complications of surgical and medical care|Late effect of complications of surgical and medical care
C0160816|T037|AB|909.4|ICD9CM|Late eff cert ext cause|Late eff cert ext cause
C0160816|T037|PT|909.4|ICD9CM|Late effect of certain other external causes|Late effect of certain other external causes
C0375668|T037|PT|909.5|ICD9CM|Late effect of adverse effect of drug, medicinal or biological substance|Late effect of adverse effect of drug, medicinal or biological substance
C0375668|T037|AB|909.5|ICD9CM|Lte efct advrs efct drug|Lte efct advrs efct drug
C2240395|T037|AB|909.9|ICD9CM|Late eff exter cause NEC|Late eff exter cause NEC
C2240395|T037|PT|909.9|ICD9CM|Late effect of other and unspecified external causes|Late effect of other and unspecified external causes
C0160818|T037|HT|910|ICD9CM|Superficial injury of face, neck, and scalp except eye|Superficial injury of face, neck, and scalp except eye
C0332671|T037|HT|910-919.99|ICD9CM|SUPERFICIAL INJURY|SUPERFICIAL INJURY
C0160819|T037|AB|910.0|ICD9CM|Abrasion head|Abrasion head
C0160819|T037|PT|910.0|ICD9CM|Abrasion or friction burn of face, neck, and scalp except eye, without mention of infection|Abrasion or friction burn of face, neck, and scalp except eye, without mention of infection
C0160820|T037|AB|910.1|ICD9CM|Abrasion head-infected|Abrasion head-infected
C0160820|T037|PT|910.1|ICD9CM|Abrasion or friction burn of face, neck, and scalp except eye, infected|Abrasion or friction burn of face, neck, and scalp except eye, infected
C0160821|T037|AB|910.2|ICD9CM|Blister head|Blister head
C0160821|T037|PT|910.2|ICD9CM|Blister of face, neck, and scalp except eye, without mention of infection|Blister of face, neck, and scalp except eye, without mention of infection
C0160822|T046|AB|910.3|ICD9CM|Blister head-infected|Blister head-infected
C0160822|T046|PT|910.3|ICD9CM|Blister of face, neck, and scalp except eye, infected|Blister of face, neck, and scalp except eye, infected
C0160823|T037|AB|910.4|ICD9CM|Insect bite head|Insect bite head
C0160823|T037|PT|910.4|ICD9CM|Insect bite, nonvenomous of face, neck, and scalp except eye, without mention of infection|Insect bite, nonvenomous of face, neck, and scalp except eye, without mention of infection
C0160824|T037|AB|910.5|ICD9CM|Insect bite head-infect|Insect bite head-infect
C0160824|T037|PT|910.5|ICD9CM|Insect bite, nonvenomous of face, neck, and scalp except eye, infected|Insect bite, nonvenomous of face, neck, and scalp except eye, infected
C0160825|T037|AB|910.6|ICD9CM|Foreign body head|Foreign body head
C0160826|T037|AB|910.7|ICD9CM|Foreign body head-infect|Foreign body head-infect
C0160827|T037|PT|910.8|ICD9CM|Other and unspecified superficial injury of face, neck, and scalp, without mention of infection|Other and unspecified superficial injury of face, neck, and scalp, without mention of infection
C0160827|T037|AB|910.8|ICD9CM|Superfic inj head NEC|Superfic inj head NEC
C0160828|T037|PT|910.9|ICD9CM|Other and unspecified superficial injury of face, neck, and scalp, infected|Other and unspecified superficial injury of face, neck, and scalp, infected
C0160828|T037|AB|910.9|ICD9CM|Superf inj head NEC-inf|Superf inj head NEC-inf
C0160829|T037|HT|911|ICD9CM|Superficial injury of trunk|Superficial injury of trunk
C0160830|T037|PT|911.0|ICD9CM|Abrasion or friction burn of trunk, without mention of infection|Abrasion or friction burn of trunk, without mention of infection
C0160830|T037|AB|911.0|ICD9CM|Abrasion trunk|Abrasion trunk
C0160831|T037|PT|911.1|ICD9CM|Abrasion or friction burn of trunk, infected|Abrasion or friction burn of trunk, infected
C0160831|T037|AB|911.1|ICD9CM|Abrasion trunk-infected|Abrasion trunk-infected
C0160832|T037|PT|911.2|ICD9CM|Blister of trunk, without mention of infection|Blister of trunk, without mention of infection
C0160832|T037|AB|911.2|ICD9CM|Blister trunk|Blister trunk
C0160833|T037|PT|911.3|ICD9CM|Blister of trunk, infected|Blister of trunk, infected
C0160833|T037|AB|911.3|ICD9CM|Blister trunk-infected|Blister trunk-infected
C0273631|T037|AB|911.4|ICD9CM|Insect bite trunk|Insect bite trunk
C0273631|T037|PT|911.4|ICD9CM|Insect bite, nonvenomous of trunk, without mention of infection|Insect bite, nonvenomous of trunk, without mention of infection
C0273632|T037|AB|911.5|ICD9CM|Insect bite trunk-infec|Insect bite trunk-infec
C0273632|T037|PT|911.5|ICD9CM|Insect bite, nonvenomous of trunk, infected|Insect bite, nonvenomous of trunk, infected
C0160836|T037|AB|911.6|ICD9CM|Foreign body trunk|Foreign body trunk
C0160837|T037|AB|911.7|ICD9CM|Foreign body trunk-infec|Foreign body trunk-infec
C0160837|T037|PT|911.7|ICD9CM|Superficial foreign body (splinter) of trunk, without major open wound, infected|Superficial foreign body (splinter) of trunk, without major open wound, infected
C0840764|T037|PT|911.8|ICD9CM|Other and unspecified superficial injury of trunk, without mention of infection|Other and unspecified superficial injury of trunk, without mention of infection
C0840764|T037|AB|911.8|ICD9CM|Superfic inj trunk NEC|Superfic inj trunk NEC
C0160839|T037|PT|911.9|ICD9CM|Other and unspecified superficial injury of trunk, infected|Other and unspecified superficial injury of trunk, infected
C0160839|T037|AB|911.9|ICD9CM|Superf inj trnk NEC-inf|Superf inj trnk NEC-inf
C0160840|T037|HT|912|ICD9CM|Superficial injury of shoulder and upper arm|Superficial injury of shoulder and upper arm
C0160841|T037|PT|912.0|ICD9CM|Abrasion or friction burn of shoulder and upper arm, without mention of infection|Abrasion or friction burn of shoulder and upper arm, without mention of infection
C0160841|T037|AB|912.0|ICD9CM|Abrasion shoulder/arm|Abrasion shoulder/arm
C0160842|T037|PT|912.1|ICD9CM|Abrasion or friction burn of shoulder and upper arm, infected|Abrasion or friction burn of shoulder and upper arm, infected
C0160842|T037|AB|912.1|ICD9CM|Abrasion shldr/arm-infec|Abrasion shldr/arm-infec
C0160843|T037|PT|912.2|ICD9CM|Blister of shoulder and upper arm, without mention of infection|Blister of shoulder and upper arm, without mention of infection
C0160843|T037|AB|912.2|ICD9CM|Blister shoulder & arm|Blister shoulder & arm
C0160844|T037|PT|912.3|ICD9CM|Blister of shoulder and upper arm, infected|Blister of shoulder and upper arm, infected
C0160844|T037|AB|912.3|ICD9CM|Blister shoulder/arm-inf|Blister shoulder/arm-inf
C0160845|T037|AB|912.4|ICD9CM|Insect bite shoulder/arm|Insect bite shoulder/arm
C0160845|T037|PT|912.4|ICD9CM|Insect bite, nonvenomous of shoulder and upper arm, without mention of infection|Insect bite, nonvenomous of shoulder and upper arm, without mention of infection
C0160846|T037|AB|912.5|ICD9CM|Insect bite shld/arm-inf|Insect bite shld/arm-inf
C0160846|T037|PT|912.5|ICD9CM|Insect bite, nonvenomous of shoulder and upper arm, infected|Insect bite, nonvenomous of shoulder and upper arm, infected
C0160847|T037|AB|912.6|ICD9CM|Foreign body shouldr/arm|Foreign body shouldr/arm
C0160848|T037|AB|912.7|ICD9CM|FB shoulder/arm-infect|FB shoulder/arm-infect
C0160848|T037|PT|912.7|ICD9CM|Superficial foreign body (splinter) of shoulder and upper arm, without major open wound, infected|Superficial foreign body (splinter) of shoulder and upper arm, without major open wound, infected
C0478269|T037|PT|912.8|ICD9CM|Other and unspecified superficial injury of shoulder and upper arm, without mention of infection|Other and unspecified superficial injury of shoulder and upper arm, without mention of infection
C0478269|T037|AB|912.8|ICD9CM|Superf inj shldr/arm NEC|Superf inj shldr/arm NEC
C0160850|T037|PT|912.9|ICD9CM|Other and unspecified superficial injury of shoulder and upper arm, infected|Other and unspecified superficial injury of shoulder and upper arm, infected
C0160850|T037|AB|912.9|ICD9CM|Superf inj shldr NEC-inf|Superf inj shldr NEC-inf
C0160851|T037|HT|913|ICD9CM|Superficial injury of elbow, forearm, and wrist|Superficial injury of elbow, forearm, and wrist
C0160852|T037|AB|913.0|ICD9CM|Abrasion forearm|Abrasion forearm
C0160852|T037|PT|913.0|ICD9CM|Abrasion or friction burn of elbow, forearm, and wrist, without mention of infection|Abrasion or friction burn of elbow, forearm, and wrist, without mention of infection
C0160853|T037|AB|913.1|ICD9CM|Abrasion forearm-infect|Abrasion forearm-infect
C0160853|T037|PT|913.1|ICD9CM|Abrasion or friction burn of elbow, forearm, and wrist, infected|Abrasion or friction burn of elbow, forearm, and wrist, infected
C0160854|T037|AB|913.2|ICD9CM|Blister forearm|Blister forearm
C0160854|T037|PT|913.2|ICD9CM|Blister of elbow, forearm, and wrist, without mention of infection|Blister of elbow, forearm, and wrist, without mention of infection
C0160855|T037|AB|913.3|ICD9CM|Blister forearm-infected|Blister forearm-infected
C0160855|T037|PT|913.3|ICD9CM|Blister of elbow, forearm, and wrist, infected|Blister of elbow, forearm, and wrist, infected
C0160856|T037|AB|913.4|ICD9CM|Insect bite forearm|Insect bite forearm
C0160856|T037|PT|913.4|ICD9CM|Insect bite, nonvenomous of elbow, forearm, and wrist, without mention of infection|Insect bite, nonvenomous of elbow, forearm, and wrist, without mention of infection
C0160857|T037|AB|913.5|ICD9CM|Insect bite forearm-inf|Insect bite forearm-inf
C0160857|T037|PT|913.5|ICD9CM|Insect bite, nonvenomous, of elbow, forearm, and wrist, infected|Insect bite, nonvenomous, of elbow, forearm, and wrist, infected
C0160858|T037|AB|913.6|ICD9CM|Foreign body forearm|Foreign body forearm
C0160859|T037|AB|913.7|ICD9CM|Foreign body forearm-inf|Foreign body forearm-inf
C0160859|T037|PT|913.7|ICD9CM|Superficial foreign body (splinter) of elbow, forearm, and wrist, without major open wound, infected|Superficial foreign body (splinter) of elbow, forearm, and wrist, without major open wound, infected
C0160860|T037|PT|913.8|ICD9CM|Other and unspecified superficial injury of elbow, forearm, and wrist, without mention of infection|Other and unspecified superficial injury of elbow, forearm, and wrist, without mention of infection
C0160860|T037|AB|913.8|ICD9CM|Superf inj forearm NEC|Superf inj forearm NEC
C0160861|T037|PT|913.9|ICD9CM|Other and unspecified superficial injury of elbow, forearm, and wrist, infected|Other and unspecified superficial injury of elbow, forearm, and wrist, infected
C0160861|T037|AB|913.9|ICD9CM|Suprf inj forarm NEC-inf|Suprf inj forarm NEC-inf
C0432721|T037|HT|914|ICD9CM|Superficial injury of hand(s) except finger(s) alone|Superficial injury of hand(s) except finger(s) alone
C0160863|T037|AB|914.0|ICD9CM|Abrasion hand|Abrasion hand
C0160863|T037|PT|914.0|ICD9CM|Abrasion or friction burn of hand(s) except finger(s) alone, without mention of infection|Abrasion or friction burn of hand(s) except finger(s) alone, without mention of infection
C0160864|T037|AB|914.1|ICD9CM|Abrasion hand-infected|Abrasion hand-infected
C0160864|T037|PT|914.1|ICD9CM|Abrasion or friction burn of hand(s) except finger(s) alone, infected|Abrasion or friction burn of hand(s) except finger(s) alone, infected
C0160865|T037|AB|914.2|ICD9CM|Blister hand|Blister hand
C0160865|T037|PT|914.2|ICD9CM|Blister of hand(s) except finger(s) alone, without mention of infection|Blister of hand(s) except finger(s) alone, without mention of infection
C0160866|T037|AB|914.3|ICD9CM|Blister hand-infected|Blister hand-infected
C0160866|T037|PT|914.3|ICD9CM|Blister of hand(s) except finger(s) alone, infected|Blister of hand(s) except finger(s) alone, infected
C0160867|T037|AB|914.4|ICD9CM|Insect bite hand|Insect bite hand
C0160867|T037|PT|914.4|ICD9CM|Insect bite, nonvenomous, of hand(s) except finger(s) alone, without mention of infection|Insect bite, nonvenomous, of hand(s) except finger(s) alone, without mention of infection
C0160868|T037|AB|914.5|ICD9CM|Insect bite hand-infect|Insect bite hand-infect
C0160868|T037|PT|914.5|ICD9CM|Insect bite, nonvenomous, of hand(s) except finger(s) alone, infected|Insect bite, nonvenomous, of hand(s) except finger(s) alone, infected
C0160869|T037|AB|914.6|ICD9CM|Foreign body hand|Foreign body hand
C0160870|T037|AB|914.7|ICD9CM|Foreign body hand-infect|Foreign body hand-infect
C0160871|T037|AB|914.8|ICD9CM|Superficial inj hand NEC|Superficial inj hand NEC
C0160872|T037|PT|914.9|ICD9CM|Other and unspecified superficial injury of hand(s) except finger(s) alone, infected|Other and unspecified superficial injury of hand(s) except finger(s) alone, infected
C0160872|T037|AB|914.9|ICD9CM|Superf inj hand NEC-inf|Superf inj hand NEC-inf
C0558421|T037|HT|915|ICD9CM|Superficial injury of finger(s)|Superficial injury of finger(s)
C0273867|T037|AB|915.0|ICD9CM|Abrasion finger|Abrasion finger
C0273867|T037|PT|915.0|ICD9CM|Abrasion or friction burn of finger(s), without mention of infection|Abrasion or friction burn of finger(s), without mention of infection
C0160875|T037|AB|915.1|ICD9CM|Abrasion finger-infected|Abrasion finger-infected
C0160875|T037|PT|915.1|ICD9CM|Abrasion or friction burn of finger(s), infected|Abrasion or friction burn of finger(s), infected
C0160876|T037|AB|915.2|ICD9CM|Blister finger|Blister finger
C0160876|T037|PT|915.2|ICD9CM|Blister of finger(s), without mention of infection|Blister of finger(s), without mention of infection
C0160877|T037|AB|915.3|ICD9CM|Blister finger-infected|Blister finger-infected
C0160877|T037|PT|915.3|ICD9CM|Blister of finger(s), infected|Blister of finger(s), infected
C0273869|T037|AB|915.4|ICD9CM|Insect bite finger|Insect bite finger
C0273869|T037|PT|915.4|ICD9CM|Insect bite, nonvenomous, of finger(s), without mention of infection|Insect bite, nonvenomous, of finger(s), without mention of infection
C0160879|T037|AB|915.5|ICD9CM|Insect bite finger-infec|Insect bite finger-infec
C0160879|T037|PT|915.5|ICD9CM|Insect bite, nonvenomous of finger(s), infected|Insect bite, nonvenomous of finger(s), infected
C0160880|T037|AB|915.6|ICD9CM|Foreign body finger|Foreign body finger
C0160881|T037|AB|915.7|ICD9CM|Foreign body finger-inf|Foreign body finger-inf
C0160881|T037|PT|915.7|ICD9CM|Superficial foreign body (splinter) of finger(s), without major open wound, infected|Superficial foreign body (splinter) of finger(s), without major open wound, infected
C0160882|T037|PT|915.8|ICD9CM|Other and unspecified superficial injury of fingers without mention of infection|Other and unspecified superficial injury of fingers without mention of infection
C0160882|T037|AB|915.8|ICD9CM|Superfic inj finger-NEC|Superfic inj finger-NEC
C0160883|T037|PT|915.9|ICD9CM|Other and unspecified superficial injury of fingers, infected|Other and unspecified superficial injury of fingers, infected
C0160883|T037|AB|915.9|ICD9CM|Suprf inj finger NEC-inf|Suprf inj finger NEC-inf
C0160884|T037|HT|916|ICD9CM|Superficial injury of hip, thigh, leg, and ankle|Superficial injury of hip, thigh, leg, and ankle
C0160885|T037|AB|916.0|ICD9CM|Abrasion hip & leg|Abrasion hip & leg
C0160885|T037|PT|916.0|ICD9CM|Abrasion or friction burn of hip, thigh, leg, and ankle, without mention of infection|Abrasion or friction burn of hip, thigh, leg, and ankle, without mention of infection
C0160886|T037|AB|916.1|ICD9CM|Abrasion hip/leg-infect|Abrasion hip/leg-infect
C0160886|T037|PT|916.1|ICD9CM|Abrasion or friction burn of hip, thigh, leg, and ankle, infected|Abrasion or friction burn of hip, thigh, leg, and ankle, infected
C0160887|T037|AB|916.2|ICD9CM|Blister hip & leg|Blister hip & leg
C0160887|T037|PT|916.2|ICD9CM|Blister of hip, thigh, leg, and ankle, without mention of infection|Blister of hip, thigh, leg, and ankle, without mention of infection
C0160888|T037|AB|916.3|ICD9CM|Blister hip & leg-infect|Blister hip & leg-infect
C0160888|T037|PT|916.3|ICD9CM|Blister of hip, thigh, leg, and ankle, infected|Blister of hip, thigh, leg, and ankle, infected
C0160889|T037|AB|916.4|ICD9CM|Insect bite hip & leg|Insect bite hip & leg
C0160889|T037|PT|916.4|ICD9CM|Insect bite, nonvenomous, of hip, thigh, leg, and ankle, without mention of infection|Insect bite, nonvenomous, of hip, thigh, leg, and ankle, without mention of infection
C0160890|T037|AB|916.5|ICD9CM|Insect bite hip/leg-inf|Insect bite hip/leg-inf
C0160890|T037|PT|916.5|ICD9CM|Insect bite, nonvenomous of hip, thigh, leg, and ankle, infected|Insect bite, nonvenomous of hip, thigh, leg, and ankle, infected
C0160891|T037|AB|916.6|ICD9CM|Foreign body hip/leg|Foreign body hip/leg
C0160892|T037|AB|916.7|ICD9CM|Foreign bdy hip/leg-inf|Foreign bdy hip/leg-inf
C0160893|T037|PT|916.8|ICD9CM|Other and unspecified superficial injury of hip, thigh, leg, and ankle, without mention of infection|Other and unspecified superficial injury of hip, thigh, leg, and ankle, without mention of infection
C0160893|T037|AB|916.8|ICD9CM|Superfic inj hip/leg NEC|Superfic inj hip/leg NEC
C0160894|T037|PT|916.9|ICD9CM|Other and unspecified superficial injury of hip, thigh, leg, and ankle, infected|Other and unspecified superficial injury of hip, thigh, leg, and ankle, infected
C0160894|T037|AB|916.9|ICD9CM|Superf inj leg NEC-infec|Superf inj leg NEC-infec
C0160895|T037|HT|917|ICD9CM|Superficial injury of foot and toe(s)|Superficial injury of foot and toe(s)
C0432869|T037|AB|917.0|ICD9CM|Abrasion foot & toe|Abrasion foot & toe
C0432869|T037|PT|917.0|ICD9CM|Abrasion or friction burn of foot and toe(s), without mention of infection|Abrasion or friction burn of foot and toe(s), without mention of infection
C0432873|T037|AB|917.1|ICD9CM|Abrasion foot/toe-infec|Abrasion foot/toe-infec
C0432873|T037|PT|917.1|ICD9CM|Abrasion or friction burn of foot and toe(s), infected|Abrasion or friction burn of foot and toe(s), infected
C0432918|T037|AB|917.2|ICD9CM|Blister foot & toe|Blister foot & toe
C0432918|T037|PT|917.2|ICD9CM|Blister of foot and toe(s), without mention of infection|Blister of foot and toe(s), without mention of infection
C0432922|T037|AB|917.3|ICD9CM|Blister foot & toe-infec|Blister foot & toe-infec
C0432922|T037|PT|917.3|ICD9CM|Blister of foot and toe(s), infected|Blister of foot and toe(s), infected
C0433039|T037|AB|917.4|ICD9CM|Insect bite foot/toe|Insect bite foot/toe
C0433039|T037|PT|917.4|ICD9CM|Insect bite, nonvenomous, of foot and toe(s), without mention of infection|Insect bite, nonvenomous, of foot and toe(s), without mention of infection
C0433050|T037|AB|917.5|ICD9CM|Insect bite foot/toe-inf|Insect bite foot/toe-inf
C0433050|T037|PT|917.5|ICD9CM|Insect bite, nonvenomous, of foot and toe(s), infected|Insect bite, nonvenomous, of foot and toe(s), infected
C0160902|T037|AB|917.6|ICD9CM|Foreign body foot & toe|Foreign body foot & toe
C0160903|T037|AB|917.7|ICD9CM|Foreign bdy foot/toe-inf|Foreign bdy foot/toe-inf
C0160903|T037|PT|917.7|ICD9CM|Superficial foreign body (splinter) of foot and toe(s), without major open wound, infected|Superficial foreign body (splinter) of foot and toe(s), without major open wound, infected
C0160904|T037|PT|917.8|ICD9CM|Other and unspecified superficial injury of foot and toes, without mention of infection|Other and unspecified superficial injury of foot and toes, without mention of infection
C0160904|T037|AB|917.8|ICD9CM|Superf inj foot/toe NEC|Superf inj foot/toe NEC
C0160905|T037|PT|917.9|ICD9CM|Other and unspecified superficial injury of foot and toes, infected|Other and unspecified superficial injury of foot and toes, infected
C0160905|T037|AB|917.9|ICD9CM|Superf inj foot NEC-inf|Superf inj foot NEC-inf
C0160906|T037|HT|918|ICD9CM|Superficial injury of eye and adnexa|Superficial injury of eye and adnexa
C0160907|T037|AB|918.0|ICD9CM|Superfic inj periocular|Superfic inj periocular
C0160907|T037|PT|918.0|ICD9CM|Superficial injury of eyelids and periocular area|Superficial injury of eyelids and periocular area
C0038824|T037|AB|918.1|ICD9CM|Superficial inj cornea|Superficial inj cornea
C0038824|T037|PT|918.1|ICD9CM|Superficial injury of cornea|Superficial injury of cornea
C0160908|T037|AB|918.2|ICD9CM|Superfic inj conjunctiva|Superfic inj conjunctiva
C0160908|T037|PT|918.2|ICD9CM|Superficial injury of conjunctiva|Superficial injury of conjunctiva
C0160909|T037|PT|918.9|ICD9CM|Other and unspecified superficial injuries of eye|Other and unspecified superficial injuries of eye
C0160909|T037|AB|918.9|ICD9CM|Superficial inj eye NEC|Superficial inj eye NEC
C0160910|T037|HT|919|ICD9CM|Superficial injury of other, multiple, and unspecified sites|Superficial injury of other, multiple, and unspecified sites
C0000827|T037|AB|919.0|ICD9CM|Abrasion NEC|Abrasion NEC
C0000827|T037|PT|919.0|ICD9CM|Abrasion or friction burn of other, multiple, and unspecified sites, without mention of infection|Abrasion or friction burn of other, multiple, and unspecified sites, without mention of infection
C0160911|T037|AB|919.1|ICD9CM|Abrasion NEC-infected|Abrasion NEC-infected
C0160911|T037|PT|919.1|ICD9CM|Abrasion or friction burn of other, multiple, and unspecified sites, infected|Abrasion or friction burn of other, multiple, and unspecified sites, infected
C0005761|T037|AB|919.2|ICD9CM|Blister NEC|Blister NEC
C0005761|T037|PT|919.2|ICD9CM|Blister of other, multiple, and unspecified sites, without mention of infection|Blister of other, multiple, and unspecified sites, without mention of infection
C0160912|T037|AB|919.3|ICD9CM|Blister NEC-infected|Blister NEC-infected
C0160912|T037|PT|919.3|ICD9CM|Blister of other, multiple, and unspecified sites, infected|Blister of other, multiple, and unspecified sites, infected
C0021567|T037|AB|919.4|ICD9CM|Insect bite NEC|Insect bite NEC
C0021567|T037|PT|919.4|ICD9CM|Insect bite, nonvenomous, of other, multiple, and unspecified sites, without mention of infection|Insect bite, nonvenomous, of other, multiple, and unspecified sites, without mention of infection
C0160913|T037|AB|919.5|ICD9CM|Insect bite NEC-infected|Insect bite NEC-infected
C0160913|T037|PT|919.5|ICD9CM|Insect bite, nonvenomous, of other, multiple, and unspecified sites, infected|Insect bite, nonvenomous, of other, multiple, and unspecified sites, infected
C0160914|T037|AB|919.6|ICD9CM|Superfic foreign bdy NEC|Superfic foreign bdy NEC
C0160915|T037|AB|919.7|ICD9CM|Superficial FB NEC-infec|Superficial FB NEC-infec
C0160916|T037|AB|919.8|ICD9CM|Superficial injury NEC|Superficial injury NEC
C0160917|T037|PT|919.9|ICD9CM|Other and unspecified superficial injury of other, multiple, and unspecified sites, infected|Other and unspecified superficial injury of other, multiple, and unspecified sites, infected
C0160917|T037|AB|919.9|ICD9CM|Superfic inj NEC-infect|Superfic inj NEC-infect
C0160918|T037|AB|920|ICD9CM|Contusion face/scalp/nck|Contusion face/scalp/nck
C0160918|T037|PT|920|ICD9CM|Contusion of face, scalp, and neck except eye(s)|Contusion of face, scalp, and neck except eye(s)
C0178327|T037|HT|920-924.99|ICD9CM|CONTUSION WITH INTACT SKIN SURFACE|CONTUSION WITH INTACT SKIN SURFACE
C0160919|T037|HT|921|ICD9CM|Contusion of eye and adnexa|Contusion of eye and adnexa
C1442861|T033|AB|921.0|ICD9CM|Black eye NOS|Black eye NOS
C1442861|T033|PT|921.0|ICD9CM|Black eye, not otherwise specified|Black eye, not otherwise specified
C0160920|T037|PT|921.1|ICD9CM|Contusion of eyelids and periocular area|Contusion of eyelids and periocular area
C0160920|T037|AB|921.1|ICD9CM|Contusion periocular|Contusion periocular
C0160921|T037|PT|921.2|ICD9CM|Contusion of orbital tissues|Contusion of orbital tissues
C0160921|T037|AB|921.2|ICD9CM|Contusion orbital tissue|Contusion orbital tissue
C2939443|T037|AB|921.3|ICD9CM|Contusion of eyeball|Contusion of eyeball
C2939443|T037|PT|921.3|ICD9CM|Contusion of eyeball|Contusion of eyeball
C0438624|T037|AB|921.9|ICD9CM|Contusion of eye NOS|Contusion of eye NOS
C0438624|T037|PT|921.9|ICD9CM|Unspecified contusion of eye|Unspecified contusion of eye
C0160923|T037|HT|922|ICD9CM|Contusion of trunk|Contusion of trunk
C0160924|T037|AB|922.0|ICD9CM|Contusion of breast|Contusion of breast
C0160924|T037|PT|922.0|ICD9CM|Contusion of breast|Contusion of breast
C0160925|T037|AB|922.1|ICD9CM|Contusion of chest wall|Contusion of chest wall
C0160925|T037|PT|922.1|ICD9CM|Contusion of chest wall|Contusion of chest wall
C0160926|T037|AB|922.2|ICD9CM|Contusion abdominal wall|Contusion abdominal wall
C0160926|T037|PT|922.2|ICD9CM|Contusion of abdominal wall|Contusion of abdominal wall
C0160927|T037|HT|922.3|ICD9CM|Contusion of back|Contusion of back
C0160927|T037|AB|922.31|ICD9CM|Back contusion|Back contusion
C0160927|T037|PT|922.31|ICD9CM|Contusion of back|Contusion of back
C0274220|T037|AB|922.32|ICD9CM|Buttock contusion|Buttock contusion
C0274220|T037|PT|922.32|ICD9CM|Contusion of buttock|Contusion of buttock
C0274221|T037|PT|922.33|ICD9CM|Contusion of interscapular region|Contusion of interscapular region
C0274221|T037|AB|922.33|ICD9CM|Interscplr reg contusion|Interscplr reg contusion
C0160928|T037|AB|922.4|ICD9CM|Contusion genital organs|Contusion genital organs
C0160928|T037|PT|922.4|ICD9CM|Contusion of genital organs|Contusion of genital organs
C0160929|T037|PT|922.8|ICD9CM|Contusion of multiple sites of trunk|Contusion of multiple sites of trunk
C0160929|T037|AB|922.8|ICD9CM|Multiple contusion trunk|Multiple contusion trunk
C0160923|T037|PT|922.9|ICD9CM|Contusion of unspecified part of trunk|Contusion of unspecified part of trunk
C0160923|T037|AB|922.9|ICD9CM|Contusion trunk NOS|Contusion trunk NOS
C0160931|T037|HT|923|ICD9CM|Contusion of upper limb|Contusion of upper limb
C0160932|T037|HT|923.0|ICD9CM|Contusion of shoulder and upper arm|Contusion of shoulder and upper arm
C0160933|T037|PT|923.00|ICD9CM|Contusion of shoulder region|Contusion of shoulder region
C0160933|T037|AB|923.00|ICD9CM|Contusion shoulder reg|Contusion shoulder reg
C0160934|T037|PT|923.01|ICD9CM|Contusion of scapular region|Contusion of scapular region
C0160934|T037|AB|923.01|ICD9CM|Contusion scapul region|Contusion scapul region
C0160935|T037|AB|923.02|ICD9CM|Contusion axillary reg|Contusion axillary reg
C0160935|T037|PT|923.02|ICD9CM|Contusion of axillary region|Contusion of axillary region
C0160936|T037|AB|923.03|ICD9CM|Contusion of upper arm|Contusion of upper arm
C0160936|T037|PT|923.03|ICD9CM|Contusion of upper arm|Contusion of upper arm
C0160937|T037|PT|923.09|ICD9CM|Contusion of multiple sites of shoulder and upper arm|Contusion of multiple sites of shoulder and upper arm
C0160937|T037|AB|923.09|ICD9CM|Contusion shoulder & arm|Contusion shoulder & arm
C0160938|T037|HT|923.1|ICD9CM|Contusion of elbow and forearm|Contusion of elbow and forearm
C0432762|T037|AB|923.10|ICD9CM|Contusion of forearm|Contusion of forearm
C0432762|T037|PT|923.10|ICD9CM|Contusion of forearm|Contusion of forearm
C0432763|T037|AB|923.11|ICD9CM|Contusion of elbow|Contusion of elbow
C0432763|T037|PT|923.11|ICD9CM|Contusion of elbow|Contusion of elbow
C0160941|T037|HT|923.2|ICD9CM|Contusion of wrist and hand(s), except finger(s) alone|Contusion of wrist and hand(s), except finger(s) alone
C0432769|T037|AB|923.20|ICD9CM|Contusion of hand(s)|Contusion of hand(s)
C0432769|T037|PT|923.20|ICD9CM|Contusion of hand(s)|Contusion of hand(s)
C0160943|T037|AB|923.21|ICD9CM|Contusion of wrist|Contusion of wrist
C0160943|T037|PT|923.21|ICD9CM|Contusion of wrist|Contusion of wrist
C0432773|T037|AB|923.3|ICD9CM|Contusion of finger|Contusion of finger
C0432773|T037|PT|923.3|ICD9CM|Contusion of finger|Contusion of finger
C0160945|T037|PT|923.8|ICD9CM|Contusion of multiple sites of upper limb|Contusion of multiple sites of upper limb
C0160945|T037|AB|923.8|ICD9CM|Multiple contusion arm|Multiple contusion arm
C0160931|T037|PT|923.9|ICD9CM|Contusion of unspecified part of upper limb|Contusion of unspecified part of upper limb
C0160931|T037|AB|923.9|ICD9CM|Contusion upper limb NOS|Contusion upper limb NOS
C0160947|T037|HT|924|ICD9CM|Contusion of lower limb and of other and unspecified sites|Contusion of lower limb and of other and unspecified sites
C0160948|T037|HT|924.0|ICD9CM|Contusion of hip and thigh|Contusion of hip and thigh
C0160949|T037|AB|924.00|ICD9CM|Contusion of thigh|Contusion of thigh
C0160949|T037|PT|924.00|ICD9CM|Contusion of thigh|Contusion of thigh
C0160950|T037|AB|924.01|ICD9CM|Contusion of hip|Contusion of hip
C0160950|T037|PT|924.01|ICD9CM|Contusion of hip|Contusion of hip
C0160951|T037|HT|924.1|ICD9CM|Contusion of knee and lower leg|Contusion of knee and lower leg
C0160952|T037|AB|924.10|ICD9CM|Contusion of lower leg|Contusion of lower leg
C0160952|T037|PT|924.10|ICD9CM|Contusion of lower leg|Contusion of lower leg
C0160953|T037|AB|924.11|ICD9CM|Contusion of knee|Contusion of knee
C0160953|T037|PT|924.11|ICD9CM|Contusion of knee|Contusion of knee
C0274237|T037|HT|924.2|ICD9CM|Contusion of ankle and foot, excluding toe(s)|Contusion of ankle and foot, excluding toe(s)
C0160955|T033|AB|924.20|ICD9CM|Contusion of foot|Contusion of foot
C0160955|T033|PT|924.20|ICD9CM|Contusion of foot|Contusion of foot
C0160956|T037|AB|924.21|ICD9CM|Contusion of ankle|Contusion of ankle
C0160956|T037|PT|924.21|ICD9CM|Contusion of ankle|Contusion of ankle
C0160957|T037|AB|924.3|ICD9CM|Contusion of toe|Contusion of toe
C0160957|T037|PT|924.3|ICD9CM|Contusion of toe|Contusion of toe
C0160958|T037|PT|924.4|ICD9CM|Contusion of multiple sites of lower limb|Contusion of multiple sites of lower limb
C0160958|T037|AB|924.4|ICD9CM|Multiple contusion leg|Multiple contusion leg
C0274236|T037|AB|924.5|ICD9CM|Contusion leg NOS|Contusion leg NOS
C0274236|T037|PT|924.5|ICD9CM|Contusion of unspecified part of lower limb|Contusion of unspecified part of lower limb
C0160960|T037|PT|924.8|ICD9CM|Contusion of multiple sites, not elsewhere classified|Contusion of multiple sites, not elsewhere classified
C0160960|T037|AB|924.8|ICD9CM|Multiple contusions NEC|Multiple contusions NEC
C0009938|T037|AB|924.9|ICD9CM|Contusion NOS|Contusion NOS
C0009938|T037|PT|924.9|ICD9CM|Contusion of unspecified site|Contusion of unspecified site
C0160961|T037|HT|925|ICD9CM|Crushing injury of face, scalp, and neck|Crushing injury of face, scalp, and neck
C0332679|T037|HT|925-929.99|ICD9CM|CRUSHING INJURY|CRUSHING INJURY
C0375669|T037|AB|925.1|ICD9CM|Crush inj face scalp|Crush inj face scalp
C0375669|T037|PT|925.1|ICD9CM|Crushing injury of face and scalp|Crushing injury of face and scalp
C0273433|T037|AB|925.2|ICD9CM|Crush inj neck|Crush inj neck
C0273433|T037|PT|925.2|ICD9CM|Crushing injury of neck|Crushing injury of neck
C0160962|T037|HT|926|ICD9CM|Crushing injury of trunk|Crushing injury of trunk
C0160963|T037|AB|926.0|ICD9CM|Crush inj ext genitalia|Crush inj ext genitalia
C0160963|T037|PT|926.0|ICD9CM|Crushing injury of external genitalia|Crushing injury of external genitalia
C0160964|T037|HT|926.1|ICD9CM|Crushing injury of other specified sites of trunk|Crushing injury of other specified sites of trunk
C0160965|T037|AB|926.11|ICD9CM|Crushing injury back|Crushing injury back
C0160965|T037|PT|926.11|ICD9CM|Crushing injury of back|Crushing injury of back
C0160966|T037|AB|926.12|ICD9CM|Crushing injury buttock|Crushing injury buttock
C0160966|T037|PT|926.12|ICD9CM|Crushing injury of buttock|Crushing injury of buttock
C0160964|T037|AB|926.19|ICD9CM|Crushing inj trunk NEC|Crushing inj trunk NEC
C0160964|T037|PT|926.19|ICD9CM|Crushing injury of other specified sites of trunk|Crushing injury of other specified sites of trunk
C0160967|T037|PT|926.8|ICD9CM|Crushing injury of multiple sites of trunk|Crushing injury of multiple sites of trunk
C0160967|T037|AB|926.8|ICD9CM|Mult crushing inj trunk|Mult crushing inj trunk
C0160962|T037|AB|926.9|ICD9CM|Crushing inj trunk NOS|Crushing inj trunk NOS
C0160962|T037|PT|926.9|ICD9CM|Crushing injury of unspecified site of trunk|Crushing injury of unspecified site of trunk
C0160969|T037|HT|927|ICD9CM|Crushing injury of upper limb|Crushing injury of upper limb
C0160970|T037|HT|927.0|ICD9CM|Crushing injury of shoulder and upper arm|Crushing injury of shoulder and upper arm
C0160971|T037|AB|927.00|ICD9CM|Crush inj shoulder reg|Crush inj shoulder reg
C0160971|T037|PT|927.00|ICD9CM|Crushing injury of shoulder region|Crushing injury of shoulder region
C0160972|T037|AB|927.01|ICD9CM|Crush inj scapul region|Crush inj scapul region
C0160972|T037|PT|927.01|ICD9CM|Crushing injury of scapular region|Crushing injury of scapular region
C0160973|T037|AB|927.02|ICD9CM|Crush inj axillary reg|Crush inj axillary reg
C0160973|T037|PT|927.02|ICD9CM|Crushing injury of axillary region|Crushing injury of axillary region
C0160974|T037|AB|927.03|ICD9CM|Crushing inj upper arm|Crushing inj upper arm
C0160974|T037|PT|927.03|ICD9CM|Crushing injury of upper arm|Crushing injury of upper arm
C0160975|T037|AB|927.09|ICD9CM|Crush inj shoulder & arm|Crush inj shoulder & arm
C0160975|T037|PT|927.09|ICD9CM|Crushing injury of multiple sites of upper arm|Crushing injury of multiple sites of upper arm
C0160976|T037|HT|927.1|ICD9CM|Crushing injury of elbow and forearm|Crushing injury of elbow and forearm
C0160977|T037|AB|927.10|ICD9CM|Crushing injury forearm|Crushing injury forearm
C0160977|T037|PT|927.10|ICD9CM|Crushing injury of forearm|Crushing injury of forearm
C0160978|T037|AB|927.11|ICD9CM|Crushing injury elbow|Crushing injury elbow
C0160978|T037|PT|927.11|ICD9CM|Crushing injury of elbow|Crushing injury of elbow
C0160979|T037|HT|927.2|ICD9CM|Crushing injury of wrist and hand(s), except finger(s) alone|Crushing injury of wrist and hand(s), except finger(s) alone
C0273444|T037|AB|927.20|ICD9CM|Crushing injury of hand|Crushing injury of hand
C0273444|T037|PT|927.20|ICD9CM|Crushing injury of hand(s)|Crushing injury of hand(s)
C0160981|T037|AB|927.21|ICD9CM|Crushing injury of wrist|Crushing injury of wrist
C0160981|T037|PT|927.21|ICD9CM|Crushing injury of wrist|Crushing injury of wrist
C0273445|T037|AB|927.3|ICD9CM|Crushing injury finger|Crushing injury finger
C0273445|T037|PT|927.3|ICD9CM|Crushing injury of finger(s)|Crushing injury of finger(s)
C0160983|T037|PT|927.8|ICD9CM|Crushing injury of multiple sites of upper limb|Crushing injury of multiple sites of upper limb
C0160983|T037|AB|927.8|ICD9CM|Mult crushing injury arm|Mult crushing injury arm
C0160969|T037|AB|927.9|ICD9CM|Crushing injury arm NOS|Crushing injury arm NOS
C0160969|T037|PT|927.9|ICD9CM|Crushing injury of unspecified site of upper limb|Crushing injury of unspecified site of upper limb
C0160985|T037|HT|928|ICD9CM|Crushing injury of lower limb|Crushing injury of lower limb
C0160986|T037|HT|928.0|ICD9CM|Crushing injury of hip and thigh|Crushing injury of hip and thigh
C0160987|T037|PT|928.00|ICD9CM|Crushing injury of thigh|Crushing injury of thigh
C0160987|T037|AB|928.00|ICD9CM|Crushing injury thigh|Crushing injury thigh
C0160988|T037|AB|928.01|ICD9CM|Crushing injury hip|Crushing injury hip
C0160988|T037|PT|928.01|ICD9CM|Crushing injury of hip|Crushing injury of hip
C0160989|T037|HT|928.1|ICD9CM|Crushing injury of knee and lower leg|Crushing injury of knee and lower leg
C0160990|T037|AB|928.10|ICD9CM|Crushing inj lower leg|Crushing inj lower leg
C0160990|T037|PT|928.10|ICD9CM|Crushing injury of lower leg|Crushing injury of lower leg
C0160991|T037|AB|928.11|ICD9CM|Crushing injury knee|Crushing injury knee
C0160991|T037|PT|928.11|ICD9CM|Crushing injury of knee|Crushing injury of knee
C0160992|T037|HT|928.2|ICD9CM|Crushing injury of ankle and foot, excluding toe(s) alone|Crushing injury of ankle and foot, excluding toe(s) alone
C0160993|T037|AB|928.20|ICD9CM|Crushing injury foot|Crushing injury foot
C0160993|T037|PT|928.20|ICD9CM|Crushing injury of foot|Crushing injury of foot
C0160994|T037|AB|928.21|ICD9CM|Crushing injury ankle|Crushing injury ankle
C0160994|T037|PT|928.21|ICD9CM|Crushing injury of ankle|Crushing injury of ankle
C0273448|T037|PT|928.3|ICD9CM|Crushing injury of toe(s)|Crushing injury of toe(s)
C0273448|T037|AB|928.3|ICD9CM|Crushing injury toe|Crushing injury toe
C0160996|T037|PT|928.8|ICD9CM|Crushing injury of multiple sites of lower limb|Crushing injury of multiple sites of lower limb
C0160996|T037|AB|928.8|ICD9CM|Mult crushing injury leg|Mult crushing injury leg
C0160985|T037|AB|928.9|ICD9CM|Crushing injury leg NOS|Crushing injury leg NOS
C0160985|T037|PT|928.9|ICD9CM|Crushing injury of unspecified site of lower limb|Crushing injury of unspecified site of lower limb
C0451984|T037|HT|929|ICD9CM|Crushing injury of multiple and unspecified sites|Crushing injury of multiple and unspecified sites
C0868762|T037|AB|929.0|ICD9CM|Crush inj mult site NEC|Crush inj mult site NEC
C0868762|T037|PT|929.0|ICD9CM|Crushing injury of multiple sites, not elsewhere classified|Crushing injury of multiple sites, not elsewhere classified
C0332679|T037|AB|929.9|ICD9CM|Crushing injury NOS|Crushing injury NOS
C0332679|T037|PT|929.9|ICD9CM|Crushing injury of unspecified site|Crushing injury of unspecified site
C0161001|T037|HT|930|ICD9CM|Foreign body on external eye|Foreign body on external eye
C0178329|T037|HT|930-939.99|ICD9CM|EFFECTS OF FOREIGN BODY ENTERING THROUGH ORIFICE|EFFECTS OF FOREIGN BODY ENTERING THROUGH ORIFICE
C0161002|T037|AB|930.0|ICD9CM|Corneal foreign body|Corneal foreign body
C0161002|T037|PT|930.0|ICD9CM|Corneal foreign body|Corneal foreign body
C0161003|T037|AB|930.1|ICD9CM|FB in conjunctival sac|FB in conjunctival sac
C0161003|T037|PT|930.1|ICD9CM|Foreign body in conjunctival sac|Foreign body in conjunctival sac
C0161004|T037|AB|930.2|ICD9CM|FB in lacrimal punctum|FB in lacrimal punctum
C0161004|T037|PT|930.2|ICD9CM|Foreign body in lacrimal punctum|Foreign body in lacrimal punctum
C0161005|T037|AB|930.8|ICD9CM|Foreign bdy ext eye NEC|Foreign bdy ext eye NEC
C0161005|T037|PT|930.8|ICD9CM|Foreign body in other and combined sites on external eye|Foreign body in other and combined sites on external eye
C0161001|T037|AB|930.9|ICD9CM|Foreign bdy ext eye NOS|Foreign bdy ext eye NOS
C0161001|T037|PT|930.9|ICD9CM|Foreign body in unspecified site on external eye|Foreign body in unspecified site on external eye
C0161007|T037|AB|931|ICD9CM|Foreign body in ear|Foreign body in ear
C0161007|T037|PT|931|ICD9CM|Foreign body in ear|Foreign body in ear
C0161008|T033|AB|932|ICD9CM|Foreign body in nose|Foreign body in nose
C0161008|T033|PT|932|ICD9CM|Foreign body in nose|Foreign body in nose
C0161009|T037|HT|933|ICD9CM|Foreign body in pharynx and larynx|Foreign body in pharynx and larynx
C0161010|T037|AB|933.0|ICD9CM|Foreign body in pharynx|Foreign body in pharynx
C0161010|T037|PT|933.0|ICD9CM|Foreign body in pharynx|Foreign body in pharynx
C0161011|T037|AB|933.1|ICD9CM|Foreign body in larynx|Foreign body in larynx
C0161011|T037|PT|933.1|ICD9CM|Foreign body in larynx|Foreign body in larynx
C0686705|T037|HT|934|ICD9CM|Foreign body in trachea, bronchus, and lung|Foreign body in trachea, bronchus, and lung
C0161013|T037|AB|934.0|ICD9CM|Foreign body in trachea|Foreign body in trachea
C0161013|T037|PT|934.0|ICD9CM|Foreign body in trachea|Foreign body in trachea
C0161014|T037|AB|934.1|ICD9CM|Foreign body bronchus|Foreign body bronchus
C0161014|T037|PT|934.1|ICD9CM|Foreign body in main bronchus|Foreign body in main bronchus
C0161015|T037|AB|934.8|ICD9CM|FB trach/bronch/lung NEC|FB trach/bronch/lung NEC
C0161015|T037|PT|934.8|ICD9CM|Foreign body in other specified parts bronchus and lung|Foreign body in other specified parts bronchus and lung
C0161016|T037|AB|934.9|ICD9CM|FB respiratory tree NOS|FB respiratory tree NOS
C0161016|T037|PT|934.9|ICD9CM|Foreign body in respiratory tree, unspecified|Foreign body in respiratory tree, unspecified
C0161017|T037|HT|935|ICD9CM|Foreign body in mouth, esophagus, and stomach|Foreign body in mouth, esophagus, and stomach
C0161018|T037|AB|935.0|ICD9CM|Foreign body in mouth|Foreign body in mouth
C0161018|T037|PT|935.0|ICD9CM|Foreign body in mouth|Foreign body in mouth
C0149532|T037|AB|935.1|ICD9CM|Foreign body esophagus|Foreign body esophagus
C0149532|T037|PT|935.1|ICD9CM|Foreign body in esophagus|Foreign body in esophagus
C0161019|T037|AB|935.2|ICD9CM|Foreign body in stomach|Foreign body in stomach
C0161019|T037|PT|935.2|ICD9CM|Foreign body in stomach|Foreign body in stomach
C0161020|T033|AB|936|ICD9CM|FB in intestine & colon|FB in intestine & colon
C0161020|T033|PT|936|ICD9CM|Foreign body in intestine and colon|Foreign body in intestine and colon
C0161021|T037|AB|937|ICD9CM|Foreign body anus/rectum|Foreign body anus/rectum
C0161021|T037|PT|937|ICD9CM|Foreign body in anus and rectum|Foreign body in anus and rectum
C0016546|T037|AB|938|ICD9CM|Foreign body GI NOS|Foreign body GI NOS
C0016546|T037|PT|938|ICD9CM|Foreign body in digestive system, unspecified|Foreign body in digestive system, unspecified
C0161022|T037|HT|939|ICD9CM|Foreign body in genitourinary tract|Foreign body in genitourinary tract
C0161023|T037|AB|939.0|ICD9CM|FB bladder & urethra|FB bladder & urethra
C0161023|T037|PT|939.0|ICD9CM|Foreign body in bladder and urethra|Foreign body in bladder and urethra
C0433686|T037|PT|939.1|ICD9CM|Foreign body in uterus, any part|Foreign body in uterus, any part
C0433686|T037|AB|939.1|ICD9CM|Foreign body uterus|Foreign body uterus
C0161025|T037|AB|939.2|ICD9CM|Foreign bdy vulva/vagina|Foreign bdy vulva/vagina
C0161025|T037|PT|939.2|ICD9CM|Foreign body in vulva and vagina|Foreign body in vulva and vagina
C0161026|T037|PT|939.3|ICD9CM|Foreign body in penis|Foreign body in penis
C0161026|T037|AB|939.3|ICD9CM|Foreign body penis|Foreign body penis
C0161022|T037|AB|939.9|ICD9CM|Foreign bdy gu tract NOS|Foreign bdy gu tract NOS
C0161022|T037|PT|939.9|ICD9CM|Foreign body in unspecified site in genitourinary tract|Foreign body in unspecified site in genitourinary tract
C0273934|T037|HT|940|ICD9CM|Burn confined to eye and adnexa|Burn confined to eye and adnexa
C0006434|T037|HT|940-949.99|ICD9CM|BURNS|BURNS
C1306015|T037|PT|940.0|ICD9CM|Chemical burn of eyelids and periocular area|Chemical burn of eyelids and periocular area
C1306015|T037|AB|940.0|ICD9CM|Chemical burn periocular|Chemical burn periocular
C0161029|T037|AB|940.1|ICD9CM|Burn periocular area NEC|Burn periocular area NEC
C0161029|T037|PT|940.1|ICD9CM|Other burns of eyelids and periocular area|Other burns of eyelids and periocular area
C0161030|T037|AB|940.2|ICD9CM|Alkal burn cornea/conjun|Alkal burn cornea/conjun
C0161030|T037|PT|940.2|ICD9CM|Alkaline chemical burn of cornea and conjunctival sac|Alkaline chemical burn of cornea and conjunctival sac
C0161031|T037|AB|940.3|ICD9CM|Acid burn cornea/conjunc|Acid burn cornea/conjunc
C0161031|T037|PT|940.3|ICD9CM|Acid chemical burn of cornea and conjunctival sac|Acid chemical burn of cornea and conjunctival sac
C3665446|T037|AB|940.4|ICD9CM|Burn cornea/conjunct NEC|Burn cornea/conjunct NEC
C3665446|T037|PT|940.4|ICD9CM|Other burn of cornea and conjunctival sac|Other burn of cornea and conjunctival sac
C0161033|T037|AB|940.5|ICD9CM|Burn w eyeball destruct|Burn w eyeball destruct
C0161033|T037|PT|940.5|ICD9CM|Burn with resulting rupture and destruction of eyeball|Burn with resulting rupture and destruction of eyeball
C0273934|T037|AB|940.9|ICD9CM|Burn eye & adnexa NOS|Burn eye & adnexa NOS
C0273934|T037|PT|940.9|ICD9CM|Unspecified burn of eye and adnexa|Unspecified burn of eye and adnexa
C2004482|T037|HT|941|ICD9CM|Burn of face, head, and neck|Burn of face, head, and neck
C0496029|T037|HT|941.0|ICD9CM|Burn of face, head, and neck, unspecified degree|Burn of face, head, and neck, unspecified degree
C0273940|T037|AB|941.00|ICD9CM|Burn NOS head-unspec|Burn NOS head-unspec
C0273940|T037|PT|941.00|ICD9CM|Burn of unspecified degree of face and head, unspecified site|Burn of unspecified degree of face and head, unspecified site
C0161036|T037|AB|941.01|ICD9CM|Burn NOS ear|Burn NOS ear
C0161036|T037|PT|941.01|ICD9CM|Burn of unspecified degree of ear [any part]|Burn of unspecified degree of ear [any part]
C0006421|T037|AB|941.02|ICD9CM|Burn NOS eye|Burn NOS eye
C0006421|T037|PT|941.02|ICD9CM|Burn of unspecified degree of eye (with other parts of face, head, and neck)|Burn of unspecified degree of eye (with other parts of face, head, and neck)
C0161037|T037|AB|941.03|ICD9CM|Burn NOS lip|Burn NOS lip
C0161037|T037|PT|941.03|ICD9CM|Burn of unspecified degree of lip(s)|Burn of unspecified degree of lip(s)
C0161038|T037|AB|941.04|ICD9CM|Burn NOS chin|Burn NOS chin
C0161038|T037|PT|941.04|ICD9CM|Burn of unspecified degree of chin|Burn of unspecified degree of chin
C0869240|T037|AB|941.05|ICD9CM|Burn NOS nose|Burn NOS nose
C0869240|T037|PT|941.05|ICD9CM|Burn of unspecified degree of nose (septum)|Burn of unspecified degree of nose (septum)
C0273970|T037|AB|941.06|ICD9CM|Burn NOS scalp|Burn NOS scalp
C0273970|T037|PT|941.06|ICD9CM|Burn of unspecified degree of scalp [any part]|Burn of unspecified degree of scalp [any part]
C0161041|T037|AB|941.07|ICD9CM|Burn NOS face NEC|Burn NOS face NEC
C0161041|T037|PT|941.07|ICD9CM|Burn of unspecified degree of forehead and cheek|Burn of unspecified degree of forehead and cheek
C0273982|T037|AB|941.08|ICD9CM|Burn NOS neck|Burn NOS neck
C0273982|T037|PT|941.08|ICD9CM|Burn of unspecified degree of neck|Burn of unspecified degree of neck
C0161043|T037|AB|941.09|ICD9CM|Burn NOS head-mult|Burn NOS head-mult
C0161043|T037|PT|941.09|ICD9CM|Burn of unspecified degree of multiple sites [except with eye] of face, head, and neck|Burn of unspecified degree of multiple sites [except with eye] of face, head, and neck
C0161044|T037|HT|941.1|ICD9CM|Erythema due to burn [first degree] of face, head, and neck|Erythema due to burn [first degree] of face, head, and neck
C0273941|T037|AB|941.10|ICD9CM|1st deg burn head NOS|1st deg burn head NOS
C0273941|T037|PT|941.10|ICD9CM|Erythema [first degree] of face and head, unspecified site|Erythema [first degree] of face and head, unspecified site
C0161046|T037|AB|941.11|ICD9CM|1st deg burn ear|1st deg burn ear
C0161046|T037|PT|941.11|ICD9CM|Erythema [first degree] of ear [any part]|Erythema [first degree] of ear [any part]
C0161047|T037|AB|941.12|ICD9CM|1st deg burn eye|1st deg burn eye
C0161047|T037|PT|941.12|ICD9CM|Erythema [first degree] of eye (with other parts face, head, and neck)|Erythema [first degree] of eye (with other parts face, head, and neck)
C0161048|T037|AB|941.13|ICD9CM|1st deg burn lip|1st deg burn lip
C0161048|T037|PT|941.13|ICD9CM|Erythema [first degree] of lip(s)|Erythema [first degree] of lip(s)
C0433307|T037|AB|941.14|ICD9CM|1st deg burn chin|1st deg burn chin
C0433307|T037|PT|941.14|ICD9CM|Erythema [first degree] of chin|Erythema [first degree] of chin
C0161050|T037|AB|941.15|ICD9CM|1st deg burn nose|1st deg burn nose
C0161050|T037|PT|941.15|ICD9CM|Erythema [first degree] of nose (septum)|Erythema [first degree] of nose (septum)
C0375673|T037|AB|941.16|ICD9CM|1st deg burn scalp|1st deg burn scalp
C0375673|T037|PT|941.16|ICD9CM|Erythema [first degree] of scalp [any part]|Erythema [first degree] of scalp [any part]
C0161052|T037|AB|941.17|ICD9CM|1st deg burn face NEC|1st deg burn face NEC
C0161052|T037|PT|941.17|ICD9CM|Erythema [first degree] of forehead and cheek|Erythema [first degree] of forehead and cheek
C0161053|T037|AB|941.18|ICD9CM|1st deg burn neck|1st deg burn neck
C0161053|T037|PT|941.18|ICD9CM|Erythema [first degree] of neck|Erythema [first degree] of neck
C0161054|T037|AB|941.19|ICD9CM|1st deg burn head-mult|1st deg burn head-mult
C0161054|T037|PT|941.19|ICD9CM|Erythema [first degree] of multiple sites [except with eye] of face, head, and neck|Erythema [first degree] of multiple sites [except with eye] of face, head, and neck
C0161055|T037|HT|941.2|ICD9CM|Blisters with epidermal loss due to burn [second degree] of face, head, and neck|Blisters with epidermal loss due to burn [second degree] of face, head, and neck
C0375674|T037|AB|941.20|ICD9CM|2nd deg burn head NOS|2nd deg burn head NOS
C0375674|T037|PT|941.20|ICD9CM|Blisters, epidermal loss [second degree] of face and head, unspecified site|Blisters, epidermal loss [second degree] of face and head, unspecified site
C0273948|T037|AB|941.21|ICD9CM|2nd deg burn ear|2nd deg burn ear
C0273948|T037|PT|941.21|ICD9CM|Blisters, epidermal loss [second degree] of ear [any part]|Blisters, epidermal loss [second degree] of ear [any part]
C0161058|T037|AB|941.22|ICD9CM|2nd deg burn eye|2nd deg burn eye
C0161058|T037|PT|941.22|ICD9CM|Blisters, epidermal loss [second degree] of eye (with other parts of face, head, and neck)|Blisters, epidermal loss [second degree] of eye (with other parts of face, head, and neck)
C0161059|T037|AB|941.23|ICD9CM|2nd deg burn lip|2nd deg burn lip
C0161059|T037|PT|941.23|ICD9CM|Blisters, epidermal loss [second degree] of lip(s)|Blisters, epidermal loss [second degree] of lip(s)
C0161060|T037|AB|941.24|ICD9CM|2nd deg burn chin|2nd deg burn chin
C0161060|T037|PT|941.24|ICD9CM|Blisters, epidermal loss [second degree] of chin|Blisters, epidermal loss [second degree] of chin
C0161061|T037|AB|941.25|ICD9CM|2nd deg burn nose|2nd deg burn nose
C0161061|T037|PT|941.25|ICD9CM|Blisters, epidermal loss [second degree] of nose (septum)|Blisters, epidermal loss [second degree] of nose (septum)
C0161062|T037|AB|941.26|ICD9CM|2nd deg burn scalp|2nd deg burn scalp
C0161062|T037|PT|941.26|ICD9CM|Blisters, epidermal loss [second degree] of scalp [any part]|Blisters, epidermal loss [second degree] of scalp [any part]
C0161063|T037|AB|941.27|ICD9CM|2nd deg burn face NEC|2nd deg burn face NEC
C0161063|T037|PT|941.27|ICD9CM|Blisters, epidermal loss [second degree] of forehead and cheek|Blisters, epidermal loss [second degree] of forehead and cheek
C0161064|T037|AB|941.28|ICD9CM|2nd deg burn neck|2nd deg burn neck
C0161064|T037|PT|941.28|ICD9CM|Blisters, epidermal loss [second degree] of neck|Blisters, epidermal loss [second degree] of neck
C0161065|T037|AB|941.29|ICD9CM|2nd deg burn head-mult|2nd deg burn head-mult
C0161065|T037|PT|941.29|ICD9CM|Blisters, epidermal loss [second degree] of multiple sites [except with eye] of face, head, and neck|Blisters, epidermal loss [second degree] of multiple sites [except with eye] of face, head, and neck
C0161066|T037|HT|941.3|ICD9CM|Full-thickness skin loss due to burn [third degree NOS] of face, head, and neck|Full-thickness skin loss due to burn [third degree NOS] of face, head, and neck
C0161067|T037|AB|941.30|ICD9CM|3rd deg burn head NOS|3rd deg burn head NOS
C0161067|T037|PT|941.30|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of face and head, unspecified site|Full-thickness skin loss [third degree, not otherwise specified] of face and head, unspecified site
C0161068|T037|AB|941.31|ICD9CM|3rd deg burn ear|3rd deg burn ear
C0161068|T037|PT|941.31|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of ear [any part]|Full-thickness skin loss [third degree, not otherwise specified] of ear [any part]
C0161069|T037|AB|941.32|ICD9CM|3rd deg burn eye|3rd deg burn eye
C0161070|T037|AB|941.33|ICD9CM|3rd deg burn lip|3rd deg burn lip
C0161070|T037|PT|941.33|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of lip(s)|Full-thickness skin loss [third degree, not otherwise specified] of lip(s)
C0161071|T037|AB|941.34|ICD9CM|3rd deg burn chin|3rd deg burn chin
C0161071|T037|PT|941.34|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of chin|Full-thickness skin loss [third degree, not otherwise specified] of chin
C0161072|T037|AB|941.35|ICD9CM|3rd deg burn nose|3rd deg burn nose
C0161072|T037|PT|941.35|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of nose (septum)|Full-thickness skin loss [third degree, not otherwise specified] of nose (septum)
C0161073|T037|AB|941.36|ICD9CM|3rd deg burn scalp|3rd deg burn scalp
C0161073|T037|PT|941.36|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of scalp [any part]|Full-thickness skin loss [third degree, not otherwise specified] of scalp [any part]
C0161074|T037|AB|941.37|ICD9CM|3rd deg burn face NEC|3rd deg burn face NEC
C0161074|T037|PT|941.37|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of forehead and cheek|Full-thickness skin loss [third degree, not otherwise specified] of forehead and cheek
C0161075|T037|AB|941.38|ICD9CM|3rd deg burn neck|3rd deg burn neck
C0161075|T037|PT|941.38|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of neck|Full-thickness skin loss [third degree, not otherwise specified] of neck
C0161076|T037|AB|941.39|ICD9CM|3rd deg burn head-mult|3rd deg burn head-mult
C0161078|T037|AB|941.40|ICD9CM|Deep 3 deg burn head NOS|Deep 3 deg burn head NOS
C0161079|T037|AB|941.41|ICD9CM|Deep 3rd deg burn ear|Deep 3rd deg burn ear
C0161080|T037|AB|941.42|ICD9CM|Deep 3rd deg burn eye|Deep 3rd deg burn eye
C0161081|T037|AB|941.43|ICD9CM|Deep 3rd deg burn lip|Deep 3rd deg burn lip
C0161082|T037|AB|941.44|ICD9CM|Deep 3rd deg burn chin|Deep 3rd deg burn chin
C0161083|T037|AB|941.45|ICD9CM|Deep 3rd deg burn nose|Deep 3rd deg burn nose
C0161084|T037|AB|941.46|ICD9CM|Deep 3rd deg burn scalp|Deep 3rd deg burn scalp
C0161085|T037|AB|941.47|ICD9CM|Deep 3rd burn face NEC|Deep 3rd burn face NEC
C0161086|T037|AB|941.48|ICD9CM|Deep 3rd deg burn neck|Deep 3rd deg burn neck
C0161087|T037|AB|941.49|ICD9CM|Deep 3 deg brn head-mult|Deep 3 deg brn head-mult
C0161089|T037|AB|941.50|ICD9CM|3rd burn w loss-head NOS|3rd burn w loss-head NOS
C0161090|T037|AB|941.51|ICD9CM|3rd deg burn w loss-ear|3rd deg burn w loss-ear
C0161090|T037|PT|941.51|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of ear [any part]|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of ear [any part]
C0161091|T037|AB|941.52|ICD9CM|3rd deg burn w loss-eye|3rd deg burn w loss-eye
C0161092|T037|AB|941.53|ICD9CM|3rd deg burn w loss-lip|3rd deg burn w loss-lip
C0161092|T037|PT|941.53|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of lip(s)|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of lip(s)
C0161093|T037|AB|941.54|ICD9CM|3rd deg burn w loss-chin|3rd deg burn w loss-chin
C0161093|T037|PT|941.54|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of chin|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of chin
C0161094|T037|AB|941.55|ICD9CM|3rd deg burn w loss-nose|3rd deg burn w loss-nose
C0161094|T037|PT|941.55|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of nose (septum)|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of nose (septum)
C0161095|T037|AB|941.56|ICD9CM|3rd deg brn w loss-scalp|3rd deg brn w loss-scalp
C0161096|T037|AB|941.57|ICD9CM|3rd burn w loss-face NEC|3rd burn w loss-face NEC
C0161097|T037|AB|941.58|ICD9CM|3rd deg burn w loss-neck|3rd deg burn w loss-neck
C0161097|T037|PT|941.58|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of neck|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of neck
C0161098|T037|AB|941.59|ICD9CM|3rd brn w loss-head mult|3rd brn w loss-head mult
C0161099|T037|HT|942|ICD9CM|Burn of trunk|Burn of trunk
C1812614|T037|HT|942.0|ICD9CM|Burn of trunk, unspecified degree|Burn of trunk, unspecified degree
C1812615|T037|AB|942.00|ICD9CM|Burn NOS trunk-unspec|Burn NOS trunk-unspec
C1812615|T037|PT|942.00|ICD9CM|Burn of unspecified degree of trunk, unspecified site|Burn of unspecified degree of trunk, unspecified site
C0273993|T037|AB|942.01|ICD9CM|Burn NOS breast|Burn NOS breast
C0273993|T037|PT|942.01|ICD9CM|Burn of unspecified degree of breast|Burn of unspecified degree of breast
C0840791|T037|AB|942.02|ICD9CM|Burn NOS chest wall|Burn NOS chest wall
C0840791|T037|PT|942.02|ICD9CM|Burn of unspecified degree of chest wall, excluding breast and nipple|Burn of unspecified degree of chest wall, excluding breast and nipple
C0274005|T037|AB|942.03|ICD9CM|Burn NOS abdominal wall|Burn NOS abdominal wall
C0274005|T037|PT|942.03|ICD9CM|Burn of unspecified degree of abdominal wall|Burn of unspecified degree of abdominal wall
C0274011|T037|AB|942.04|ICD9CM|Burn NOS back|Burn NOS back
C0274011|T037|PT|942.04|ICD9CM|Burn of unspecified degree of back [any part]|Burn of unspecified degree of back [any part]
C0161105|T037|AB|942.05|ICD9CM|Burn NOS genitalia|Burn NOS genitalia
C0161105|T037|PT|942.05|ICD9CM|Burn of unspecified degree of genitalia|Burn of unspecified degree of genitalia
C0161106|T037|AB|942.09|ICD9CM|Burn NOS trunk NEC|Burn NOS trunk NEC
C0161106|T037|PT|942.09|ICD9CM|Burn of unspecified degree of other and multiple sites of trunk|Burn of unspecified degree of other and multiple sites of trunk
C0161107|T037|HT|942.1|ICD9CM|Erythema due to burn [first degree] of trunk|Erythema due to burn [first degree] of trunk
C0840795|T037|AB|942.10|ICD9CM|1st deg burn trunk NOS|1st deg burn trunk NOS
C0840795|T037|PT|942.10|ICD9CM|Erythema [first degree] of trunk, unspecified site|Erythema [first degree] of trunk, unspecified site
C0161109|T037|AB|942.11|ICD9CM|1st deg burn breast|1st deg burn breast
C0161109|T037|PT|942.11|ICD9CM|Erythema [first degree] of breast|Erythema [first degree] of breast
C0161110|T037|AB|942.12|ICD9CM|1st deg burn chest wall|1st deg burn chest wall
C0161110|T037|PT|942.12|ICD9CM|Erythema [first degree] of chest wall, excluding breast and nipple|Erythema [first degree] of chest wall, excluding breast and nipple
C0840797|T037|AB|942.13|ICD9CM|1st deg burn abdomn wall|1st deg burn abdomn wall
C0840797|T037|PT|942.13|ICD9CM|Erythema [first degree] of abdominal wall|Erythema [first degree] of abdominal wall
C0840798|T037|AB|942.14|ICD9CM|1st deg burn back|1st deg burn back
C0840798|T037|PT|942.14|ICD9CM|Erythema [first degree] of back [any part]|Erythema [first degree] of back [any part]
C0161113|T037|AB|942.15|ICD9CM|1st deg burn genitalia|1st deg burn genitalia
C0161113|T037|PT|942.15|ICD9CM|Erythema [first degree] of genitalia|Erythema [first degree] of genitalia
C0161114|T037|AB|942.19|ICD9CM|1st deg burn trunk NEC|1st deg burn trunk NEC
C0161114|T037|PT|942.19|ICD9CM|Erythema [first degree] of other and multiple sites of trunk|Erythema [first degree] of other and multiple sites of trunk
C0433353|T037|HT|942.2|ICD9CM|Blisters with epidermal loss due to burn [second degree] of trunk|Blisters with epidermal loss due to burn [second degree] of trunk
C0840801|T037|AB|942.20|ICD9CM|2nd deg burn trunk NOS|2nd deg burn trunk NOS
C0840801|T037|PT|942.20|ICD9CM|Blisters, epidermal loss [second degree] of trunk, unspecified site|Blisters, epidermal loss [second degree] of trunk, unspecified site
C0840802|T037|AB|942.21|ICD9CM|2nd deg burn breast|2nd deg burn breast
C0840802|T037|PT|942.21|ICD9CM|Blisters, epidermal loss [second degree] of breast|Blisters, epidermal loss [second degree] of breast
C0161118|T037|AB|942.22|ICD9CM|2nd deg burn chest wall|2nd deg burn chest wall
C0161118|T037|PT|942.22|ICD9CM|Blisters, epidermal loss [second degree] of chest wall, excluding breast and nipple|Blisters, epidermal loss [second degree] of chest wall, excluding breast and nipple
C0840804|T037|AB|942.23|ICD9CM|2nd deg burn abdomn wall|2nd deg burn abdomn wall
C0840804|T037|PT|942.23|ICD9CM|Blisters, epidermal loss [second degree] of abdominal wall|Blisters, epidermal loss [second degree] of abdominal wall
C0840805|T037|AB|942.24|ICD9CM|2nd deg burn back|2nd deg burn back
C0840805|T037|PT|942.24|ICD9CM|Blisters, epidermal loss [second degree] of back [any part]|Blisters, epidermal loss [second degree] of back [any part]
C0161121|T037|AB|942.25|ICD9CM|2nd deg burn genitalia|2nd deg burn genitalia
C0161121|T037|PT|942.25|ICD9CM|Blisters, epidermal loss [second degree] of genitalia|Blisters, epidermal loss [second degree] of genitalia
C0161122|T037|AB|942.29|ICD9CM|2nd deg burn trunk NEC|2nd deg burn trunk NEC
C0161122|T037|PT|942.29|ICD9CM|Blisters, epidermal loss [second degree] of other and multiple sites of trunk|Blisters, epidermal loss [second degree] of other and multiple sites of trunk
C0161123|T037|HT|942.3|ICD9CM|Full-thickness skin loss due to burn [third degree NOS] of trunk|Full-thickness skin loss due to burn [third degree NOS] of trunk
C0840808|T037|AB|942.30|ICD9CM|3rd deg burn trunk NOS|3rd deg burn trunk NOS
C0840808|T037|PT|942.30|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of trunk, unspecified site|Full-thickness skin loss [third degree, not otherwise specified] of trunk, unspecified site
C0433480|T037|AB|942.31|ICD9CM|3rd deg burn breast|3rd deg burn breast
C0433480|T037|PT|942.31|ICD9CM|Full-thickness skin loss [third degree,not otherwise specified] of breast|Full-thickness skin loss [third degree,not otherwise specified] of breast
C0161126|T037|AB|942.32|ICD9CM|3rd deg burn chest wall|3rd deg burn chest wall
C0433482|T037|AB|942.33|ICD9CM|3rd deg burn abdomn wall|3rd deg burn abdomn wall
C0433482|T037|PT|942.33|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of abdominal wall|Full-thickness skin loss [third degree, not otherwise specified] of abdominal wall
C0840810|T037|AB|942.34|ICD9CM|3rd deg burn back|3rd deg burn back
C0840810|T037|PT|942.34|ICD9CM|Full-thickness skin loss [third degree,not otherwise specified] of back [any part]|Full-thickness skin loss [third degree,not otherwise specified] of back [any part]
C0161129|T037|AB|942.35|ICD9CM|3rd deg burn genitalia|3rd deg burn genitalia
C0161129|T037|PT|942.35|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of genitalia|Full-thickness skin loss [third degree, not otherwise specified] of genitalia
C0161130|T037|AB|942.39|ICD9CM|3rd deg burn trunk NEC|3rd deg burn trunk NEC
C0161132|T037|AB|942.40|ICD9CM|Deep 3rd burn trunk NOS|Deep 3rd burn trunk NOS
C0161133|T037|AB|942.41|ICD9CM|Deep 3rd deg burn breast|Deep 3rd deg burn breast
C0161134|T037|AB|942.42|ICD9CM|Deep 3rd burn chest wall|Deep 3rd burn chest wall
C0375675|T037|AB|942.43|ICD9CM|Deep 3rd burn abdom wall|Deep 3rd burn abdom wall
C0375676|T047|AB|942.44|ICD9CM|Deep 3rd deg burn back|Deep 3rd deg burn back
C0375677|T047|AB|942.45|ICD9CM|Deep 3rd burn genitalia|Deep 3rd burn genitalia
C0161138|T037|AB|942.49|ICD9CM|Deep 3rd burn trunk NEC|Deep 3rd burn trunk NEC
C0161140|T037|AB|942.50|ICD9CM|3rd brn w loss-trunk NOS|3rd brn w loss-trunk NOS
C0161141|T037|AB|942.51|ICD9CM|3rd burn w loss-breast|3rd burn w loss-breast
C0161141|T037|PT|942.51|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of breast|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of breast
C0161142|T037|AB|942.52|ICD9CM|3rd brn w loss-chest wll|3rd brn w loss-chest wll
C0375678|T037|AB|942.53|ICD9CM|3rd brn w loss-abdom wll|3rd brn w loss-abdom wll
C0375678|T037|PT|942.53|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of abdominal wall|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of abdominal wall
C0375679|T037|AB|942.54|ICD9CM|3rd deg burn w loss-back|3rd deg burn w loss-back
C0375679|T037|PT|942.54|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of back [any part]|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of back [any part]
C0375680|T037|AB|942.55|ICD9CM|3rd brn w loss-genitalia|3rd brn w loss-genitalia
C0375680|T037|PT|942.55|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of genitalia|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of genitalia
C0161146|T037|AB|942.59|ICD9CM|3rd brn w loss-trunk NEC|3rd brn w loss-trunk NEC
C0433193|T037|HT|943|ICD9CM|Burn of upper limb, except wrist and hand|Burn of upper limb, except wrist and hand
C0375681|T037|HT|943.0|ICD9CM|Burn of upper limb, except wrist and hand, unspecified degree|Burn of upper limb, except wrist and hand, unspecified degree
C0274035|T037|AB|943.00|ICD9CM|Burn NOS arm-unspec|Burn NOS arm-unspec
C0274035|T037|PT|943.00|ICD9CM|Burn of unspecified degree of upper limb, except wrist and hand, unspecified site|Burn of unspecified degree of upper limb, except wrist and hand, unspecified site
C0274071|T037|AB|943.01|ICD9CM|Burn NOS forearm|Burn NOS forearm
C0274071|T037|PT|943.01|ICD9CM|Burn of unspecified degree of forearm|Burn of unspecified degree of forearm
C0274065|T037|AB|943.02|ICD9CM|Burn NOS elbow|Burn NOS elbow
C0274065|T037|PT|943.02|ICD9CM|Burn of unspecified degree of elbow|Burn of unspecified degree of elbow
C0161151|T037|AB|943.03|ICD9CM|Burn NOS upper arm|Burn NOS upper arm
C0161151|T037|PT|943.03|ICD9CM|Burn of unspecified degree of upper arm|Burn of unspecified degree of upper arm
C0274053|T037|AB|943.04|ICD9CM|Burn NOS axilla|Burn NOS axilla
C0274053|T037|PT|943.04|ICD9CM|Burn of unspecified degree of axilla|Burn of unspecified degree of axilla
C0274041|T037|AB|943.05|ICD9CM|Burn NOS shoulder|Burn NOS shoulder
C0274041|T037|PT|943.05|ICD9CM|Burn of unspecified degree of shoulder|Burn of unspecified degree of shoulder
C0274047|T037|AB|943.06|ICD9CM|Burn NOS scapula|Burn NOS scapula
C0274047|T037|PT|943.06|ICD9CM|Burn of unspecified degree of scapular region|Burn of unspecified degree of scapular region
C0161155|T037|AB|943.09|ICD9CM|Burn NOS arm-multiple|Burn NOS arm-multiple
C0161155|T037|PT|943.09|ICD9CM|Burn of unspecified degree of multiple sites of upper limb, except wrist and hand|Burn of unspecified degree of multiple sites of upper limb, except wrist and hand
C0161156|T037|HT|943.1|ICD9CM|Erythema due to burn [first degree] of upper limb, except wrist and hand|Erythema due to burn [first degree] of upper limb, except wrist and hand
C0161157|T037|AB|943.10|ICD9CM|1st deg burn arm NOS|1st deg burn arm NOS
C0161157|T037|PT|943.10|ICD9CM|Erythema [first degree] of upper limb, unspecified site|Erythema [first degree] of upper limb, unspecified site
C0161158|T037|AB|943.11|ICD9CM|1st deg burn forearm|1st deg burn forearm
C0161158|T037|PT|943.11|ICD9CM|Erythema [first degree] of forearm|Erythema [first degree] of forearm
C0161159|T037|AB|943.12|ICD9CM|1st deg burn elbow|1st deg burn elbow
C0161159|T037|PT|943.12|ICD9CM|Erythema [first degree] of elbow|Erythema [first degree] of elbow
C0161160|T037|AB|943.13|ICD9CM|1st deg burn upper arm|1st deg burn upper arm
C0161160|T037|PT|943.13|ICD9CM|Erythema [first degree] of upper arm|Erythema [first degree] of upper arm
C0161161|T037|AB|943.14|ICD9CM|1st deg burn axilla|1st deg burn axilla
C0161161|T037|PT|943.14|ICD9CM|Erythema [first degree] of axilla|Erythema [first degree] of axilla
C0161162|T037|AB|943.15|ICD9CM|1st deg burn shoulder|1st deg burn shoulder
C0161162|T037|PT|943.15|ICD9CM|Erythema [first degree] of shoulder|Erythema [first degree] of shoulder
C0161163|T037|AB|943.16|ICD9CM|1st deg burn scapula|1st deg burn scapula
C0161163|T037|PT|943.16|ICD9CM|Erythema [first degree] of scapular region|Erythema [first degree] of scapular region
C0161164|T037|AB|943.19|ICD9CM|1st deg burn arm-mult|1st deg burn arm-mult
C0161164|T037|PT|943.19|ICD9CM|Erythema [first degree] of multiple sites of upper limb, except wrist and hand|Erythema [first degree] of multiple sites of upper limb, except wrist and hand
C0161165|T037|HT|943.2|ICD9CM|Blisters with epidermal loss due to burn [second degree] of upper limb, except wrist and hand|Blisters with epidermal loss due to burn [second degree] of upper limb, except wrist and hand
C0161166|T037|AB|943.20|ICD9CM|2nd deg burn arm NOS|2nd deg burn arm NOS
C0161166|T037|PT|943.20|ICD9CM|Blisters, epidermal loss [second degree] of upper limb, unspecified site|Blisters, epidermal loss [second degree] of upper limb, unspecified site
C0161167|T037|AB|943.21|ICD9CM|2nd deg burn forearm|2nd deg burn forearm
C0161167|T037|PT|943.21|ICD9CM|Blisters, epidermal loss [second degree] of forearm|Blisters, epidermal loss [second degree] of forearm
C0161168|T037|AB|943.22|ICD9CM|2nd deg burn elbow|2nd deg burn elbow
C0161168|T037|PT|943.22|ICD9CM|Blisters, epidermal loss [second degree] of elbow|Blisters, epidermal loss [second degree] of elbow
C0161169|T037|AB|943.23|ICD9CM|2nd deg burn upper arm|2nd deg burn upper arm
C0161169|T037|PT|943.23|ICD9CM|Blisters, epidermal loss [second degree] of upper arm|Blisters, epidermal loss [second degree] of upper arm
C0161170|T037|AB|943.24|ICD9CM|2nd deg burn axilla|2nd deg burn axilla
C0161170|T037|PT|943.24|ICD9CM|Blisters, epidermal loss [second degree] of axilla|Blisters, epidermal loss [second degree] of axilla
C0161171|T037|AB|943.25|ICD9CM|2nd deg burn shoulder|2nd deg burn shoulder
C0161171|T037|PT|943.25|ICD9CM|Blisters, epidermal loss [second degree] of shoulder|Blisters, epidermal loss [second degree] of shoulder
C0161172|T037|AB|943.26|ICD9CM|2nd deg burn scapula|2nd deg burn scapula
C0161172|T037|PT|943.26|ICD9CM|Blisters, epidermal loss [second degree] of scapular region|Blisters, epidermal loss [second degree] of scapular region
C0161173|T037|AB|943.29|ICD9CM|2nd deg burn arm-mult|2nd deg burn arm-mult
C0161173|T037|PT|943.29|ICD9CM|Blisters, epidermal loss [second degree] of multiple sites of upper limb, except wrist and hand|Blisters, epidermal loss [second degree] of multiple sites of upper limb, except wrist and hand
C0161174|T037|HT|943.3|ICD9CM|Full-thickness skin loss due to burn [third degree NOS] of upper limb, except wrist and hand|Full-thickness skin loss due to burn [third degree NOS] of upper limb, except wrist and hand
C0161175|T037|AB|943.30|ICD9CM|3rd deg burn arm NOS|3rd deg burn arm NOS
C0161175|T037|PT|943.30|ICD9CM|Full-thickness skin [third degree, not otherwise specified] of upper limb, unspecified site|Full-thickness skin [third degree, not otherwise specified] of upper limb, unspecified site
C0161176|T037|AB|943.31|ICD9CM|3rd deg burn forearm|3rd deg burn forearm
C0161176|T037|PT|943.31|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of forearm|Full-thickness skin loss [third degree, not otherwise specified] of forearm
C0161177|T037|AB|943.32|ICD9CM|3rd deg burn elbow|3rd deg burn elbow
C0161177|T037|PT|943.32|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of elbow|Full-thickness skin loss [third degree, not otherwise specified] of elbow
C0161178|T037|AB|943.33|ICD9CM|3rd deg burn upper arm|3rd deg burn upper arm
C0161178|T037|PT|943.33|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of upper arm|Full-thickness skin loss [third degree, not otherwise specified] of upper arm
C0274056|T037|AB|943.34|ICD9CM|3rd deg burn axilla|3rd deg burn axilla
C0274056|T037|PT|943.34|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of axilla|Full-thickness skin loss [third degree, not otherwise specified] of axilla
C0161180|T037|AB|943.35|ICD9CM|3rd deg burn shoulder|3rd deg burn shoulder
C0161180|T037|PT|943.35|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of shoulder|Full-thickness skin loss [third degree, not otherwise specified] of shoulder
C0161181|T037|AB|943.36|ICD9CM|3rd deg burn scapula|3rd deg burn scapula
C0161181|T037|PT|943.36|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of scapular region|Full-thickness skin loss [third degree, not otherwise specified] of scapular region
C0161182|T037|AB|943.39|ICD9CM|3rd deg burn arm-mult|3rd deg burn arm-mult
C0161184|T037|AB|943.40|ICD9CM|Deep 3 deg burn arm NOS|Deep 3 deg burn arm NOS
C0161185|T037|AB|943.41|ICD9CM|Deep 3 deg burn forearm|Deep 3 deg burn forearm
C0161186|T037|AB|943.42|ICD9CM|Deep 3 deg burn elbow|Deep 3 deg burn elbow
C0161187|T037|AB|943.43|ICD9CM|Deep 3 deg brn upper arm|Deep 3 deg brn upper arm
C0161188|T037|AB|943.44|ICD9CM|Deep 3 deg burn axilla|Deep 3 deg burn axilla
C0161189|T037|AB|943.45|ICD9CM|Deep 3 deg burn shoulder|Deep 3 deg burn shoulder
C0161190|T037|AB|943.46|ICD9CM|Deep 3 deg burn scapula|Deep 3 deg burn scapula
C0161191|T037|AB|943.49|ICD9CM|Deep 3 deg burn arm-mult|Deep 3 deg burn arm-mult
C0161193|T037|AB|943.50|ICD9CM|3rd burn w loss-arm NOS|3rd burn w loss-arm NOS
C0161194|T037|AB|943.51|ICD9CM|3rd burn w loss-forearm|3rd burn w loss-forearm
C0161194|T037|PT|943.51|ICD9CM|Deep necrosis of underlying tissues [deep third degree) with loss of a body part, of forearm|Deep necrosis of underlying tissues [deep third degree) with loss of a body part, of forearm
C0161195|T037|AB|943.52|ICD9CM|3rd burn w loss-elbow|3rd burn w loss-elbow
C0161195|T037|PT|943.52|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of elbow|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of elbow
C0161196|T037|AB|943.53|ICD9CM|3rd brn w loss-upper arm|3rd brn w loss-upper arm
C0161196|T037|PT|943.53|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of upper arm|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of upper arm
C0161197|T037|AB|943.54|ICD9CM|3rd burn w loss-axilla|3rd burn w loss-axilla
C0161197|T037|PT|943.54|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of axilla|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of axilla
C0161198|T037|AB|943.55|ICD9CM|3rd burn w loss-shoulder|3rd burn w loss-shoulder
C0161198|T037|PT|943.55|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of shoulder|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of shoulder
C0161199|T037|AB|943.56|ICD9CM|3rd burn w loss-scapula|3rd burn w loss-scapula
C0161199|T037|PT|943.56|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of scapular region|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of scapular region
C0161200|T037|AB|943.59|ICD9CM|3rd burn w loss arm-mult|3rd burn w loss arm-mult
C0433205|T037|HT|944|ICD9CM|Burn of wrist(s) and hand(s)|Burn of wrist(s) and hand(s)
C1812619|T037|HT|944.0|ICD9CM|Burn of wrist(s) and hand(s), unspecified degree|Burn of wrist(s) and hand(s), unspecified degree
C0274089|T037|AB|944.00|ICD9CM|Burn NOS hand-unspec|Burn NOS hand-unspec
C0274089|T037|PT|944.00|ICD9CM|Burn of unspecified degree of hand, unspecified site|Burn of unspecified degree of hand, unspecified site
C0161203|T037|AB|944.01|ICD9CM|Burn NOS finger|Burn NOS finger
C0161203|T037|PT|944.01|ICD9CM|Burn of unspecified degree of single digit (finger (nail) other than thumb|Burn of unspecified degree of single digit (finger (nail) other than thumb
C0161204|T037|AB|944.02|ICD9CM|Burn NOS thumb|Burn NOS thumb
C0161204|T037|PT|944.02|ICD9CM|Burn of unspecified degree of thumb (nail)|Burn of unspecified degree of thumb (nail)
C0161205|T037|AB|944.03|ICD9CM|Burn NOS mult fingers|Burn NOS mult fingers
C0161205|T037|PT|944.03|ICD9CM|Burn of unspecified degree of two or more digits of hand, not including thumb|Burn of unspecified degree of two or more digits of hand, not including thumb
C0161206|T037|AB|944.04|ICD9CM|Burn NOS finger w thumb|Burn NOS finger w thumb
C0161206|T037|PT|944.04|ICD9CM|Burn of unspecified degree of two or more digits of hand, including thumb|Burn of unspecified degree of two or more digits of hand, including thumb
C0161207|T037|AB|944.05|ICD9CM|Burn NOS palm|Burn NOS palm
C0161207|T037|PT|944.05|ICD9CM|Burn of unspecified degree of palm|Burn of unspecified degree of palm
C0161208|T037|AB|944.06|ICD9CM|Burn NOS back of hand|Burn NOS back of hand
C0161208|T037|PT|944.06|ICD9CM|Burn of unspecified degree of back of hand|Burn of unspecified degree of back of hand
C0274083|T037|AB|944.07|ICD9CM|Burn NOS wrist|Burn NOS wrist
C0274083|T037|PT|944.07|ICD9CM|Burn of unspecified degree of wrist|Burn of unspecified degree of wrist
C0161210|T037|AB|944.08|ICD9CM|Burn NOS hand-multiple|Burn NOS hand-multiple
C0161210|T037|PT|944.08|ICD9CM|Burn of unspecified degree of multiple sites of wrist(s) and hand(s)|Burn of unspecified degree of multiple sites of wrist(s) and hand(s)
C0161211|T037|HT|944.1|ICD9CM|Erythema due to burn [first degree] of wrist(s) and hand(s)|Erythema due to burn [first degree] of wrist(s) and hand(s)
C0274090|T037|AB|944.10|ICD9CM|1st deg burn hand NOS|1st deg burn hand NOS
C0274090|T037|PT|944.10|ICD9CM|Erythema [first degree] of hand, unspecified site|Erythema [first degree] of hand, unspecified site
C0161213|T037|AB|944.11|ICD9CM|1st deg burn finger|1st deg burn finger
C0161213|T037|PT|944.11|ICD9CM|Erythema [first degree] of single digit (finger (nail)) other than thumb|Erythema [first degree] of single digit (finger (nail)) other than thumb
C0161214|T037|AB|944.12|ICD9CM|1st deg burn thumb|1st deg burn thumb
C0161214|T037|PT|944.12|ICD9CM|Erythema [first degree] of thumb (nail)|Erythema [first degree] of thumb (nail)
C0161215|T037|AB|944.13|ICD9CM|1st deg burn mult finger|1st deg burn mult finger
C0161215|T037|PT|944.13|ICD9CM|Erythema [first degree] of two or more digits of hand, not including thumb|Erythema [first degree] of two or more digits of hand, not including thumb
C1112529|T037|AB|944.14|ICD9CM|1 deg burn fingr w thumb|1 deg burn fingr w thumb
C1112529|T037|PT|944.14|ICD9CM|Erythema [first degree] of two or more digits of hand including thumb|Erythema [first degree] of two or more digits of hand including thumb
C0161217|T037|AB|944.15|ICD9CM|1st deg burn palm|1st deg burn palm
C0161217|T037|PT|944.15|ICD9CM|Erythema [first degree] of palm|Erythema [first degree] of palm
C0433333|T037|AB|944.16|ICD9CM|1 deg burn back of hand|1 deg burn back of hand
C0433333|T037|PT|944.16|ICD9CM|Erythema [first degree] of back of hand|Erythema [first degree] of back of hand
C0274084|T037|AB|944.17|ICD9CM|1st deg burn wrist|1st deg burn wrist
C0274084|T037|PT|944.17|ICD9CM|Erythema [first degree] of wrist|Erythema [first degree] of wrist
C0161220|T037|AB|944.18|ICD9CM|1st deg burn hand-mult|1st deg burn hand-mult
C0161220|T037|PT|944.18|ICD9CM|Erythema [first degree] of multiple sites of wrist(s) and hand(s)|Erythema [first degree] of multiple sites of wrist(s) and hand(s)
C0161221|T037|HT|944.2|ICD9CM|Blisters with epidermal loss due to burn [second degree] of wrist(s) and hand(s)|Blisters with epidermal loss due to burn [second degree] of wrist(s) and hand(s)
C0433361|T037|AB|944.20|ICD9CM|2nd deg burn hand NOS|2nd deg burn hand NOS
C0433361|T037|PT|944.20|ICD9CM|Blisters, epidermal loss [second degree] of hand, unspecified site|Blisters, epidermal loss [second degree] of hand, unspecified site
C0161223|T037|AB|944.21|ICD9CM|2nd deg burn finger|2nd deg burn finger
C0161223|T037|PT|944.21|ICD9CM|Blisters, epidermal loss [second degree] of single digit [finger (nail)] other than thumb|Blisters, epidermal loss [second degree] of single digit [finger (nail)] other than thumb
C0161224|T037|AB|944.22|ICD9CM|2nd deg burn thumb|2nd deg burn thumb
C0161224|T037|PT|944.22|ICD9CM|Blisters, epidermal loss [second degree] of thumb (nail)|Blisters, epidermal loss [second degree] of thumb (nail)
C0161225|T037|AB|944.23|ICD9CM|2nd deg burn mult finger|2nd deg burn mult finger
C0161225|T037|PT|944.23|ICD9CM|Blisters, epidermal loss [second degree] of two or more digits of hand, not including thumb|Blisters, epidermal loss [second degree] of two or more digits of hand, not including thumb
C0161226|T037|AB|944.24|ICD9CM|2 deg burn fingr w thumb|2 deg burn fingr w thumb
C0161226|T037|PT|944.24|ICD9CM|Blisters, epidermal loss [second degree] of two or more digits of hand including thumb|Blisters, epidermal loss [second degree] of two or more digits of hand including thumb
C0161227|T037|AB|944.25|ICD9CM|2nd deg burn palm|2nd deg burn palm
C0161227|T037|PT|944.25|ICD9CM|Blisters, epidermal loss [second degree] of palm|Blisters, epidermal loss [second degree] of palm
C0161228|T037|AB|944.26|ICD9CM|2 deg burn back of hand|2 deg burn back of hand
C0161228|T037|PT|944.26|ICD9CM|Blisters , epidermal loss [second degree] of back of hand|Blisters , epidermal loss [second degree] of back of hand
C1443011|T037|AB|944.27|ICD9CM|2nd deg burn wrist|2nd deg burn wrist
C1443011|T037|PT|944.27|ICD9CM|Blisters, epidermal loss [second degree] of wrist|Blisters, epidermal loss [second degree] of wrist
C0161230|T037|AB|944.28|ICD9CM|2nd deg burn hand-mult|2nd deg burn hand-mult
C0161230|T037|PT|944.28|ICD9CM|Blisters, epidermal loss [second degree] of multiple sites of wrist(s) and hand(s)|Blisters, epidermal loss [second degree] of multiple sites of wrist(s) and hand(s)
C0274134|T037|HT|944.3|ICD9CM|Full-thickness skin loss due to burn [third degree NOS] of wrist(s) and hand(s)|Full-thickness skin loss due to burn [third degree NOS] of wrist(s) and hand(s)
C0161232|T037|AB|944.30|ICD9CM|3rd deg burn hand NOS|3rd deg burn hand NOS
C0161232|T037|PT|944.30|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of hand, unspecified site|Full-thickness skin loss [third degree, not otherwise specified] of hand, unspecified site
C0161233|T037|AB|944.31|ICD9CM|3rd deg burn finger|3rd deg burn finger
C0161234|T037|AB|944.32|ICD9CM|3rd deg burn thumb|3rd deg burn thumb
C0161234|T037|PT|944.32|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of thumb (nail)|Full-thickness skin loss [third degree, not otherwise specified] of thumb (nail)
C0161235|T037|AB|944.33|ICD9CM|3rd deg burn mult finger|3rd deg burn mult finger
C0161236|T037|AB|944.34|ICD9CM|3 deg burn fingr w thumb|3 deg burn fingr w thumb
C0161237|T037|AB|944.35|ICD9CM|3rd deg burn palm|3rd deg burn palm
C0161237|T037|PT|944.35|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of palm of hand|Full-thickness skin loss [third degree, not otherwise specified] of palm of hand
C0161238|T037|AB|944.36|ICD9CM|3 deg burn back of hand|3 deg burn back of hand
C0161238|T037|PT|944.36|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of back of hand|Full-thickness skin loss [third degree, not otherwise specified] of back of hand
C1443010|T037|AB|944.37|ICD9CM|3rd deg burn wrist|3rd deg burn wrist
C1443010|T037|PT|944.37|ICD9CM|Full-thickness skin loss [third degree, not otherwise specified] of wrist|Full-thickness skin loss [third degree, not otherwise specified] of wrist
C0161240|T037|AB|944.38|ICD9CM|3rd deg burn hand-mult|3rd deg burn hand-mult
C0161242|T037|AB|944.40|ICD9CM|Deep 3 deg brn hand NOS|Deep 3 deg brn hand NOS
C0161243|T037|AB|944.41|ICD9CM|Deep 3 deg burn finger|Deep 3 deg burn finger
C0161244|T037|AB|944.42|ICD9CM|Deep 3 deg burn thumb|Deep 3 deg burn thumb
C0161245|T037|AB|944.43|ICD9CM|Deep 3rd brn mult finger|Deep 3rd brn mult finger
C0161246|T037|AB|944.44|ICD9CM|Deep 3rd brn fngr w thmb|Deep 3rd brn fngr w thmb
C0161247|T037|AB|944.45|ICD9CM|Deep 3 deg burn palm|Deep 3 deg burn palm
C0161248|T037|AB|944.46|ICD9CM|Deep 3rd brn back of hnd|Deep 3rd brn back of hnd
C0161249|T037|AB|944.47|ICD9CM|Deep 3 deg burn wrist|Deep 3 deg burn wrist
C0161250|T037|AB|944.48|ICD9CM|Deep 3 deg brn hand-mult|Deep 3 deg brn hand-mult
C0161252|T037|AB|944.50|ICD9CM|3rd brn w loss-hand NOS|3rd brn w loss-hand NOS
C0161253|T037|AB|944.51|ICD9CM|3rd burn w loss-finger|3rd burn w loss-finger
C0161254|T037|AB|944.52|ICD9CM|3rd burn w loss-thumb|3rd burn w loss-thumb
C0161254|T037|PT|944.52|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of thumb (nail)|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of thumb (nail)
C0161255|T037|AB|944.53|ICD9CM|3rd brn w loss-mult fngr|3rd brn w loss-mult fngr
C0161256|T037|AB|944.54|ICD9CM|3rd brn w loss-fngr/thmb|3rd brn w loss-fngr/thmb
C0161257|T037|AB|944.55|ICD9CM|3rd burn w loss-palm|3rd burn w loss-palm
C0161257|T037|PT|944.55|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of palm of hand|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of palm of hand
C0161258|T037|AB|944.56|ICD9CM|3rd brn w loss-bk of hnd|3rd brn w loss-bk of hnd
C0161258|T037|PT|944.56|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of back of hand|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of back of hand
C0161259|T037|AB|944.57|ICD9CM|3rd burn w loss-wrist|3rd burn w loss-wrist
C0161259|T037|PT|944.57|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of wrist|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of wrist
C0161260|T037|AB|944.58|ICD9CM|3rd brn w loss hand-mult|3rd brn w loss hand-mult
C0274137|T037|HT|945|ICD9CM|Burn of lower limb(s)|Burn of lower limb(s)
C1812618|T037|HT|945.0|ICD9CM|Burn of lower limb(s), unspecified degree|Burn of lower limb(s), unspecified degree
C1812617|T037|AB|945.00|ICD9CM|Burn NOS leg-unspec|Burn NOS leg-unspec
C1812617|T037|PT|945.00|ICD9CM|Burn of unspecified degree of lower limb [leg], unspecified site|Burn of unspecified degree of lower limb [leg], unspecified site
C0161263|T037|AB|945.01|ICD9CM|Burn NOS toe|Burn NOS toe
C0161263|T037|PT|945.01|ICD9CM|Burn of unspecified degree of toe(s) (nail)|Burn of unspecified degree of toe(s) (nail)
C0274167|T037|AB|945.02|ICD9CM|Burn NOS foot|Burn NOS foot
C0274167|T037|PT|945.02|ICD9CM|Burn of unspecified degree of foot|Burn of unspecified degree of foot
C0274161|T037|AB|945.03|ICD9CM|Burn NOS ankle|Burn NOS ankle
C0274161|T037|PT|945.03|ICD9CM|Burn of unspecified degree of ankle|Burn of unspecified degree of ankle
C0274155|T037|AB|945.04|ICD9CM|Burn NOS lower leg|Burn NOS lower leg
C0274155|T037|PT|945.04|ICD9CM|Burn of unspecified degree of lower leg|Burn of unspecified degree of lower leg
C0274149|T037|AB|945.05|ICD9CM|Burn NOS knee|Burn NOS knee
C0274149|T037|PT|945.05|ICD9CM|Burn of unspecified degree of knee|Burn of unspecified degree of knee
C0274143|T037|AB|945.06|ICD9CM|Burn NOS thigh|Burn NOS thigh
C0274143|T037|PT|945.06|ICD9CM|Burn of unspecified degree of thigh [any part]|Burn of unspecified degree of thigh [any part]
C0161269|T037|AB|945.09|ICD9CM|Burn NOS leg-multiple|Burn NOS leg-multiple
C0161269|T037|PT|945.09|ICD9CM|Burn of unspecified degree of multiple sites of lower limb(s)|Burn of unspecified degree of multiple sites of lower limb(s)
C0161270|T037|HT|945.1|ICD9CM|Erythema due to burn [first degree] of lower limb(s)|Erythema due to burn [first degree] of lower limb(s)
C0161271|T037|AB|945.10|ICD9CM|1st deg burn leg NOS|1st deg burn leg NOS
C0161271|T037|PT|945.10|ICD9CM|Erythema [first degree] of lower limb [leg], unspecified site|Erythema [first degree] of lower limb [leg], unspecified site
C0161272|T037|AB|945.11|ICD9CM|1st deg burn toe|1st deg burn toe
C0161272|T037|PT|945.11|ICD9CM|Erythema [first degree] of toe(s) (nail)|Erythema [first degree] of toe(s) (nail)
C0161273|T037|AB|945.12|ICD9CM|1st deg burn foot|1st deg burn foot
C0161273|T037|PT|945.12|ICD9CM|Erythema [first degree] of foot|Erythema [first degree] of foot
C0161274|T037|AB|945.13|ICD9CM|1st deg burn ankle|1st deg burn ankle
C0161274|T037|PT|945.13|ICD9CM|Erythema [first degree] of ankle|Erythema [first degree] of ankle
C0161275|T037|AB|945.14|ICD9CM|1st deg burn lower leg|1st deg burn lower leg
C0161275|T037|PT|945.14|ICD9CM|Erythema [first degree] of lower leg|Erythema [first degree] of lower leg
C0161276|T037|AB|945.15|ICD9CM|1st deg burn knee|1st deg burn knee
C0161276|T037|PT|945.15|ICD9CM|Erythema [first degree] of knee|Erythema [first degree] of knee
C0161277|T037|AB|945.16|ICD9CM|1st deg burn thigh|1st deg burn thigh
C0161277|T037|PT|945.16|ICD9CM|Erythema [first degree] of thigh [any part]|Erythema [first degree] of thigh [any part]
C0161278|T037|AB|945.19|ICD9CM|1st deg burn leg-mult|1st deg burn leg-mult
C0161278|T037|PT|945.19|ICD9CM|Erythema [first degree] of multiple sites of lower limb(s)|Erythema [first degree] of multiple sites of lower limb(s)
C0161279|T037|HT|945.2|ICD9CM|Blisters with epidermal loss due to burn [second degree] of lower limb(s)|Blisters with epidermal loss due to burn [second degree] of lower limb(s)
C0161280|T037|AB|945.20|ICD9CM|2nd deg burn leg NOS|2nd deg burn leg NOS
C0161280|T037|PT|945.20|ICD9CM|Blisters, epidermal loss [second degree] of lower limb [leg], unspecified site|Blisters, epidermal loss [second degree] of lower limb [leg], unspecified site
C0161281|T037|AB|945.21|ICD9CM|2nd deg burn toe|2nd deg burn toe
C0161281|T037|PT|945.21|ICD9CM|Blisters, epidermal loss [second degree] of toe(s) (nail)|Blisters, epidermal loss [second degree] of toe(s) (nail)
C0161282|T037|AB|945.22|ICD9CM|2nd deg burn foot|2nd deg burn foot
C0161282|T037|PT|945.22|ICD9CM|Blisters, epidermal loss [second degree] of foot|Blisters, epidermal loss [second degree] of foot
C0161283|T037|AB|945.23|ICD9CM|2nd deg burn ankle|2nd deg burn ankle
C0161283|T037|PT|945.23|ICD9CM|Blisters, epidermal loss [second degree] of ankle|Blisters, epidermal loss [second degree] of ankle
C0161284|T037|AB|945.24|ICD9CM|2nd deg burn lower leg|2nd deg burn lower leg
C0161284|T037|PT|945.24|ICD9CM|Blisters, epidermal loss [second degree] of lower leg|Blisters, epidermal loss [second degree] of lower leg
C0161285|T037|AB|945.25|ICD9CM|2nd deg burn knee|2nd deg burn knee
C0161285|T037|PT|945.25|ICD9CM|Blisters, epidermal loss [second degree] of knee|Blisters, epidermal loss [second degree] of knee
C0161286|T037|AB|945.26|ICD9CM|2nd deg burn thigh|2nd deg burn thigh
C0161286|T037|PT|945.26|ICD9CM|Blisters, epidermal loss [second degree] of thigh [any part]|Blisters, epidermal loss [second degree] of thigh [any part]
C0161287|T037|AB|945.29|ICD9CM|2nd deg burn leg-mult|2nd deg burn leg-mult
C0161287|T037|PT|945.29|ICD9CM|Blisters, epidermal loss [second degree] of multiple sites of lower limb(s)|Blisters, epidermal loss [second degree] of multiple sites of lower limb(s)
C0161288|T037|HT|945.3|ICD9CM|Full-thickness skin loss due to burn [third degree NOS] of lower limb(s)|Full-thickness skin loss due to burn [third degree NOS] of lower limb(s)
C0161289|T037|AB|945.30|ICD9CM|3rd deg burn leg NOS|3rd deg burn leg NOS
C0161289|T037|PT|945.30|ICD9CM|Full-thickness skin loss [third degree NOS] of lower limb [leg] unspecified site|Full-thickness skin loss [third degree NOS] of lower limb [leg] unspecified site
C0161290|T037|AB|945.31|ICD9CM|3rd deg burn toe|3rd deg burn toe
C0161290|T037|PT|945.31|ICD9CM|Full-thickness skin loss [third degree NOS] of toe(s) (nail)|Full-thickness skin loss [third degree NOS] of toe(s) (nail)
C0161291|T037|AB|945.32|ICD9CM|3rd deg burn foot|3rd deg burn foot
C0161291|T037|PT|945.32|ICD9CM|Full-thickness skin loss [third degree NOS] of foot|Full-thickness skin loss [third degree NOS] of foot
C0161292|T037|AB|945.33|ICD9CM|3rd deg burn ankle|3rd deg burn ankle
C0161292|T037|PT|945.33|ICD9CM|Full-thickness skin loss [third degree NOS] of ankle|Full-thickness skin loss [third degree NOS] of ankle
C0161293|T037|AB|945.34|ICD9CM|3rd deg burn low leg|3rd deg burn low leg
C0161293|T037|PT|945.34|ICD9CM|Full-thickness skin loss [third degree nos] of lower leg|Full-thickness skin loss [third degree nos] of lower leg
C0161294|T037|AB|945.35|ICD9CM|3rd deg burn knee|3rd deg burn knee
C0161294|T037|PT|945.35|ICD9CM|Full-thickness skin loss [third degree NOS] of knee|Full-thickness skin loss [third degree NOS] of knee
C0161295|T037|AB|945.36|ICD9CM|3rd deg burn thigh|3rd deg burn thigh
C0161295|T037|PT|945.36|ICD9CM|Full-thickness skin loss [third degree NOS] of thigh [any part]|Full-thickness skin loss [third degree NOS] of thigh [any part]
C0161296|T037|AB|945.39|ICD9CM|3rd deg burn leg-mult|3rd deg burn leg-mult
C0161296|T037|PT|945.39|ICD9CM|Full-thickness skin loss [third degree NOS] of multiple sites of lower limb(s)|Full-thickness skin loss [third degree NOS] of multiple sites of lower limb(s)
C0161298|T037|AB|945.40|ICD9CM|Deep 3rd deg brn leg NOS|Deep 3rd deg brn leg NOS
C0375683|T037|AB|945.41|ICD9CM|Deep 3rd deg burn toe|Deep 3rd deg burn toe
C0161300|T037|AB|945.42|ICD9CM|Deep 3rd deg burn foot|Deep 3rd deg burn foot
C0161301|T037|AB|945.43|ICD9CM|Deep 3rd deg burn ankle|Deep 3rd deg burn ankle
C0161302|T037|AB|945.44|ICD9CM|Deep 3rd deg brn low leg|Deep 3rd deg brn low leg
C0161303|T037|AB|945.45|ICD9CM|Deep 3rd deg burn knee|Deep 3rd deg burn knee
C0161304|T037|AB|945.46|ICD9CM|Deep 3rd deg burn thigh|Deep 3rd deg burn thigh
C0161305|T037|AB|945.49|ICD9CM|Deep 3 deg burn leg-mult|Deep 3 deg burn leg-mult
C0161307|T037|AB|945.50|ICD9CM|3 deg brn w loss-leg NOS|3 deg brn w loss-leg NOS
C0375684|T037|AB|945.51|ICD9CM|3 deg burn w loss-toe|3 deg burn w loss-toe
C0375684|T037|PT|945.51|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of toe(s) (nail)|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of toe(s) (nail)
C0161309|T037|AB|945.52|ICD9CM|3 deg burn w loss-foot|3 deg burn w loss-foot
C0161309|T037|PT|945.52|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of foot|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of foot
C0161310|T037|AB|945.53|ICD9CM|3 deg burn w loss-ankle|3 deg burn w loss-ankle
C0161310|T037|PT|945.53|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of ankle|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of ankle
C0161311|T037|AB|945.54|ICD9CM|3 deg brn w loss-low leg|3 deg brn w loss-low leg
C0161311|T037|PT|945.54|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of lower leg|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of lower leg
C0161312|T037|AB|945.55|ICD9CM|3 deg burn w loss-knee|3 deg burn w loss-knee
C0161312|T037|PT|945.55|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of knee|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of knee
C0161313|T037|AB|945.56|ICD9CM|3 deg burn w loss-thigh|3 deg burn w loss-thigh
C0161314|T037|AB|945.59|ICD9CM|3 deg brn w loss leg-mlt|3 deg brn w loss leg-mlt
C3665447|T037|HT|946|ICD9CM|Burns of multiple specified sites|Burns of multiple specified sites
C1812616|T037|AB|946.0|ICD9CM|Burn NOS multiple site|Burn NOS multiple site
C1812616|T037|PT|946.0|ICD9CM|Burns of multiple specified sites, unspecified degree|Burns of multiple specified sites, unspecified degree
C0161316|T037|AB|946.1|ICD9CM|1st deg burn mult site|1st deg burn mult site
C0161316|T037|PT|946.1|ICD9CM|Erythema [first degree] of multiple specified sites|Erythema [first degree] of multiple specified sites
C0161317|T037|AB|946.2|ICD9CM|2nd deg burn mult site|2nd deg burn mult site
C0161317|T037|PT|946.2|ICD9CM|Blisters, epidermal loss [second degree] of multiple specified sites|Blisters, epidermal loss [second degree] of multiple specified sites
C0161318|T037|AB|946.3|ICD9CM|3rd deg burn mult site|3rd deg burn mult site
C0161318|T037|PT|946.3|ICD9CM|Full-thickness skin loss [third degree NOS] of multiple specified sites|Full-thickness skin loss [third degree NOS] of multiple specified sites
C0161319|T037|AB|946.4|ICD9CM|Deep 3 deg brn mult site|Deep 3 deg brn mult site
C0161320|T037|AB|946.5|ICD9CM|3rd brn w loss-mult site|3rd brn w loss-mult site
C0006420|T037|HT|947|ICD9CM|Burn of internal organs|Burn of internal organs
C0161321|T037|AB|947.0|ICD9CM|Burn of mouth & pharynx|Burn of mouth & pharynx
C0161321|T037|PT|947.0|ICD9CM|Burn of mouth and pharynx|Burn of mouth and pharynx
C0161322|T037|AB|947.1|ICD9CM|Burn larynx/trachea/lung|Burn larynx/trachea/lung
C0161322|T037|PT|947.1|ICD9CM|Burn of larynx, trachea, and lung|Burn of larynx, trachea, and lung
C0162286|T037|AB|947.2|ICD9CM|Burn of esophagus|Burn of esophagus
C0162286|T037|PT|947.2|ICD9CM|Burn of esophagus|Burn of esophagus
C0161323|T037|PT|947.3|ICD9CM|Burn of gastrointestinal tract|Burn of gastrointestinal tract
C0161323|T037|AB|947.3|ICD9CM|Burn of GI tract|Burn of GI tract
C0433217|T037|AB|947.4|ICD9CM|Burn of vagina & uterus|Burn of vagina & uterus
C0433217|T037|PT|947.4|ICD9CM|Burn of vagina and uterus|Burn of vagina and uterus
C0161325|T037|AB|947.8|ICD9CM|Burn internal organ NEC|Burn internal organ NEC
C0161325|T037|PT|947.8|ICD9CM|Burn of other specified sites of internal organs|Burn of other specified sites of internal organs
C0006420|T037|AB|947.9|ICD9CM|Burn internal organ NOS|Burn internal organ NOS
C0006420|T037|PT|947.9|ICD9CM|Burn of internal organs, unspecified site|Burn of internal organs, unspecified site
C0433219|T037|HT|948|ICD9CM|Burns classified according to extent of body surface involved|Burns classified according to extent of body surface involved
C0161327|T037|HT|948.0|ICD9CM|Burn [any degree] involving less than 10 percent of body surface|Burn [any degree] involving less than 10 percent of body surface
C0161328|T037|AB|948.00|ICD9CM|Bdy brn < 10%/3d deg NOS|Bdy brn < 10%/3d deg NOS
C0161329|T037|HT|948.1|ICD9CM|Burn [any degree] involving 10-19 percent of body surface|Burn [any degree] involving 10-19 percent of body surface
C0161330|T037|AB|948.10|ICD9CM|10-19% bdy brn/3 deg NOS|10-19% bdy brn/3 deg NOS
C0161331|T037|AB|948.11|ICD9CM|10-19% bdy brn/10-19% 3d|10-19% bdy brn/10-19% 3d
C0161331|T037|PT|948.11|ICD9CM|Burn [any degree] involving 10-19 percent of body surface with third degree burn, 10-19%|Burn [any degree] involving 10-19 percent of body surface with third degree burn, 10-19%
C0161332|T037|HT|948.2|ICD9CM|Burn [any degree] involving 20-29 percent of body surface|Burn [any degree] involving 20-29 percent of body surface
C0161333|T037|AB|948.20|ICD9CM|20-29% bdy brn/3 deg NOS|20-29% bdy brn/3 deg NOS
C0161334|T037|AB|948.21|ICD9CM|20-29% bdy brn/10-19% 3d|20-29% bdy brn/10-19% 3d
C0161334|T037|PT|948.21|ICD9CM|Burn [any degree] involving 20-29 percent of body surface with third degree burn, 10-19%|Burn [any degree] involving 20-29 percent of body surface with third degree burn, 10-19%
C0161335|T037|AB|948.22|ICD9CM|20-29% bdy brn/20-29% 3d|20-29% bdy brn/20-29% 3d
C0161335|T037|PT|948.22|ICD9CM|Burn [any degree] involving 20-29 percent of body surface with third degree burn, 20-29%|Burn [any degree] involving 20-29 percent of body surface with third degree burn, 20-29%
C0161336|T037|HT|948.3|ICD9CM|Burn [any degree] involving 30-39 percent of body surface|Burn [any degree] involving 30-39 percent of body surface
C0161337|T037|AB|948.30|ICD9CM|30-39% bdy brn/3 deg NOS|30-39% bdy brn/3 deg NOS
C0161338|T037|AB|948.31|ICD9CM|30-39% bdy brn/10-19% 3d|30-39% bdy brn/10-19% 3d
C0161338|T037|PT|948.31|ICD9CM|Burn [any degree] involving 30-39 percent of body surface with third degree burn, 10-19%|Burn [any degree] involving 30-39 percent of body surface with third degree burn, 10-19%
C0161339|T037|AB|948.32|ICD9CM|30-39% bdy brn/20-29% 3d|30-39% bdy brn/20-29% 3d
C0161339|T037|PT|948.32|ICD9CM|Burn [any degree] involving 30-39 percent of body surface with third degree burn, 20-29%|Burn [any degree] involving 30-39 percent of body surface with third degree burn, 20-29%
C0161340|T037|AB|948.33|ICD9CM|30-39% bdy brn/30-39% 3d|30-39% bdy brn/30-39% 3d
C0161340|T037|PT|948.33|ICD9CM|Burn [any degree] involving 30-39 percent of body surface with third degree burn, 30-39%|Burn [any degree] involving 30-39 percent of body surface with third degree burn, 30-39%
C0161341|T037|HT|948.4|ICD9CM|Burn [any degree] involving 40-49 percent of body surface|Burn [any degree] involving 40-49 percent of body surface
C0161342|T037|AB|948.40|ICD9CM|40-49% bdy brn/3 deg NOS|40-49% bdy brn/3 deg NOS
C0161343|T037|AB|948.41|ICD9CM|40-49% bdy brn/10-19% 3d|40-49% bdy brn/10-19% 3d
C0161343|T037|PT|948.41|ICD9CM|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 10-19%|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 10-19%
C0161344|T037|AB|948.42|ICD9CM|40-49% bdy brn/20-29% 3d|40-49% bdy brn/20-29% 3d
C0161344|T037|PT|948.42|ICD9CM|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 20-29%|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 20-29%
C0161345|T037|AB|948.43|ICD9CM|40-49% bdy brn/30-39% 3d|40-49% bdy brn/30-39% 3d
C0161345|T037|PT|948.43|ICD9CM|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 30-39%|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 30-39%
C0161346|T037|AB|948.44|ICD9CM|40-49% bdy brn/40-49% 3d|40-49% bdy brn/40-49% 3d
C0161346|T037|PT|948.44|ICD9CM|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 40-49%|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 40-49%
C0161347|T037|HT|948.5|ICD9CM|Burn [any degree] involving 50-59 percent of body surface|Burn [any degree] involving 50-59 percent of body surface
C0161348|T037|AB|948.50|ICD9CM|50-59% bdy brn/3 deg NOS|50-59% bdy brn/3 deg NOS
C0161349|T037|AB|948.51|ICD9CM|50-59% bdy brn/10-19% 3d|50-59% bdy brn/10-19% 3d
C0161349|T037|PT|948.51|ICD9CM|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 10-19%|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 10-19%
C0161350|T037|AB|948.52|ICD9CM|50-59% bdy brn/20-29% 3d|50-59% bdy brn/20-29% 3d
C0161350|T037|PT|948.52|ICD9CM|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 20-29%|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 20-29%
C0161351|T037|AB|948.53|ICD9CM|50-59% bdy brn/30-39% 3d|50-59% bdy brn/30-39% 3d
C0161351|T037|PT|948.53|ICD9CM|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 30-39%|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 30-39%
C0161352|T037|AB|948.54|ICD9CM|50-59% bdy brn/40-49% 3d|50-59% bdy brn/40-49% 3d
C0161352|T037|PT|948.54|ICD9CM|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 40-49%|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 40-49%
C0161353|T037|AB|948.55|ICD9CM|50-59% bdy brn/50-59% 3d|50-59% bdy brn/50-59% 3d
C0161353|T037|PT|948.55|ICD9CM|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 50-59%|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 50-59%
C0161354|T037|HT|948.6|ICD9CM|Burn [any degree] involving 60-69 percent of body surface|Burn [any degree] involving 60-69 percent of body surface
C0161355|T037|AB|948.60|ICD9CM|60-69% bdy brn/3 deg NOS|60-69% bdy brn/3 deg NOS
C0161356|T037|AB|948.61|ICD9CM|60-69% bdy brn/10-19% 3d|60-69% bdy brn/10-19% 3d
C0161356|T037|PT|948.61|ICD9CM|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 10-19%|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 10-19%
C0161357|T037|AB|948.62|ICD9CM|60-69% bdy brn/20-29% 3d|60-69% bdy brn/20-29% 3d
C0161357|T037|PT|948.62|ICD9CM|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 20-29%|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 20-29%
C0161358|T037|AB|948.63|ICD9CM|60-69% bdy brn/30-39% 3d|60-69% bdy brn/30-39% 3d
C0161358|T037|PT|948.63|ICD9CM|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 30-39%|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 30-39%
C0161359|T037|AB|948.64|ICD9CM|60-69% bdy brn/40-49% 3d|60-69% bdy brn/40-49% 3d
C0161359|T037|PT|948.64|ICD9CM|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 40-49%|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 40-49%
C0161360|T037|AB|948.65|ICD9CM|60-69% bdy brn/50-59% 3d|60-69% bdy brn/50-59% 3d
C0161360|T037|PT|948.65|ICD9CM|Burn (any degree) involving 60-69 percent of body surface with third degree burn, 50-59%|Burn (any degree) involving 60-69 percent of body surface with third degree burn, 50-59%
C0161361|T037|AB|948.66|ICD9CM|60-69% bdy brn/60-69% 3d|60-69% bdy brn/60-69% 3d
C0161361|T037|PT|948.66|ICD9CM|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 60-69%|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 60-69%
C0161362|T037|HT|948.7|ICD9CM|Burn [any degree] involving 70-79 percent of body surface|Burn [any degree] involving 70-79 percent of body surface
C0161363|T037|AB|948.70|ICD9CM|70-79% bdy brn/3 deg NOS|70-79% bdy brn/3 deg NOS
C0161364|T037|AB|948.71|ICD9CM|70-79% bdy brn/10-19% 3d|70-79% bdy brn/10-19% 3d
C0161364|T037|PT|948.71|ICD9CM|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 10-19%|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 10-19%
C0161365|T037|AB|948.72|ICD9CM|70-79% bdy brn/20-29% 3d|70-79% bdy brn/20-29% 3d
C0161365|T037|PT|948.72|ICD9CM|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 20-29%|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 20-29%
C0161366|T037|AB|948.73|ICD9CM|70-79% bdy brn/30-39% 3d|70-79% bdy brn/30-39% 3d
C0161366|T037|PT|948.73|ICD9CM|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 30-39%|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 30-39%
C0161367|T037|AB|948.74|ICD9CM|70-79% bdy brn/40-49% 3d|70-79% bdy brn/40-49% 3d
C0161367|T037|PT|948.74|ICD9CM|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 40-49%|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 40-49%
C0161368|T037|AB|948.75|ICD9CM|70-79% bdy brn/50-59% 3d|70-79% bdy brn/50-59% 3d
C0161368|T037|PT|948.75|ICD9CM|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 50-59%|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 50-59%
C0161369|T037|AB|948.76|ICD9CM|70-79% bdy brn/60-69% 3d|70-79% bdy brn/60-69% 3d
C0161369|T037|PT|948.76|ICD9CM|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 60-69%|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 60-69%
C0161370|T037|AB|948.77|ICD9CM|70-79% bdy brn/70-79% 3d|70-79% bdy brn/70-79% 3d
C0161370|T037|PT|948.77|ICD9CM|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 70-79%|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 70-79%
C0161371|T037|HT|948.8|ICD9CM|Burn [any degree] involving 80-89 percent of body surface|Burn [any degree] involving 80-89 percent of body surface
C0161372|T037|AB|948.80|ICD9CM|80-89% bdy brn/3 deg NOS|80-89% bdy brn/3 deg NOS
C0161373|T037|AB|948.81|ICD9CM|80-89% bdy brn/10-19% 3d|80-89% bdy brn/10-19% 3d
C0161373|T037|PT|948.81|ICD9CM|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 10-19%|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 10-19%
C0161374|T037|AB|948.82|ICD9CM|80-89% bdy brn/20-29% 3d|80-89% bdy brn/20-29% 3d
C0161374|T037|PT|948.82|ICD9CM|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 20-29%|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 20-29%
C0161375|T037|AB|948.83|ICD9CM|80-89% bdy brn/30-39% 3d|80-89% bdy brn/30-39% 3d
C0161375|T037|PT|948.83|ICD9CM|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 30-39%|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 30-39%
C0161376|T037|AB|948.84|ICD9CM|80-89% bdy brn/40-49% 3d|80-89% bdy brn/40-49% 3d
C0161376|T037|PT|948.84|ICD9CM|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 40-49%|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 40-49%
C0161377|T037|AB|948.85|ICD9CM|80-89% bdy brn/50-59% 3d|80-89% bdy brn/50-59% 3d
C0161377|T037|PT|948.85|ICD9CM|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 50-59%|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 50-59%
C0161378|T037|AB|948.86|ICD9CM|80-89% bdy brn/60-69% 3d|80-89% bdy brn/60-69% 3d
C0161378|T037|PT|948.86|ICD9CM|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 60-69%|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 60-69%
C0161379|T037|AB|948.87|ICD9CM|80-89% bdy brn/70-79% 3d|80-89% bdy brn/70-79% 3d
C0161379|T037|PT|948.87|ICD9CM|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 70-79%|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 70-79%
C0161380|T037|AB|948.88|ICD9CM|80-89% bdy brn/80-89% 3d|80-89% bdy brn/80-89% 3d
C0161380|T037|PT|948.88|ICD9CM|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 80-89%|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 80-89%
C0161381|T037|HT|948.9|ICD9CM|Burn [any degree] involving 90 percent or more of body surface|Burn [any degree] involving 90 percent or more of body surface
C0161382|T037|AB|948.90|ICD9CM|90% + bdy brn/3d deg NOS|90% + bdy brn/3d deg NOS
C0161383|T037|AB|948.91|ICD9CM|90% + bdy brn/10-19% 3rd|90% + bdy brn/10-19% 3rd
C0161383|T037|PT|948.91|ICD9CM|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 10-19%|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 10-19%
C0161384|T037|AB|948.92|ICD9CM|90% + bdy brn/20-29% 3rd|90% + bdy brn/20-29% 3rd
C0161384|T037|PT|948.92|ICD9CM|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 20-29%|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 20-29%
C0161385|T037|AB|948.93|ICD9CM|90% + bdy brn/30-39% 3rd|90% + bdy brn/30-39% 3rd
C0161385|T037|PT|948.93|ICD9CM|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 30-39%|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 30-39%
C0161386|T037|AB|948.94|ICD9CM|90% + bdy brn/40-49% 3rd|90% + bdy brn/40-49% 3rd
C0161386|T037|PT|948.94|ICD9CM|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 40-49%|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 40-49%
C0161387|T037|AB|948.95|ICD9CM|90% + bdy brn/50-59% 3rd|90% + bdy brn/50-59% 3rd
C0161387|T037|PT|948.95|ICD9CM|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 50-59%|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 50-59%
C0161388|T037|AB|948.96|ICD9CM|90% + bdy brn/60-69% 3rd|90% + bdy brn/60-69% 3rd
C0161388|T037|PT|948.96|ICD9CM|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 60-69%|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 60-69%
C0161389|T037|AB|948.97|ICD9CM|90% + bdy brn/70-79% 3rd|90% + bdy brn/70-79% 3rd
C0161389|T037|PT|948.97|ICD9CM|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 70-79%|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 70-79%
C0161390|T037|AB|948.98|ICD9CM|90% + bdy brn/80-89% 3rd|90% + bdy brn/80-89% 3rd
C0161390|T037|PT|948.98|ICD9CM|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 80-89%|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 80-89%
C0161391|T037|AB|948.99|ICD9CM|90% + bdy brn/90% + 3rd|90% + bdy brn/90% + 3rd
C1812606|T037|HT|949|ICD9CM|Burn, unspecified site|Burn, unspecified site
C0006434|T037|AB|949.0|ICD9CM|Burn NOS|Burn NOS
C0006434|T037|PT|949.0|ICD9CM|Burn of unspecified site, unspecified degree|Burn of unspecified site, unspecified degree
C0332686|T037|AB|949.1|ICD9CM|1st degree burn NOS|1st degree burn NOS
C0332686|T037|PT|949.1|ICD9CM|Erythema [first degree], unspecified site|Erythema [first degree], unspecified site
C0332687|T037|AB|949.2|ICD9CM|2nd degree burn NOS|2nd degree burn NOS
C0332687|T037|PT|949.2|ICD9CM|Blisters, epidermal loss [second degree], unspecified site|Blisters, epidermal loss [second degree], unspecified site
C0375688|T037|AB|949.3|ICD9CM|3rd degree burn NOS|3rd degree burn NOS
C0375688|T037|PT|949.3|ICD9CM|Full-thickness skin loss [third degree nos]|Full-thickness skin loss [third degree nos]
C0161395|T037|AB|949.4|ICD9CM|Deep 3rd deg burn NOS|Deep 3rd deg burn NOS
C0161396|T037|AB|949.5|ICD9CM|3rd burn w loss-site NOS|3rd burn w loss-site NOS
C0161396|T037|PT|949.5|ICD9CM|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, unspecified|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, unspecified
C0161397|T037|HT|950|ICD9CM|Injury to optic nerve and pathways|Injury to optic nerve and pathways
C0178330|T037|HT|950-957.99|ICD9CM|INJURY TO NERVES AND SPINAL CORD|INJURY TO NERVES AND SPINAL CORD
C0161398|T037|AB|950.0|ICD9CM|Optic nerve injury|Optic nerve injury
C0161398|T037|PT|950.0|ICD9CM|Optic nerve injury|Optic nerve injury
C0161399|T037|AB|950.1|ICD9CM|Injury to optic chiasm|Injury to optic chiasm
C0161399|T037|PT|950.1|ICD9CM|Injury to optic chiasm|Injury to optic chiasm
C0161400|T037|AB|950.2|ICD9CM|Injury to optic pathways|Injury to optic pathways
C0161400|T037|PT|950.2|ICD9CM|Injury to optic pathways|Injury to optic pathways
C0161401|T037|AB|950.3|ICD9CM|Injury to visual cortex|Injury to visual cortex
C0161401|T037|PT|950.3|ICD9CM|Injury to visual cortex|Injury to visual cortex
C0161397|T037|AB|950.9|ICD9CM|Inj optic nerv/path NOS|Inj optic nerv/path NOS
C0161397|T037|PT|950.9|ICD9CM|Injury to unspecified optic nerve and pathways|Injury to unspecified optic nerve and pathways
C0478205|T037|HT|951|ICD9CM|Injury to other cranial nerve(s)|Injury to other cranial nerve(s)
C1321926|T037|AB|951.0|ICD9CM|Injury oculomotor nerve|Injury oculomotor nerve
C1321926|T037|PT|951.0|ICD9CM|Injury to oculomotor nerve|Injury to oculomotor nerve
C0161405|T037|PT|951.1|ICD9CM|Injury to trochlear nerve|Injury to trochlear nerve
C0161405|T037|AB|951.1|ICD9CM|Injury trochlear nerve|Injury trochlear nerve
C0161406|T037|PT|951.2|ICD9CM|Injury to trigeminal nerve|Injury to trigeminal nerve
C0161406|T037|AB|951.2|ICD9CM|Injury trigeminal nerve|Injury trigeminal nerve
C0161407|T037|AB|951.3|ICD9CM|Injury abducens nerve|Injury abducens nerve
C0161407|T037|PT|951.3|ICD9CM|Injury to abducens nerve|Injury to abducens nerve
C0161408|T037|AB|951.4|ICD9CM|Injury to facial nerve|Injury to facial nerve
C0161408|T037|PT|951.4|ICD9CM|Injury to facial nerve|Injury to facial nerve
C0161409|T037|AB|951.5|ICD9CM|Injury to acoustic nerve|Injury to acoustic nerve
C0161409|T037|PT|951.5|ICD9CM|Injury to acoustic nerve|Injury to acoustic nerve
C0161410|T037|AB|951.6|ICD9CM|Injury accessory nerve|Injury accessory nerve
C0161410|T037|PT|951.6|ICD9CM|Injury to accessory nerve|Injury to accessory nerve
C0161411|T037|AB|951.7|ICD9CM|Injury hypoglossal nerve|Injury hypoglossal nerve
C0161411|T037|PT|951.7|ICD9CM|Injury to hypoglossal nerve|Injury to hypoglossal nerve
C0161412|T037|AB|951.8|ICD9CM|Injury cranial nerve NEC|Injury cranial nerve NEC
C0161412|T037|PT|951.8|ICD9CM|Injury to other specified cranial nerves|Injury to other specified cranial nerves
C0273483|T037|AB|951.9|ICD9CM|Injury cranial nerve NOS|Injury cranial nerve NOS
C0273483|T037|PT|951.9|ICD9CM|Injury to unspecified cranial nerve|Injury to unspecified cranial nerve
C0161414|T037|HT|952|ICD9CM|Spinal cord injury without evidence of spinal bone injury|Spinal cord injury without evidence of spinal bone injury
C0433858|T037|HT|952.0|ICD9CM|Cervical spinal cord injury without evidence of spinal bone injury|Cervical spinal cord injury without evidence of spinal bone injury
C0161416|T037|PT|952.00|ICD9CM|C1-C4 level with unspecified spinal cord injury|C1-C4 level with unspecified spinal cord injury
C0161416|T037|AB|952.00|ICD9CM|C1-c4 spin cord inj NOS|C1-c4 spin cord inj NOS
C0161417|T037|PT|952.01|ICD9CM|C1-C4 level with complete lesion of spinal cord|C1-C4 level with complete lesion of spinal cord
C0161417|T037|AB|952.01|ICD9CM|Complete les cord/c1-c4|Complete les cord/c1-c4
C0161418|T037|AB|952.02|ICD9CM|Anterior cord synd/c1-c4|Anterior cord synd/c1-c4
C0161418|T037|PT|952.02|ICD9CM|C1-C4 level with anterior cord syndrome|C1-C4 level with anterior cord syndrome
C0161419|T037|PT|952.03|ICD9CM|C1-C4 level with central cord syndrome|C1-C4 level with central cord syndrome
C0161419|T037|AB|952.03|ICD9CM|Central cord synd/c1-c4|Central cord synd/c1-c4
C0161420|T037|PT|952.04|ICD9CM|C1-C4 level with other specified spinal cord injury|C1-C4 level with other specified spinal cord injury
C0161420|T037|AB|952.04|ICD9CM|C1-c4 spin cord inj NEC|C1-c4 spin cord inj NEC
C0161421|T037|PT|952.05|ICD9CM|C5-C7 level with unspecified spinal cord injury|C5-C7 level with unspecified spinal cord injury
C0161421|T037|AB|952.05|ICD9CM|C5-c7 spin cord inj NOS|C5-c7 spin cord inj NOS
C0161422|T037|PT|952.06|ICD9CM|C5-C7 level with complete lesion of spinal cord|C5-C7 level with complete lesion of spinal cord
C0161422|T037|AB|952.06|ICD9CM|Complete les cord/c5-c7|Complete les cord/c5-c7
C0161423|T037|AB|952.07|ICD9CM|Anterior cord synd/c5-c7|Anterior cord synd/c5-c7
C0161423|T037|PT|952.07|ICD9CM|C5-C7 level with anterior cord syndrome|C5-C7 level with anterior cord syndrome
C0161424|T037|PT|952.08|ICD9CM|C5-C7 level with central cord syndrome|C5-C7 level with central cord syndrome
C0161424|T037|AB|952.08|ICD9CM|Central cord synd/c5-c7|Central cord synd/c5-c7
C0161425|T037|PT|952.09|ICD9CM|C5-C7 level with other specified spinal cord injury|C5-C7 level with other specified spinal cord injury
C0161425|T037|AB|952.09|ICD9CM|C5-c7 spin cord inj NEC|C5-c7 spin cord inj NEC
C0161426|T037|HT|952.1|ICD9CM|Dorsal [thoracic] spinal cord injury without evidence of spinal bone injury|Dorsal [thoracic] spinal cord injury without evidence of spinal bone injury
C0161427|T037|PT|952.10|ICD9CM|T1-T6 level with unspecified spinal cord injury|T1-T6 level with unspecified spinal cord injury
C0161427|T037|AB|952.10|ICD9CM|T1-t6 spin cord inj NOS|T1-t6 spin cord inj NOS
C0859375|T037|AB|952.11|ICD9CM|Complete les cord/t1-t6|Complete les cord/t1-t6
C0859375|T037|PT|952.11|ICD9CM|T1-T6 level with complete lesion of spinal cord|T1-T6 level with complete lesion of spinal cord
C0859376|T037|AB|952.12|ICD9CM|Anterior cord synd/t1-t6|Anterior cord synd/t1-t6
C0859376|T037|PT|952.12|ICD9CM|T1-T6 level with anterior cord syndrome|T1-T6 level with anterior cord syndrome
C0859377|T037|AB|952.13|ICD9CM|Central cord synd/t1-t6|Central cord synd/t1-t6
C0859377|T037|PT|952.13|ICD9CM|T1-T6 level with central cord syndrome|T1-T6 level with central cord syndrome
C0859378|T037|PT|952.14|ICD9CM|T1-T6 level with other specified spinal cord injury|T1-T6 level with other specified spinal cord injury
C0859378|T037|AB|952.14|ICD9CM|T1-t6 spin cord inj NEC|T1-t6 spin cord inj NEC
C0161432|T037|PT|952.15|ICD9CM|T7-T12 level with unspecified spinal cord injury|T7-T12 level with unspecified spinal cord injury
C0161432|T037|AB|952.15|ICD9CM|T7-t12 spin cord inj NOS|T7-t12 spin cord inj NOS
C0859379|T037|AB|952.16|ICD9CM|Complete les cord/t7-t12|Complete les cord/t7-t12
C0859379|T037|PT|952.16|ICD9CM|T7-T12 level with complete lesion of spinal cord|T7-T12 level with complete lesion of spinal cord
C0859380|T037|AB|952.17|ICD9CM|Anterior cord syn/t7-t12|Anterior cord syn/t7-t12
C0859380|T037|PT|952.17|ICD9CM|T7-T12 level with anterior cord syndrome|T7-T12 level with anterior cord syndrome
C0859381|T037|AB|952.18|ICD9CM|Central cord syn/t7-t12|Central cord syn/t7-t12
C0859381|T037|PT|952.18|ICD9CM|T7-T12 level with central cord syndrome|T7-T12 level with central cord syndrome
C0161436|T037|PT|952.19|ICD9CM|T7-T12 level with other specified spinal cord injury|T7-T12 level with other specified spinal cord injury
C0161436|T037|AB|952.19|ICD9CM|T7-t12 spin cord inj NEC|T7-t12 spin cord inj NEC
C0273520|T037|AB|952.2|ICD9CM|Lumbar spinal cord injur|Lumbar spinal cord injur
C0273520|T037|PT|952.2|ICD9CM|Lumbar spinal cord injury without evidence of spinal bone injury|Lumbar spinal cord injury without evidence of spinal bone injury
C0273521|T037|AB|952.3|ICD9CM|Sacral spinal cord injur|Sacral spinal cord injur
C0273521|T037|PT|952.3|ICD9CM|Sacral spinal cord injury without evidence of spinal bone injury|Sacral spinal cord injury without evidence of spinal bone injury
C0161439|T037|AB|952.4|ICD9CM|Cauda equina injury|Cauda equina injury
C0161439|T037|PT|952.4|ICD9CM|Cauda equina spinal cord injury without evidence of spinal bone injury|Cauda equina spinal cord injury without evidence of spinal bone injury
C0161440|T037|PT|952.8|ICD9CM|Multiple sites of spinal cord injury without evidence of spinal bone injury|Multiple sites of spinal cord injury without evidence of spinal bone injury
C0161440|T037|AB|952.8|ICD9CM|Spin cord inj-mult site|Spin cord inj-mult site
C0859273|T037|AB|952.9|ICD9CM|Spinal cord injury NOS|Spinal cord injury NOS
C0859273|T037|PT|952.9|ICD9CM|Unspecified site of spinal cord injury without evidence of spinal bone injury|Unspecified site of spinal cord injury without evidence of spinal bone injury
C0161441|T037|HT|953|ICD9CM|Injury to nerve roots and spinal plexus|Injury to nerve roots and spinal plexus
C0161442|T037|AB|953.0|ICD9CM|Cervical root injury|Cervical root injury
C0161442|T037|PT|953.0|ICD9CM|Injury to cervical nerve root|Injury to cervical nerve root
C1536686|T037|AB|953.1|ICD9CM|Dorsal root injury|Dorsal root injury
C1536686|T037|PT|953.1|ICD9CM|Injury to dorsal nerve root|Injury to dorsal nerve root
C0161444|T037|PT|953.2|ICD9CM|Injury to lumbar nerve root|Injury to lumbar nerve root
C0161444|T037|AB|953.2|ICD9CM|Lumbar root injury|Lumbar root injury
C0161445|T037|PT|953.3|ICD9CM|Injury to sacral nerve root|Injury to sacral nerve root
C0161445|T037|AB|953.3|ICD9CM|Sacral root injury|Sacral root injury
C0161446|T037|AB|953.4|ICD9CM|Brachial plexus injury|Brachial plexus injury
C0161446|T037|PT|953.4|ICD9CM|Injury to brachial plexus|Injury to brachial plexus
C0161447|T037|PT|953.5|ICD9CM|Injury to lumbosacral plexus|Injury to lumbosacral plexus
C0161447|T037|AB|953.5|ICD9CM|Lumbosacral plex injury|Lumbosacral plex injury
C0161448|T037|PT|953.8|ICD9CM|Injury to multiple sites of nerve roots and spinal plexus|Injury to multiple sites of nerve roots and spinal plexus
C0161448|T037|AB|953.8|ICD9CM|Mult nerve root/plex inj|Mult nerve root/plex inj
C0161441|T037|AB|953.9|ICD9CM|Inj nerve root/plex NOS|Inj nerve root/plex NOS
C0161441|T037|PT|953.9|ICD9CM|Injury to unspecified site of nerve roots and spinal plexus|Injury to unspecified site of nerve roots and spinal plexus
C0433857|T037|HT|954|ICD9CM|Injury to other nerve(s) of trunk, excluding shoulder and pelvic girdles|Injury to other nerve(s) of trunk, excluding shoulder and pelvic girdles
C0161451|T037|AB|954.0|ICD9CM|Inj cerv sympath nerve|Inj cerv sympath nerve
C0161451|T037|PT|954.0|ICD9CM|Injury to cervical sympathetic nerve, excluding shoulder and pelvic girdles|Injury to cervical sympathetic nerve, excluding shoulder and pelvic girdles
C0161452|T037|AB|954.1|ICD9CM|Inj sympath nerve NEC|Inj sympath nerve NEC
C0161452|T037|PT|954.1|ICD9CM|Injury to other sympathetic nerve, excluding shoulder and pelvic girdles|Injury to other sympathetic nerve, excluding shoulder and pelvic girdles
C0161453|T037|PT|954.8|ICD9CM|Injury to other specified nerve(s) of trunk, excluding shoulder and pelvic girdles|Injury to other specified nerve(s) of trunk, excluding shoulder and pelvic girdles
C0161453|T037|AB|954.8|ICD9CM|Injury trunk nerve NEC|Injury trunk nerve NEC
C0161454|T037|PT|954.9|ICD9CM|Injury to unspecified nerve of trunk, excluding shoulder and pelvic girdles|Injury to unspecified nerve of trunk, excluding shoulder and pelvic girdles
C0161454|T037|AB|954.9|ICD9CM|Injury trunk nerve NOS|Injury trunk nerve NOS
C0273529|T037|HT|955|ICD9CM|Injury to peripheral nerve(s) of shoulder girdle and upper limb|Injury to peripheral nerve(s) of shoulder girdle and upper limb
C0161456|T037|AB|955.0|ICD9CM|Injury axillary nerve|Injury axillary nerve
C0161456|T037|PT|955.0|ICD9CM|Injury to axillary nerve|Injury to axillary nerve
C0161457|T037|AB|955.1|ICD9CM|Injury median nerve|Injury median nerve
C0161457|T037|PT|955.1|ICD9CM|Injury to median nerve|Injury to median nerve
C0161458|T037|PT|955.2|ICD9CM|Injury to ulnar nerve|Injury to ulnar nerve
C0161458|T037|AB|955.2|ICD9CM|Injury ulnar nerve|Injury ulnar nerve
C0161459|T037|AB|955.3|ICD9CM|Injury radial nerve|Injury radial nerve
C0161459|T037|PT|955.3|ICD9CM|Injury to radial nerve|Injury to radial nerve
C0161460|T037|AB|955.4|ICD9CM|Inj musculocutan nerve|Inj musculocutan nerve
C0161460|T037|PT|955.4|ICD9CM|Injury to musculocutaneous nerve|Injury to musculocutaneous nerve
C0161461|T037|AB|955.5|ICD9CM|Inj cutan senso nerv/arm|Inj cutan senso nerv/arm
C0161461|T037|PT|955.5|ICD9CM|Injury to cutaneous sensory nerve, upper limb|Injury to cutaneous sensory nerve, upper limb
C0161462|T037|AB|955.6|ICD9CM|Injury digital nerve|Injury digital nerve
C0161462|T037|PT|955.6|ICD9CM|Injury to digital nerve, upper limb|Injury to digital nerve, upper limb
C0161463|T037|AB|955.7|ICD9CM|Inj nerve shldr/arm NEC|Inj nerve shldr/arm NEC
C0161463|T037|PT|955.7|ICD9CM|Injury to other specified nerve(s) of shoulder girdle and upper limb|Injury to other specified nerve(s) of shoulder girdle and upper limb
C2053768|T037|AB|955.8|ICD9CM|Inj mult nerve shldr/arm|Inj mult nerve shldr/arm
C2053768|T037|PT|955.8|ICD9CM|Injury to multiple nerves of shoulder girdle and upper limb|Injury to multiple nerves of shoulder girdle and upper limb
C0273529|T037|AB|955.9|ICD9CM|Inj nerve shldr/arm NOS|Inj nerve shldr/arm NOS
C0273529|T037|PT|955.9|ICD9CM|Injury to unspecified nerve of shoulder girdle and upper limb|Injury to unspecified nerve of shoulder girdle and upper limb
C1260908|T037|HT|956|ICD9CM|Injury to peripheral nerve(s) of pelvic girdle and lower limb|Injury to peripheral nerve(s) of pelvic girdle and lower limb
C0161467|T037|AB|956.0|ICD9CM|Injury sciatic nerve|Injury sciatic nerve
C0161467|T037|PT|956.0|ICD9CM|Injury to sciatic nerve|Injury to sciatic nerve
C0161468|T037|AB|956.1|ICD9CM|Injury femoral nerve|Injury femoral nerve
C0161468|T037|PT|956.1|ICD9CM|Injury to femoral nerve|Injury to femoral nerve
C0273532|T037|AB|956.2|ICD9CM|Inj posterior tib nerve|Inj posterior tib nerve
C0273532|T037|PT|956.2|ICD9CM|Injury to posterior tibial nerve|Injury to posterior tibial nerve
C1321896|T037|AB|956.3|ICD9CM|Injury peroneal nerve|Injury peroneal nerve
C1321896|T037|PT|956.3|ICD9CM|Injury to peroneal nerve|Injury to peroneal nerve
C0161471|T037|AB|956.4|ICD9CM|Inj cutan senso nerv/leg|Inj cutan senso nerv/leg
C0161471|T037|PT|956.4|ICD9CM|Injury to cutaneous sensory nerve, lower limb|Injury to cutaneous sensory nerve, lower limb
C0273533|T037|AB|956.5|ICD9CM|Inj nerve pelv/leg NEC|Inj nerve pelv/leg NEC
C0273533|T037|PT|956.5|ICD9CM|Injury to other specified nerve(s) of pelvic girdle and lower limb|Injury to other specified nerve(s) of pelvic girdle and lower limb
C0161473|T037|AB|956.8|ICD9CM|Inj mult nerve pelv/leg|Inj mult nerve pelv/leg
C0161473|T037|PT|956.8|ICD9CM|Injury to multiple nerves of pelvic girdle and lower limb|Injury to multiple nerves of pelvic girdle and lower limb
C0273531|T037|AB|956.9|ICD9CM|Inj nerve pelv/leg NOS|Inj nerve pelv/leg NOS
C0273531|T037|PT|956.9|ICD9CM|Injury to unspecified nerve of pelvic girdle and lower limb|Injury to unspecified nerve of pelvic girdle and lower limb
C0161475|T037|HT|957|ICD9CM|Injury to other and unspecified nerves|Injury to other and unspecified nerves
C0161476|T037|AB|957.0|ICD9CM|Inj superf nerv head/nck|Inj superf nerv head/nck
C0161476|T037|PT|957.0|ICD9CM|Injury to superficial nerves of head and neck|Injury to superficial nerves of head and neck
C0434291|T037|AB|957.1|ICD9CM|Injury to nerve NEC|Injury to nerve NEC
C0434291|T037|PT|957.1|ICD9CM|Injury to other specified nerve(s)|Injury to other specified nerve(s)
C0161478|T037|AB|957.8|ICD9CM|Injury to mult nerves|Injury to mult nerves
C0161478|T037|PT|957.8|ICD9CM|Injury to multiple nerves in several parts|Injury to multiple nerves in several parts
C0161479|T037|AB|957.9|ICD9CM|Injury to nerve NOS|Injury to nerve NOS
C0161479|T037|PT|957.9|ICD9CM|Injury to nerves, unspecified site|Injury to nerves, unspecified site
C0161480|T046|HT|958|ICD9CM|Certain early complications of trauma|Certain early complications of trauma
C0178331|T037|HT|958-959.99|ICD9CM|CERTAIN TRAUMATIC COMPLICATIONS AND UNSPECIFIED INJURIES|CERTAIN TRAUMATIC COMPLICATIONS AND UNSPECIFIED INJURIES
C0274265|T037|AB|958.0|ICD9CM|Air embolism|Air embolism
C0274265|T037|PT|958.0|ICD9CM|Air embolism|Air embolism
C1533618|T046|AB|958.1|ICD9CM|Fat embolism|Fat embolism
C1533618|T046|PT|958.1|ICD9CM|Fat embolism|Fat embolism
C0274267|T046|PT|958.2|ICD9CM|Secondary and recurrent hemorrhage|Secondary and recurrent hemorrhage
C0274267|T046|AB|958.2|ICD9CM|Secondary/recur hemorr|Secondary/recur hemorr
C0868767|T047|AB|958.3|ICD9CM|Posttraum wnd infec NEC|Posttraum wnd infec NEC
C0868767|T047|PT|958.3|ICD9CM|Posttraumatic wound infection not elsewhere classified|Posttraumatic wound infection not elsewhere classified
C0036986|T046|AB|958.4|ICD9CM|Traumatic shock|Traumatic shock
C0036986|T046|PT|958.4|ICD9CM|Traumatic shock|Traumatic shock
C0040793|T037|AB|958.5|ICD9CM|Traumatic anuria|Traumatic anuria
C0040793|T037|PT|958.5|ICD9CM|Traumatic anuria|Traumatic anuria
C0042951|T047|AB|958.6|ICD9CM|Volkmann's isch contract|Volkmann's isch contract
C0042951|T047|PT|958.6|ICD9CM|Volkmann's ischemic contracture|Volkmann's ischemic contracture
C0040799|T037|AB|958.7|ICD9CM|Traum subcutan emphysema|Traum subcutan emphysema
C0040799|T037|PT|958.7|ICD9CM|Traumatic subcutaneous emphysema|Traumatic subcutaneous emphysema
C0029603|T037|AB|958.8|ICD9CM|Early complic trauma NEC|Early complic trauma NEC
C0029603|T037|PT|958.8|ICD9CM|Other early complications of trauma|Other early complications of trauma
C1719662|T037|HT|958.9|ICD9CM|Traumatic compartment syndrome|Traumatic compartment syndrome
C0009492|T047|AB|958.90|ICD9CM|Compartment syndrome NOS|Compartment syndrome NOS
C0009492|T047|PT|958.90|ICD9CM|Compartment syndrome, unspecified|Compartment syndrome, unspecified
C1719657|T037|AB|958.91|ICD9CM|Trauma comp synd up ext|Trauma comp synd up ext
C1719657|T037|PT|958.91|ICD9CM|Traumatic compartment syndrome of upper extremity|Traumatic compartment syndrome of upper extremity
C1719659|T037|AB|958.92|ICD9CM|Trauma comp synd low ext|Trauma comp synd low ext
C1719659|T037|PT|958.92|ICD9CM|Traumatic compartment syndrome of lower extremity|Traumatic compartment syndrome of lower extremity
C1719660|T037|AB|958.93|ICD9CM|Trauma compart synd abd|Trauma compart synd abd
C1719660|T037|PT|958.93|ICD9CM|Traumatic compartment syndrome of abdomen|Traumatic compartment syndrome of abdomen
C1719661|T037|AB|958.99|ICD9CM|Trauma compart synd NEC|Trauma compart synd NEC
C1719661|T037|PT|958.99|ICD9CM|Traumatic compartment syndrome of other sites|Traumatic compartment syndrome of other sites
C0302401|T037|HT|959|ICD9CM|Injury, other and unspecified|Injury, other and unspecified
C0490041|T037|HT|959.0|ICD9CM|Other and unspecified injury to head, face, and neck|Other and unspecified injury to head, face, and neck
C0018674|T037|AB|959.01|ICD9CM|Head injury NOS|Head injury NOS
C0018674|T037|PT|959.01|ICD9CM|Head injury, unspecified|Head injury, unspecified
C0272422|T037|AB|959.09|ICD9CM|Face & neck injury|Face & neck injury
C0272422|T037|PT|959.09|ICD9CM|Injury of face and neck|Injury of face and neck
C0029508|T037|HT|959.1|ICD9CM|Other and unspecified injury to trunk|Other and unspecified injury to trunk
C0436055|T037|AB|959.11|ICD9CM|Injury of chest wall NEC|Injury of chest wall NEC
C0436055|T037|PT|959.11|ICD9CM|Other injury of chest wall|Other injury of chest wall
C1260446|T037|AB|959.12|ICD9CM|Injury of abdomen NEC|Injury of abdomen NEC
C1260446|T037|PT|959.12|ICD9CM|Other injury of abdomen|Other injury of abdomen
C1260447|T037|PT|959.13|ICD9CM|Fracture of corpus cavernosum penis|Fracture of corpus cavernosum penis
C1260447|T037|AB|959.13|ICD9CM|Fx corpus cavrnosm penis|Fx corpus cavrnosm penis
C0436064|T037|AB|959.14|ICD9CM|Inj external genital NEC|Inj external genital NEC
C0436064|T037|PT|959.14|ICD9CM|Other injury of external genitals|Other injury of external genitals
C1260449|T037|PT|959.19|ICD9CM|Other injury of other sites of trunk|Other injury of other sites of trunk
C1260449|T037|AB|959.19|ICD9CM|Trunk injury-sites NEC|Trunk injury-sites NEC
C0161483|T037|AB|959.2|ICD9CM|Shldr/upper arm inj NOS|Shldr/upper arm inj NOS
C0161483|T037|PT|959.2|ICD9CM|Shoulder and upper arm injury|Shoulder and upper arm injury
C0272443|T037|AB|959.3|ICD9CM|Elb/forearm/wrst inj NOS|Elb/forearm/wrst inj NOS
C0272443|T037|PT|959.3|ICD9CM|Elbow, forearm, and wrist injury|Elbow, forearm, and wrist injury
C0029505|T037|AB|959.4|ICD9CM|Hand injury NOS|Hand injury NOS
C0029505|T037|PT|959.4|ICD9CM|Hand, except finger injury|Hand, except finger injury
C0016124|T037|PT|959.5|ICD9CM|Finger injury|Finger injury
C0016124|T037|AB|959.5|ICD9CM|Finger injury NOS|Finger injury NOS
C0161484|T037|AB|959.6|ICD9CM|Hip & thigh injury NOS|Hip & thigh injury NOS
C0161484|T037|PT|959.6|ICD9CM|Hip and thigh injury|Hip and thigh injury
C0029506|T037|PT|959.7|ICD9CM|Knee, leg, ankle, and foot injury|Knee, leg, ankle, and foot injury
C0029506|T037|AB|959.7|ICD9CM|Lower leg injury NOS|Lower leg injury NOS
C0029507|T037|AB|959.8|ICD9CM|Injury mlt site/site NEC|Injury mlt site/site NEC
C0029507|T037|PT|959.8|ICD9CM|Other specified sites, including multiple injury|Other specified sites, including multiple injury
C0029509|T037|AB|959.9|ICD9CM|Injury-site NOS|Injury-site NOS
C0029509|T037|PT|959.9|ICD9CM|Unspecified site injury|Unspecified site injury
C0161485|T037|HT|960|ICD9CM|Poisoning by antibiotics|Poisoning by antibiotics
C0178332|T037|HT|960-979.99|ICD9CM|POISONING BY DRUGS, MEDICINAL AND BIOLOGICAL SUBSTANCES|POISONING BY DRUGS, MEDICINAL AND BIOLOGICAL SUBSTANCES
C0161486|T037|PT|960.0|ICD9CM|Poisoning by penicillins|Poisoning by penicillins
C0161486|T037|AB|960.0|ICD9CM|Poisoning-penicillins|Poisoning-penicillins
C0161487|T037|AB|960.1|ICD9CM|Pois-antifungal antibiot|Pois-antifungal antibiot
C0161487|T037|PT|960.1|ICD9CM|Poisoning by antifungal antibiotics|Poisoning by antifungal antibiotics
C0161488|T037|AB|960.2|ICD9CM|Poison-chloramphenicol|Poison-chloramphenicol
C0161488|T037|PT|960.2|ICD9CM|Poisoning by chloramphenicol group|Poisoning by chloramphenicol group
C0161489|T037|AB|960.3|ICD9CM|Pois-erythromyc/macrolid|Pois-erythromyc/macrolid
C0161489|T037|PT|960.3|ICD9CM|Poisoning by erythromycin and other macrolides|Poisoning by erythromycin and other macrolides
C0274507|T037|PT|960.4|ICD9CM|Poisoning by tetracycline group|Poisoning by tetracycline group
C0274507|T037|AB|960.4|ICD9CM|Poisoning-tetracycline|Poisoning-tetracycline
C0274511|T037|AB|960.5|ICD9CM|Pois-cephalosporin group|Pois-cephalosporin group
C0274511|T037|PT|960.5|ICD9CM|Poisoning of cephalosporin group|Poisoning of cephalosporin group
C0274484|T037|AB|960.6|ICD9CM|Pois-antimycobac antibio|Pois-antimycobac antibio
C0274484|T037|PT|960.6|ICD9CM|Poisoning of antimycobacterial antibiotics|Poisoning of antimycobacterial antibiotics
C0161493|T037|AB|960.7|ICD9CM|Pois-antineop antibiotic|Pois-antineop antibiotic
C0161493|T037|PT|960.7|ICD9CM|Poisoning by antineoplastic antibiotics|Poisoning by antineoplastic antibiotics
C0161494|T037|PT|960.8|ICD9CM|Poisoning by other specified antibiotics|Poisoning by other specified antibiotics
C0161494|T037|AB|960.8|ICD9CM|Poisoning-antibiotic NEC|Poisoning-antibiotic NEC
C0161485|T037|PT|960.9|ICD9CM|Poisoning by unspecified antibiotic|Poisoning by unspecified antibiotic
C0161485|T037|AB|960.9|ICD9CM|Poisoning-antibiotic NOS|Poisoning-antibiotic NOS
C0161496|T037|HT|961|ICD9CM|Poisoning by other anti-infectives|Poisoning by other anti-infectives
C0161497|T037|PT|961.0|ICD9CM|Poisoning by sulfonamides|Poisoning by sulfonamides
C0161497|T037|AB|961.0|ICD9CM|Poisoning-sulfonamides|Poisoning-sulfonamides
C0161498|T037|AB|961.1|ICD9CM|Pois-arsenic anti-infec|Pois-arsenic anti-infec
C0161498|T037|PT|961.1|ICD9CM|Poisoning by arsenical anti-infectives|Poisoning by arsenical anti-infectives
C0161499|T037|AB|961.2|ICD9CM|Pois-heav met anti-infec|Pois-heav met anti-infec
C0161499|T037|PT|961.2|ICD9CM|Poisoning by heavy metal anti-infectives|Poisoning by heavy metal anti-infectives
C0347966|T037|AB|961.3|ICD9CM|Pois-quinoline/hydroxyqu|Pois-quinoline/hydroxyqu
C0347966|T037|PT|961.3|ICD9CM|Poisoning by quinoline and hydroxyquinoline derivatives|Poisoning by quinoline and hydroxyquinoline derivatives
C0161501|T037|PT|961.4|ICD9CM|Poisoning by antimalarials and drugs acting on other blood protozoa|Poisoning by antimalarials and drugs acting on other blood protozoa
C0161501|T037|AB|961.4|ICD9CM|Poisoning-antimalarials|Poisoning-antimalarials
C0161502|T037|AB|961.5|ICD9CM|Pois-antiprotoz drug NEC|Pois-antiprotoz drug NEC
C0161502|T037|PT|961.5|ICD9CM|Poisoning by other antiprotozoal drugs|Poisoning by other antiprotozoal drugs
C0496964|T037|PT|961.6|ICD9CM|Poisoning by anthelmintics|Poisoning by anthelmintics
C0496964|T037|AB|961.6|ICD9CM|Poisoning-anthelmintics|Poisoning-anthelmintics
C0161504|T037|PT|961.7|ICD9CM|Poisoning by antiviral drugs|Poisoning by antiviral drugs
C0161504|T037|AB|961.7|ICD9CM|Poisoning-antiviral drug|Poisoning-antiviral drug
C0161505|T037|AB|961.8|ICD9CM|Pois-antimycobac drg NEC|Pois-antimycobac drg NEC
C0161505|T037|PT|961.8|ICD9CM|Poisoning by other antimycobacterial drugs|Poisoning by other antimycobacterial drugs
C0161506|T037|AB|961.9|ICD9CM|Pois-anti-infect NEC/NOS|Pois-anti-infect NEC/NOS
C0161506|T037|PT|961.9|ICD9CM|Poisoning by other and unspecified anti-infectives|Poisoning by other and unspecified anti-infectives
C0274526|T037|HT|962|ICD9CM|Poisoning by hormones and synthetic substitutes|Poisoning by hormones and synthetic substitutes
C0161508|T037|AB|962.0|ICD9CM|Pois-corticosteroids|Pois-corticosteroids
C0161508|T037|PT|962.0|ICD9CM|Poisoning by adrenal cortical steroids|Poisoning by adrenal cortical steroids
C0161509|T037|PT|962.1|ICD9CM|Poisoning by androgens and anabolic congeners|Poisoning by androgens and anabolic congeners
C0161509|T037|AB|962.1|ICD9CM|Poisoning-androgens|Poisoning-androgens
C0274535|T037|PT|962.2|ICD9CM|Poisoning by ovarian hormones and synthetic substitutes|Poisoning by ovarian hormones and synthetic substitutes
C0274535|T037|AB|962.2|ICD9CM|Poisoning-ovarian hormon|Poisoning-ovarian hormon
C0496967|T037|AB|962.3|ICD9CM|Poison-insulin/antidiab|Poison-insulin/antidiab
C0496967|T037|PT|962.3|ICD9CM|Poisoning by insulins and antidiabetic agents|Poisoning by insulins and antidiabetic agents
C0161512|T037|AB|962.4|ICD9CM|Pois-ant pituitary horm|Pois-ant pituitary horm
C0161512|T037|PT|962.4|ICD9CM|Poisoning by anterior pituitary hormones|Poisoning by anterior pituitary hormones
C0161513|T037|AB|962.5|ICD9CM|Pois-post pituitary horm|Pois-post pituitary horm
C0161513|T037|PT|962.5|ICD9CM|Poisoning by posterior pituitary hormones|Poisoning by posterior pituitary hormones
C0161514|T037|PT|962.6|ICD9CM|Poisoning by parathyroid and parathyroid derivatives|Poisoning by parathyroid and parathyroid derivatives
C0161514|T037|AB|962.6|ICD9CM|Poisoning-parathyroids|Poisoning-parathyroids
C0161515|T037|PT|962.7|ICD9CM|Poisoning by thyroid and thyroid derivatives|Poisoning by thyroid and thyroid derivatives
C0161515|T037|AB|962.7|ICD9CM|Poisoning-thyroid/deriv|Poisoning-thyroid/deriv
C0161516|T037|AB|962.8|ICD9CM|Poison-antithyroid agent|Poison-antithyroid agent
C0161516|T037|PT|962.8|ICD9CM|Poisoning by antithyroid agents|Poisoning by antithyroid agents
C0161517|T037|PT|962.9|ICD9CM|Poisoning by other and unspecified hormones and synthetic substitutes|Poisoning by other and unspecified hormones and synthetic substitutes
C0161517|T037|AB|962.9|ICD9CM|Poisoning hormon NEC/NOS|Poisoning hormon NEC/NOS
C0161518|T037|HT|963|ICD9CM|Poisoning by primarily systemic agents|Poisoning by primarily systemic agents
C0161519|T037|AB|963.0|ICD9CM|Pois-antiallrg/antiemet|Pois-antiallrg/antiemet
C0161519|T037|PT|963.0|ICD9CM|Poisoning by antiallergic and antiemetic drugs|Poisoning by antiallergic and antiemetic drugs
C0412836|T037|AB|963.1|ICD9CM|Pois-antineopl/immunosup|Pois-antineopl/immunosup
C0412836|T037|PT|963.1|ICD9CM|Poisoning by antineoplastic and immunosuppressive drugs|Poisoning by antineoplastic and immunosuppressive drugs
C0161521|T037|PT|963.2|ICD9CM|Poisoning by acidifying agents|Poisoning by acidifying agents
C0161521|T037|AB|963.2|ICD9CM|Poisoning-acidifying agt|Poisoning-acidifying agt
C0161522|T037|PT|963.3|ICD9CM|Poisoning by alkalizing agents|Poisoning by alkalizing agents
C0161522|T037|AB|963.3|ICD9CM|Poisoning-alkalizing agt|Poisoning-alkalizing agt
C0869507|T037|PT|963.4|ICD9CM|Poisoning by enzymes, not elsewhere classified|Poisoning by enzymes, not elsewhere classified
C0869507|T037|AB|963.4|ICD9CM|Poisoning-enzymes NEC|Poisoning-enzymes NEC
C0869511|T037|PT|963.5|ICD9CM|Poisoning by vitamins, not elsewhere classified|Poisoning by vitamins, not elsewhere classified
C0869511|T037|AB|963.5|ICD9CM|Poisoning-vitamins NEC|Poisoning-vitamins NEC
C0161525|T037|PT|963.8|ICD9CM|Poisoning by other specified systemic agents|Poisoning by other specified systemic agents
C0161525|T037|AB|963.8|ICD9CM|Poisoning-system agt NEC|Poisoning-system agt NEC
C0161518|T037|PT|963.9|ICD9CM|Poisoning by unspecified systemic agent|Poisoning by unspecified systemic agent
C0161518|T037|AB|963.9|ICD9CM|Poisoning-system agt NOS|Poisoning-system agt NOS
C0161527|T037|HT|964|ICD9CM|Poisoning by agents primarily affecting blood constituents|Poisoning by agents primarily affecting blood constituents
C0412842|T037|PT|964.0|ICD9CM|Poisoning by iron and its compounds|Poisoning by iron and its compounds
C0412842|T037|AB|964.0|ICD9CM|Poisoning-iron/compounds|Poisoning-iron/compounds
C0161529|T037|AB|964.1|ICD9CM|Poison-liver/antianemics|Poison-liver/antianemics
C0161529|T037|PT|964.1|ICD9CM|Poisoning by liver preparations and other antianemic agents|Poisoning by liver preparations and other antianemic agents
C0161530|T037|PT|964.2|ICD9CM|Poisoning by anticoagulants|Poisoning by anticoagulants
C0161530|T037|AB|964.2|ICD9CM|Poisoning-anticoagulants|Poisoning-anticoagulants
C0274594|T037|PT|964.3|ICD9CM|Poisoning by vitamin K (phytonadione)|Poisoning by vitamin K (phytonadione)
C0274594|T037|AB|964.3|ICD9CM|Poisoning-vitamin k|Poisoning-vitamin k
C0412845|T037|AB|964.4|ICD9CM|Poison-fibrinolysis agnt|Poison-fibrinolysis agnt
C0412845|T037|PT|964.4|ICD9CM|Poisoning by fibrinolysis-affecting drugs|Poisoning by fibrinolysis-affecting drugs
C0161533|T037|PT|964.5|ICD9CM|Poisoning by anticoagulant antagonists and other coagulants|Poisoning by anticoagulant antagonists and other coagulants
C0161533|T037|AB|964.5|ICD9CM|Poisoning-coagulants|Poisoning-coagulants
C0161534|T037|PT|964.6|ICD9CM|Poisoning by gamma globulin|Poisoning by gamma globulin
C0161534|T037|AB|964.6|ICD9CM|Poisoning-gamma globulin|Poisoning-gamma globulin
C0274602|T037|PT|964.7|ICD9CM|Poisoning by natural blood and blood products|Poisoning by natural blood and blood products
C0274602|T037|AB|964.7|ICD9CM|Poisoning-blood product|Poisoning-blood product
C0161536|T037|PT|964.8|ICD9CM|Poisoning by other specified agents affecting blood constituents|Poisoning by other specified agents affecting blood constituents
C0161536|T037|AB|964.8|ICD9CM|Poisoning-blood agt NEC|Poisoning-blood agt NEC
C0161537|T037|PT|964.9|ICD9CM|Poisoning by unspecified agent affecting blood constituents|Poisoning by unspecified agent affecting blood constituents
C0161537|T037|AB|964.9|ICD9CM|Poisoning-blood agt NOS|Poisoning-blood agt NOS
C0161538|T037|HT|965|ICD9CM|Poisoning by analgesics, antipyretics, and antirheumatics|Poisoning by analgesics, antipyretics, and antirheumatics
C1443030|T037|HT|965.0|ICD9CM|Poisoning by opiates and related narcotics|Poisoning by opiates and related narcotics
C0161540|T037|PT|965.00|ICD9CM|Poisoning by opium (alkaloids), unspecified|Poisoning by opium (alkaloids), unspecified
C0161540|T037|AB|965.00|ICD9CM|Poisoning-opium NOS|Poisoning-opium NOS
C0161541|T037|PT|965.01|ICD9CM|Poisoning by heroin|Poisoning by heroin
C0161541|T037|AB|965.01|ICD9CM|Poisoning-heroin|Poisoning-heroin
C0161542|T037|PT|965.02|ICD9CM|Poisoning by methadone|Poisoning by methadone
C0161542|T037|AB|965.02|ICD9CM|Poisoning-methadone|Poisoning-methadone
C0161543|T037|PT|965.09|ICD9CM|Poisoning by other opiates and related narcotics|Poisoning by other opiates and related narcotics
C0161543|T037|AB|965.09|ICD9CM|Poisoning-opiates NEC|Poisoning-opiates NEC
C0161544|T037|PT|965.1|ICD9CM|Poisoning by salicylates|Poisoning by salicylates
C0161544|T037|AB|965.1|ICD9CM|Poisoning-salicylates|Poisoning-salicylates
C0868775|T037|AB|965.4|ICD9CM|Pois-arom analgesics NEC|Pois-arom analgesics NEC
C0868775|T037|PT|965.4|ICD9CM|Poisoning by aromatic analgesics, not elsewhere classified|Poisoning by aromatic analgesics, not elsewhere classified
C0161546|T037|PT|965.5|ICD9CM|Poisoning by pyrazole derivatives|Poisoning by pyrazole derivatives
C0161546|T037|AB|965.5|ICD9CM|Poisoning-pyrazole deriv|Poisoning-pyrazole deriv
C0344128|T037|HT|965.6|ICD9CM|Poisoning by antirheumatics [antiphlogistics]|Poisoning by antirheumatics [antiphlogistics]
C0695274|T037|AB|965.61|ICD9CM|Pois-propionic acid derv|Pois-propionic acid derv
C0695274|T037|PT|965.61|ICD9CM|Poisoning by propionic acid derivatives|Poisoning by propionic acid derivatives
C0695253|T037|AB|965.69|ICD9CM|Poison-antirheumatic NEC|Poison-antirheumatic NEC
C0695253|T037|PT|965.69|ICD9CM|Poisoning by other antirheumatics|Poisoning by other antirheumatics
C0161548|T037|AB|965.7|ICD9CM|Pois-no-narc analges NEC|Pois-no-narc analges NEC
C0161548|T037|PT|965.7|ICD9CM|Poisoning by other non-narcotic analgesics|Poisoning by other non-narcotic analgesics
C0161549|T037|AB|965.8|ICD9CM|Pois-analges/antipyr NEC|Pois-analges/antipyr NEC
C0161549|T037|PT|965.8|ICD9CM|Poisoning by other specified analgesics and antipyretics|Poisoning by other specified analgesics and antipyretics
C0274609|T037|AB|965.9|ICD9CM|Pois-analges/antipyr NOS|Pois-analges/antipyr NOS
C0274609|T037|PT|965.9|ICD9CM|Poisoning by unspecified analgesic and antipyretic|Poisoning by unspecified analgesic and antipyretic
C0412928|T037|HT|966|ICD9CM|Poisoning by anticonvulsants and anti-Parkinsonism drugs|Poisoning by anticonvulsants and anti-Parkinsonism drugs
C0161552|T037|AB|966.0|ICD9CM|Poison-oxazolidine deriv|Poison-oxazolidine deriv
C0161552|T037|PT|966.0|ICD9CM|Poisoning by oxazolidine derivatives|Poisoning by oxazolidine derivatives
C0161553|T037|AB|966.1|ICD9CM|Poison-hydantoin derivat|Poison-hydantoin derivat
C0161553|T037|PT|966.1|ICD9CM|Poisoning by hydantoin derivatives|Poisoning by hydantoin derivatives
C0161554|T037|PT|966.2|ICD9CM|Poisoning by succinimides|Poisoning by succinimides
C0161554|T037|AB|966.2|ICD9CM|Poisoning-succinimides|Poisoning-succinimides
C0161555|T037|AB|966.3|ICD9CM|Pois-anticonvul NEC/NOS|Pois-anticonvul NEC/NOS
C0161555|T037|PT|966.3|ICD9CM|Poisoning by other and unspecified anticonvulsants|Poisoning by other and unspecified anticonvulsants
C0161556|T037|AB|966.4|ICD9CM|Pois-anti-parkinson drug|Pois-anti-parkinson drug
C0161556|T037|PT|966.4|ICD9CM|Poisoning by anti-Parkinsonism drugs|Poisoning by anti-Parkinsonism drugs
C0274638|T037|HT|967|ICD9CM|Poisoning by sedatives and hypnotics|Poisoning by sedatives and hypnotics
C0161558|T037|PT|967.0|ICD9CM|Poisoning by barbiturates|Poisoning by barbiturates
C0161558|T037|AB|967.0|ICD9CM|Poisoning-barbiturates|Poisoning-barbiturates
C0344156|T037|PT|967.1|ICD9CM|Poisoning by chloral hydrate group|Poisoning by chloral hydrate group
C0344156|T037|AB|967.1|ICD9CM|Poisoning-chloral hydrat|Poisoning-chloral hydrat
C0161560|T037|PT|967.2|ICD9CM|Poisoning by paraldehyde|Poisoning by paraldehyde
C0161560|T037|AB|967.2|ICD9CM|Poisoning-paraldehyde|Poisoning-paraldehyde
C1533166|T037|PT|967.3|ICD9CM|Poisoning by bromine compounds|Poisoning by bromine compounds
C1533166|T037|AB|967.3|ICD9CM|Poisoning-bromine compnd|Poisoning-bromine compnd
C0161562|T037|PT|967.4|ICD9CM|Poisoning by methaqualone compounds|Poisoning by methaqualone compounds
C0161562|T037|AB|967.4|ICD9CM|Poisoning-methaqualone|Poisoning-methaqualone
C0161563|T037|PT|967.5|ICD9CM|Poisoning by glutethimide group|Poisoning by glutethimide group
C0161563|T037|AB|967.5|ICD9CM|Poisoning-glutethimide|Poisoning-glutethimide
C0868780|T037|AB|967.6|ICD9CM|Poison-mix sedative NEC|Poison-mix sedative NEC
C0868780|T037|PT|967.6|ICD9CM|Poisoning by mixed sedatives, not elsewhere classified|Poisoning by mixed sedatives, not elsewhere classified
C0161565|T037|AB|967.8|ICD9CM|Pois-sedative/hypnot NEC|Pois-sedative/hypnot NEC
C0161565|T037|PT|967.8|ICD9CM|Poisoning by other sedatives and hypnotics|Poisoning by other sedatives and hypnotics
C0274638|T037|AB|967.9|ICD9CM|Pois-sedative/hypnot NOS|Pois-sedative/hypnot NOS
C0274638|T037|PT|967.9|ICD9CM|Poisoning by unspecified sedative or hypnotic|Poisoning by unspecified sedative or hypnotic
C0161567|T037|HT|968|ICD9CM|Poisoning by other central nervous system depressants and anesthetics|Poisoning by other central nervous system depressants and anesthetics
C0161568|T037|AB|968.0|ICD9CM|Pois-cns muscle depress|Pois-cns muscle depress
C0161568|T037|PT|968.0|ICD9CM|Poisoning by central nervous system muscle-tone depressants|Poisoning by central nervous system muscle-tone depressants
C0161569|T037|PT|968.1|ICD9CM|Poisoning by halothane|Poisoning by halothane
C0161569|T037|AB|968.1|ICD9CM|Poisoning-halothane|Poisoning-halothane
C0473975|T037|AB|968.2|ICD9CM|Poison-gas anesthet NEC|Poison-gas anesthet NEC
C0473975|T037|PT|968.2|ICD9CM|Poisoning by other gaseous anesthetics|Poisoning by other gaseous anesthetics
C0161571|T037|AB|968.3|ICD9CM|Poison-intraven anesthet|Poison-intraven anesthet
C0161571|T037|PT|968.3|ICD9CM|Poisoning by intravenous anesthetics|Poisoning by intravenous anesthetics
C0161572|T037|AB|968.4|ICD9CM|Pois-gen anesth NEC/NOS|Pois-gen anesth NEC/NOS
C0161572|T037|PT|968.4|ICD9CM|Poisoning by other and unspecified general anesthetics|Poisoning by other and unspecified general anesthetics
C0161573|T037|PT|968.5|ICD9CM|Surface (topical) and infiltration anesthetics|Surface (topical) and infiltration anesthetics
C0161573|T037|AB|968.5|ICD9CM|Surfce-topic/infilt anes|Surfce-topic/infilt anes
C0161574|T037|AB|968.6|ICD9CM|Pois-nerve/plex-blk anes|Pois-nerve/plex-blk anes
C0161574|T037|PT|968.6|ICD9CM|Poisoning by peripheral nerve- and plexus-blocking anesthetics|Poisoning by peripheral nerve- and plexus-blocking anesthetics
C0161575|T037|AB|968.7|ICD9CM|Poison-spinal anesthetic|Poison-spinal anesthetic
C0161575|T037|PT|968.7|ICD9CM|Poisoning by spinal anesthetics|Poisoning by spinal anesthetics
C0161576|T037|AB|968.9|ICD9CM|Pois-local anest NEC/NOS|Pois-local anest NEC/NOS
C0161576|T037|PT|968.9|ICD9CM|Poisoning by other and unspecified local anesthetics|Poisoning by other and unspecified local anesthetics
C0161577|T037|HT|969|ICD9CM|Poisoning by psychotropic agents|Poisoning by psychotropic agents
C0161578|T037|HT|969.0|ICD9CM|Poisoning by antidepressants|Poisoning by antidepressants
C2712374|T037|AB|969.00|ICD9CM|Poison-antidepresnt NOS|Poison-antidepresnt NOS
C2712374|T037|PT|969.00|ICD9CM|Poisoning by antidepressant, unspecified|Poisoning by antidepressant, unspecified
C0274669|T037|AB|969.01|ICD9CM|Pois monoamine oxidase|Pois monoamine oxidase
C0274669|T037|PT|969.01|ICD9CM|Poisoning by monoamine oxidase inhibitors|Poisoning by monoamine oxidase inhibitors
C2712375|T037|AB|969.02|ICD9CM|Pois serotn/norepinephrn|Pois serotn/norepinephrn
C2712375|T037|PT|969.02|ICD9CM|Poisoning by selective serotonin and norepinephrine reuptake inhibitors|Poisoning by selective serotonin and norepinephrine reuptake inhibitors
C2712376|T037|AB|969.03|ICD9CM|Pois serotinin reuptake|Pois serotinin reuptake
C2712376|T037|PT|969.03|ICD9CM|Poisoning by selective serotonin reuptake inhibitors|Poisoning by selective serotonin reuptake inhibitors
C2712377|T037|AB|969.04|ICD9CM|Pois tetracyclc andepres|Pois tetracyclc andepres
C2712377|T037|PT|969.04|ICD9CM|Poisoning by tetracyclic antidepressants|Poisoning by tetracyclic antidepressants
C0496978|T037|AB|969.05|ICD9CM|Pois tricyclc antidepres|Pois tricyclc antidepres
C0496978|T037|PT|969.05|ICD9CM|Poisoning by tricyclic antidepressants|Poisoning by tricyclic antidepressants
C2712378|T037|AB|969.09|ICD9CM|Pois antidepressants NEC|Pois antidepressants NEC
C2712378|T037|PT|969.09|ICD9CM|Poisoning by other antidepressants|Poisoning by other antidepressants
C0274967|T037|AB|969.1|ICD9CM|Pois-phenothiazine tranq|Pois-phenothiazine tranq
C0274967|T037|PT|969.1|ICD9CM|Poisoning by phenothiazine-based tranquilizers|Poisoning by phenothiazine-based tranquilizers
C0344133|T037|AB|969.2|ICD9CM|Pois-butyrophenone tranq|Pois-butyrophenone tranq
C0344133|T037|PT|969.2|ICD9CM|Poisoning by butyrophenone-based tranquilizers|Poisoning by butyrophenone-based tranquilizers
C0161581|T037|AB|969.3|ICD9CM|Poison-antipsychotic NEC|Poison-antipsychotic NEC
C0161581|T037|PT|969.3|ICD9CM|Poisoning by other antipsychotics, neuroleptics, and major tranquilizers|Poisoning by other antipsychotics, neuroleptics, and major tranquilizers
C0412862|T037|AB|969.4|ICD9CM|Pois-benzodiazepine tran|Pois-benzodiazepine tran
C0412862|T037|PT|969.4|ICD9CM|Poisoning by benzodiazepine-based tranquilizers|Poisoning by benzodiazepine-based tranquilizers
C0161583|T037|AB|969.5|ICD9CM|Poison-tranquilizer NEC|Poison-tranquilizer NEC
C0161583|T037|PT|969.5|ICD9CM|Poisoning by other tranquilizers|Poisoning by other tranquilizers
C0161584|T037|PT|969.6|ICD9CM|Poisoning by psychodysleptics (hallucinogens)|Poisoning by psychodysleptics (hallucinogens)
C0161584|T037|AB|969.6|ICD9CM|Poisoning-hallucinogens|Poisoning-hallucinogens
C0161585|T037|HT|969.7|ICD9CM|Poisoning by psychostimulants|Poisoning by psychostimulants
C2712379|T037|AB|969.70|ICD9CM|Pois psychostimulant NOS|Pois psychostimulant NOS
C2712379|T037|PT|969.70|ICD9CM|Poisoning by psychostimulant, unspecified|Poisoning by psychostimulant, unspecified
C0274693|T037|PT|969.71|ICD9CM|Poisoning by caffeine|Poisoning by caffeine
C0274693|T037|AB|969.71|ICD9CM|Poisoning by caffeine|Poisoning by caffeine
C0274692|T037|AB|969.72|ICD9CM|Poisoning by amphetamine|Poisoning by amphetamine
C0274692|T037|PT|969.72|ICD9CM|Poisoning by amphetamines|Poisoning by amphetamines
C2712380|T037|AB|969.73|ICD9CM|Poison by methylphendate|Poison by methylphendate
C2712380|T037|PT|969.73|ICD9CM|Poisoning by methylphenidate|Poisoning by methylphenidate
C2712381|T037|AB|969.79|ICD9CM|Poison by psychostim NEC|Poison by psychostim NEC
C2712381|T037|PT|969.79|ICD9CM|Poisoning by other psychostimulants|Poisoning by other psychostimulants
C0161586|T037|AB|969.8|ICD9CM|Poison-psychotropic NEC|Poison-psychotropic NEC
C0161586|T037|PT|969.8|ICD9CM|Poisoning by other specified psychotropic agents|Poisoning by other specified psychotropic agents
C0161577|T037|AB|969.9|ICD9CM|Poison-psychotropic NOS|Poison-psychotropic NOS
C0161577|T037|PT|969.9|ICD9CM|Poisoning by unspecified psychotropic agent|Poisoning by unspecified psychotropic agent
C0161588|T037|HT|970|ICD9CM|Poisoning by central nervous system stimulants|Poisoning by central nervous system stimulants
C0161589|T037|PT|970.0|ICD9CM|Poisoning by analeptics|Poisoning by analeptics
C0161589|T037|AB|970.0|ICD9CM|Poisoning-analeptics|Poisoning-analeptics
C0161590|T037|AB|970.1|ICD9CM|Poison-opiate antagonist|Poison-opiate antagonist
C0161590|T037|PT|970.1|ICD9CM|Poisoning by opiate antagonists|Poisoning by opiate antagonists
C0161591|T037|HT|970.8|ICD9CM|Poisoning by other specified central nervous system stimulants|Poisoning by other specified central nervous system stimulants
C0274659|T037|PT|970.81|ICD9CM|Poisoning by cocaine|Poisoning by cocaine
C0274659|T037|AB|970.81|ICD9CM|Poisoning by cocaine|Poisoning by cocaine
C0412869|T037|AB|970.89|ICD9CM|Poison-CNS stimulant NEC|Poison-CNS stimulant NEC
C0412869|T037|PT|970.89|ICD9CM|Poisoning by other central nervous system stimulants|Poisoning by other central nervous system stimulants
C0161588|T037|AB|970.9|ICD9CM|Pois-cns stimulant NOS|Pois-cns stimulant NOS
C0161588|T037|PT|970.9|ICD9CM|Poisoning by unspecified central nervous system stimulant|Poisoning by unspecified central nervous system stimulant
C0161593|T037|HT|971|ICD9CM|Poisoning by drugs primarily affecting the autonomic nervous system|Poisoning by drugs primarily affecting the autonomic nervous system
C0274702|T037|AB|971.0|ICD9CM|Pois-parasympathomimetic|Pois-parasympathomimetic
C0274702|T037|PT|971.0|ICD9CM|Poisoning by parasympathomimetics (cholinergics)|Poisoning by parasympathomimetics (cholinergics)
C0412870|T037|AB|971.1|ICD9CM|Pois-parasympatholytics|Pois-parasympatholytics
C0412870|T037|PT|971.1|ICD9CM|Poisoning by parasympatholytics (anticholinergics and antimuscarinics) and spasmolytics|Poisoning by parasympatholytics (anticholinergics and antimuscarinics) and spasmolytics
C0274714|T037|AB|971.2|ICD9CM|Poison-sympathomimetics|Poison-sympathomimetics
C0274714|T037|PT|971.2|ICD9CM|Poisoning by sympathomimetics [adrenergics]|Poisoning by sympathomimetics [adrenergics]
C0274717|T037|PT|971.3|ICD9CM|Poisoning by sympatholytics [antiadrenergics]|Poisoning by sympatholytics [antiadrenergics]
C0274717|T037|AB|971.3|ICD9CM|Poisoning-sympatholytics|Poisoning-sympatholytics
C0161598|T037|AB|971.9|ICD9CM|Pois-autonomic agent NOS|Pois-autonomic agent NOS
C0161598|T037|PT|971.9|ICD9CM|Poisoning by unspecified drug primarily affecting autonomic nervous system|Poisoning by unspecified drug primarily affecting autonomic nervous system
C0161599|T037|HT|972|ICD9CM|Poisoning by agents primarily affecting the cardiovascular system|Poisoning by agents primarily affecting the cardiovascular system
C0412873|T037|AB|972.0|ICD9CM|Pois-card rhythm regulat|Pois-card rhythm regulat
C0412873|T037|PT|972.0|ICD9CM|Poisoning by cardiac rhythm regulators|Poisoning by cardiac rhythm regulators
C0161601|T037|PT|972.1|ICD9CM|Poisoning by cardiotonic glycosides and drugs of similar action|Poisoning by cardiotonic glycosides and drugs of similar action
C0161601|T037|AB|972.1|ICD9CM|Poisoning-cardiotonics|Poisoning-cardiotonics
C0161602|T037|PT|972.2|ICD9CM|Poisoning by antilipemic and antiarteriosclerotic drugs|Poisoning by antilipemic and antiarteriosclerotic drugs
C0161602|T037|AB|972.2|ICD9CM|Poisoning-antilipemics|Poisoning-antilipemics
C0161603|T037|AB|972.3|ICD9CM|Pois-ganglion block agt|Pois-ganglion block agt
C0161603|T037|PT|972.3|ICD9CM|Poisoning by ganglion-blocking agents|Poisoning by ganglion-blocking agents
C0161604|T037|AB|972.4|ICD9CM|Pois-coronary vasodilat|Pois-coronary vasodilat
C0161604|T037|PT|972.4|ICD9CM|Poisoning by coronary vasodilators|Poisoning by coronary vasodilators
C0161605|T037|AB|972.5|ICD9CM|Poison-vasodilator NEC|Poison-vasodilator NEC
C0161605|T037|PT|972.5|ICD9CM|Poisoning by other vasodilators|Poisoning by other vasodilators
C0161606|T037|AB|972.6|ICD9CM|Pois-antihyperten agent|Pois-antihyperten agent
C0161606|T037|PT|972.6|ICD9CM|Poisoning by other antihypertensive agents|Poisoning by other antihypertensive agents
C0161607|T037|AB|972.7|ICD9CM|Poison-antivaricose drug|Poison-antivaricose drug
C0161607|T037|PT|972.7|ICD9CM|Poisoning by antivaricose drugs, including sclerosing agents|Poisoning by antivaricose drugs, including sclerosing agents
C0161608|T037|AB|972.8|ICD9CM|Poison-capillary act agt|Poison-capillary act agt
C0161608|T037|PT|972.8|ICD9CM|Poisoning by capillary-active drugs|Poisoning by capillary-active drugs
C0161609|T037|AB|972.9|ICD9CM|Pois-cardiovasc agt NEC|Pois-cardiovasc agt NEC
C0161609|T037|PT|972.9|ICD9CM|Poisoning by other and unspecified agents primarily affecting the cardiovascular system|Poisoning by other and unspecified agents primarily affecting the cardiovascular system
C0161610|T037|HT|973|ICD9CM|Poisoning by agents primarily affecting the gastrointestinal system|Poisoning by agents primarily affecting the gastrointestinal system
C0161611|T037|AB|973.0|ICD9CM|Pois-antacid/antigastric|Pois-antacid/antigastric
C0161611|T037|PT|973.0|ICD9CM|Poisoning by antacids and antigastric secretion drugs|Poisoning by antacids and antigastric secretion drugs
C0161612|T037|AB|973.1|ICD9CM|Pois-irritant cathartics|Pois-irritant cathartics
C0161612|T037|PT|973.1|ICD9CM|Poisoning by irritant cathartics|Poisoning by irritant cathartics
C0161613|T037|AB|973.2|ICD9CM|Pois-emollient cathartic|Pois-emollient cathartic
C0161613|T037|PT|973.2|ICD9CM|Poisoning by emollient cathartics|Poisoning by emollient cathartics
C3161460|T037|PT|973.3|ICD9CM|Poisoning by other cathartics, including intestinal atonia|Poisoning by other cathartics, including intestinal atonia
C3161460|T037|AB|973.3|ICD9CM|Poisoning-cathartic NEC|Poisoning-cathartic NEC
C0161615|T037|PT|973.4|ICD9CM|Poisoning by digestants|Poisoning by digestants
C0161615|T037|AB|973.4|ICD9CM|Poisoning-digestants|Poisoning-digestants
C0161616|T037|PT|973.5|ICD9CM|Poisoning by antidiarrheal drugs|Poisoning by antidiarrheal drugs
C0161616|T037|AB|973.5|ICD9CM|Poisoning-antidiarrh agt|Poisoning-antidiarrh agt
C0161617|T037|PT|973.6|ICD9CM|Poisoning by emetics|Poisoning by emetics
C0161617|T037|AB|973.6|ICD9CM|Poisoning-emetics|Poisoning-emetics
C0161618|T037|PT|973.8|ICD9CM|Poisoning by other specified agents primarily affecting the gastrointestinal system|Poisoning by other specified agents primarily affecting the gastrointestinal system
C0161618|T037|AB|973.8|ICD9CM|Poisoning-gi agents NEC|Poisoning-gi agents NEC
C0161619|T037|PT|973.9|ICD9CM|Poisoning by unspecified agent primarily affecting the gastrointestinal system|Poisoning by unspecified agent primarily affecting the gastrointestinal system
C0161619|T037|AB|973.9|ICD9CM|Poisoning-gi agent NOS|Poisoning-gi agent NOS
C0859760|T037|HT|974|ICD9CM|Poisoning by water, mineral, and uric acid metabolism drugs|Poisoning by water, mineral, and uric acid metabolism drugs
C0161621|T037|AB|974.0|ICD9CM|Pois-mercurial diuretics|Pois-mercurial diuretics
C0161621|T037|PT|974.0|ICD9CM|Poisoning by mercurial diuretics|Poisoning by mercurial diuretics
C0161622|T037|AB|974.1|ICD9CM|Pois-purine diuretics|Pois-purine diuretics
C0161622|T037|PT|974.1|ICD9CM|Poisoning by purine derivative diuretics|Poisoning by purine derivative diuretics
C0161623|T037|AB|974.2|ICD9CM|Pois-h2co3 anhydra inhib|Pois-h2co3 anhydra inhib
C0161623|T037|PT|974.2|ICD9CM|Poisoning by carbonic acid anhydrase inhibitors|Poisoning by carbonic acid anhydrase inhibitors
C0161624|T037|PT|974.3|ICD9CM|Poisoning by saluretics|Poisoning by saluretics
C0161624|T037|AB|974.3|ICD9CM|Poisoning-saluretics|Poisoning-saluretics
C0161625|T037|PT|974.4|ICD9CM|Poisoning by other diuretics|Poisoning by other diuretics
C0161625|T037|AB|974.4|ICD9CM|Poisoning-diuretics NEC|Poisoning-diuretics NEC
C0161626|T037|AB|974.5|ICD9CM|Pois-electro/cal/wat agt|Pois-electro/cal/wat agt
C0161626|T037|PT|974.5|ICD9CM|Poisoning by electrolytic, caloric, and water-balance agents|Poisoning by electrolytic, caloric, and water-balance agents
C0302406|T037|AB|974.6|ICD9CM|Poison-mineral salts NEC|Poison-mineral salts NEC
C0302406|T037|PT|974.6|ICD9CM|Poisoning by other mineral salts, not elsewhere classified|Poisoning by other mineral salts, not elsewhere classified
C0161628|T037|AB|974.7|ICD9CM|Pois-uric acid metabol|Pois-uric acid metabol
C0161628|T037|PT|974.7|ICD9CM|Poisoning by uric acid metabolism drugs|Poisoning by uric acid metabolism drugs
C0161629|T037|HT|975|ICD9CM|Poisoning by agents primarily acting on the smooth and skeletal muscles and respiratory system|Poisoning by agents primarily acting on the smooth and skeletal muscles and respiratory system
C0161630|T037|PT|975.0|ICD9CM|Poisoning by oxytocic agents|Poisoning by oxytocic agents
C0161630|T037|AB|975.0|ICD9CM|Poisoning-oxytocic agent|Poisoning-oxytocic agent
C0161631|T037|AB|975.1|ICD9CM|Pois-smooth muscle relax|Pois-smooth muscle relax
C0161631|T037|PT|975.1|ICD9CM|Poisoning by smooth muscle relaxants|Poisoning by smooth muscle relaxants
C0161632|T037|AB|975.2|ICD9CM|Pois-skelet muscle relax|Pois-skelet muscle relax
C0161632|T037|PT|975.2|ICD9CM|Poisoning by skeletal muscle relaxants|Poisoning by skeletal muscle relaxants
C0161633|T037|AB|975.3|ICD9CM|Poison-muscle agent NEC|Poison-muscle agent NEC
C0161633|T037|PT|975.3|ICD9CM|Poisoning by other and unspecified drugs acting on muscles|Poisoning by other and unspecified drugs acting on muscles
C0161634|T037|PT|975.4|ICD9CM|Poisoning by antitussives|Poisoning by antitussives
C0161634|T037|AB|975.4|ICD9CM|Poisoning-antitussives|Poisoning-antitussives
C0161635|T037|PT|975.5|ICD9CM|Poisoning by expectorants|Poisoning by expectorants
C0161635|T037|AB|975.5|ICD9CM|Poisoning-expectorants|Poisoning-expectorants
C0161636|T037|AB|975.6|ICD9CM|Pois-anti-cold drugs|Pois-anti-cold drugs
C0161636|T037|PT|975.6|ICD9CM|Poisoning by anti-common cold drugs|Poisoning by anti-common cold drugs
C0161637|T037|PT|975.7|ICD9CM|Poisoning by antiasthmatics|Poisoning by antiasthmatics
C0161637|T037|AB|975.7|ICD9CM|Poisoning-antiasthmatics|Poisoning-antiasthmatics
C0478453|T037|AB|975.8|ICD9CM|Pois-respir drug NEC/NOS|Pois-respir drug NEC/NOS
C0478453|T037|PT|975.8|ICD9CM|Poisoning by other and unspecified respiratory drugs|Poisoning by other and unspecified respiratory drugs
C0161640|T037|AB|976.0|ICD9CM|Pois-local anti-infect|Pois-local anti-infect
C0161640|T037|PT|976.0|ICD9CM|Poisoning by local anti-infectives and anti-inflammatory drugs|Poisoning by local anti-infectives and anti-inflammatory drugs
C0161641|T037|PT|976.1|ICD9CM|Poisoning by antipruritics|Poisoning by antipruritics
C0161641|T037|AB|976.1|ICD9CM|Poisoning-antipruritics|Poisoning-antipruritics
C0161642|T037|AB|976.2|ICD9CM|Pois-loc astring/deterg|Pois-loc astring/deterg
C0161642|T037|PT|976.2|ICD9CM|Poisoning by local astringents and local detergents|Poisoning by local astringents and local detergents
C0161643|T037|AB|976.3|ICD9CM|Pois-emol/demul/protect|Pois-emol/demul/protect
C0161643|T037|PT|976.3|ICD9CM|Poisoning by emollients, demulcents, and protectants|Poisoning by emollients, demulcents, and protectants
C0161644|T037|AB|976.4|ICD9CM|Poison-hair/scalp prep|Poison-hair/scalp prep
C0161644|T037|PT|976.4|ICD9CM|Poisoning by keratolytics, keratoplastics, other hair treatment drugs and preparations|Poisoning by keratolytics, keratoplastics, other hair treatment drugs and preparations
C0161645|T037|AB|976.5|ICD9CM|Pois-eye anti-infec/drug|Pois-eye anti-infec/drug
C0161645|T037|PT|976.5|ICD9CM|Poisoning by eye anti-infectives and other eye drugs|Poisoning by eye anti-infectives and other eye drugs
C0161646|T037|AB|976.6|ICD9CM|Poison-ent preparation|Poison-ent preparation
C0161646|T037|PT|976.6|ICD9CM|Poisoning by anti-infectives and other drugs and preparations for ear, nose, and throat|Poisoning by anti-infectives and other drugs and preparations for ear, nose, and throat
C0161647|T037|AB|976.7|ICD9CM|Pois-topical dental drug|Pois-topical dental drug
C0161647|T037|PT|976.7|ICD9CM|Poisoning by dental drugs topically applied|Poisoning by dental drugs topically applied
C0161648|T037|AB|976.8|ICD9CM|Pois-skin/membr agnt NEC|Pois-skin/membr agnt NEC
C0161648|T037|PT|976.8|ICD9CM|Poisoning by other agents primarily affecting skin and mucous membrane|Poisoning by other agents primarily affecting skin and mucous membrane
C0161649|T037|AB|976.9|ICD9CM|Pois-skin/membr agnt NOS|Pois-skin/membr agnt NOS
C0161649|T037|PT|976.9|ICD9CM|Poisoning by unspecified agent primarily affecting skin and mucous membrane|Poisoning by unspecified agent primarily affecting skin and mucous membrane
C0412909|T037|HT|977|ICD9CM|Poisoning by other and unspecified drugs and medicinal substances|Poisoning by other and unspecified drugs and medicinal substances
C0161651|T037|PT|977.0|ICD9CM|Poisoning by dietetics|Poisoning by dietetics
C0161651|T037|AB|977.0|ICD9CM|Poisoning-dietetics|Poisoning-dietetics
C0161652|T037|AB|977.1|ICD9CM|Poison-lipotropic drugs|Poison-lipotropic drugs
C0161652|T037|PT|977.1|ICD9CM|Poisoning by lipotropic drugs|Poisoning by lipotropic drugs
C0869440|T037|PT|977.2|ICD9CM|Poisoning by antidotes and chelating agents, not elsewhere classified|Poisoning by antidotes and chelating agents, not elsewhere classified
C0869440|T037|AB|977.2|ICD9CM|Poisoning-antidotes NEC|Poisoning-antidotes NEC
C0161654|T037|AB|977.3|ICD9CM|Poison-alcohol deterrent|Poison-alcohol deterrent
C0161654|T037|PT|977.3|ICD9CM|Poisoning by alcohol deterrents|Poisoning by alcohol deterrents
C0161655|T037|AB|977.4|ICD9CM|Pois-pharmaceut excipien|Pois-pharmaceut excipien
C0161655|T037|PT|977.4|ICD9CM|Poisoning by pharmaceutical excipients|Poisoning by pharmaceutical excipients
C0161656|T037|AB|977.8|ICD9CM|Poison-medicinal agt NEC|Poison-medicinal agt NEC
C0161656|T037|PT|977.8|ICD9CM|Poisoning by other specified drugs and medicinal substances|Poisoning by other specified drugs and medicinal substances
C0013221|T037|AB|977.9|ICD9CM|Poison-medicinal agt NOS|Poison-medicinal agt NOS
C0013221|T037|PT|977.9|ICD9CM|Poisoning by unspecified drug or medicinal substance|Poisoning by unspecified drug or medicinal substance
C0161658|T037|HT|978|ICD9CM|Poisoning by bacterial vaccines|Poisoning by bacterial vaccines
C0161659|T037|PT|978.0|ICD9CM|Poisoning by BCG vaccine|Poisoning by BCG vaccine
C0161659|T037|AB|978.0|ICD9CM|Poisoning-bcg vaccine|Poisoning-bcg vaccine
C0412915|T037|AB|978.1|ICD9CM|Pois-typh/paratyph vacc|Pois-typh/paratyph vacc
C0412915|T037|PT|978.1|ICD9CM|Poisoning by typhoid and paratyphoid vaccine|Poisoning by typhoid and paratyphoid vaccine
C0161661|T037|PT|978.2|ICD9CM|Poisoning by cholera vaccine|Poisoning by cholera vaccine
C0161661|T037|AB|978.2|ICD9CM|Poisoning-cholera vaccin|Poisoning-cholera vaccin
C0161662|T037|PT|978.3|ICD9CM|Poisoning by plague vaccine|Poisoning by plague vaccine
C0161662|T037|AB|978.3|ICD9CM|Poisoning-plague vaccine|Poisoning-plague vaccine
C0161663|T037|PT|978.4|ICD9CM|Poisoning by tetanus vaccine|Poisoning by tetanus vaccine
C0161663|T037|AB|978.4|ICD9CM|Poisoning-tetanus vaccin|Poisoning-tetanus vaccin
C0161664|T037|AB|978.5|ICD9CM|Pois-diphtheria vaccine|Pois-diphtheria vaccine
C0161664|T037|PT|978.5|ICD9CM|Poisoning by diphtheria vaccine|Poisoning by diphtheria vaccine
C0412916|T037|AB|978.6|ICD9CM|Pois-pertussis vaccine|Pois-pertussis vaccine
C0412916|T037|PT|978.6|ICD9CM|Poisoning by pertussis vaccine, including combinations with a pertussis component|Poisoning by pertussis vaccine, including combinations with a pertussis component
C0161666|T037|AB|978.8|ICD9CM|Pois-bact vaccin NEC/NOS|Pois-bact vaccin NEC/NOS
C0161666|T037|PT|978.8|ICD9CM|Poisoning by other and unspecified bacterial vaccines|Poisoning by other and unspecified bacterial vaccines
C0412917|T037|AB|978.9|ICD9CM|Pois-mix bacter vaccines|Pois-mix bacter vaccines
C0412917|T037|PT|978.9|ICD9CM|Poisoning by mixed bacterial vaccines, except combinations with a pertussis component|Poisoning by mixed bacterial vaccines, except combinations with a pertussis component
C0161677|T037|HT|979|ICD9CM|Poisoning by other vaccines and biological substances|Poisoning by other vaccines and biological substances
C0161669|T037|AB|979.0|ICD9CM|Poison-smallpox vaccine|Poison-smallpox vaccine
C0161669|T037|PT|979.0|ICD9CM|Poisoning by smallpox vaccine|Poisoning by smallpox vaccine
C0161670|T037|AB|979.1|ICD9CM|Poison-rabies vaccine|Poison-rabies vaccine
C0161670|T037|PT|979.1|ICD9CM|Poisoning by rabies vaccine|Poisoning by rabies vaccine
C0161671|T037|AB|979.2|ICD9CM|Poison-typhus vaccine|Poison-typhus vaccine
C0161671|T037|PT|979.2|ICD9CM|Poisoning by typhus vaccine|Poisoning by typhus vaccine
C0161672|T037|AB|979.3|ICD9CM|Pois-yellow fever vaccin|Pois-yellow fever vaccin
C0161672|T037|PT|979.3|ICD9CM|Poisoning by yellow fever vaccine|Poisoning by yellow fever vaccine
C0161673|T037|PT|979.4|ICD9CM|Poisoning by measles vaccine|Poisoning by measles vaccine
C0161673|T037|AB|979.4|ICD9CM|Poisoning-measles vaccin|Poisoning-measles vaccin
C0161674|T037|AB|979.5|ICD9CM|Pois-poliomyelit vaccine|Pois-poliomyelit vaccine
C0161674|T037|PT|979.5|ICD9CM|Poisoning by poliomyelitis vaccine|Poisoning by poliomyelitis vaccine
C0161675|T037|AB|979.6|ICD9CM|Pois-viral/rick vacc NEC|Pois-viral/rick vacc NEC
C0161675|T037|PT|979.6|ICD9CM|Poisoning by other and unspecified viral and rickettsial vaccines|Poisoning by other and unspecified viral and rickettsial vaccines
C0161676|T037|AB|979.7|ICD9CM|Poisoning-mixed vaccine|Poisoning-mixed vaccine
C0161677|T037|AB|979.9|ICD9CM|Pois-vaccine/biolog NEC|Pois-vaccine/biolog NEC
C0161677|T037|PT|979.9|ICD9CM|Poisoning by other and unspecified vaccines and biological substances|Poisoning by other and unspecified vaccines and biological substances
C0161678|T037|HT|980|ICD9CM|Toxic effect of alcohol|Toxic effect of alcohol
C0274829|T037|HT|980-989.99|ICD9CM|TOXIC EFFECTS OF SUBSTANCES CHIEFLY NONMEDICINAL AS TO SOURCE|TOXIC EFFECTS OF SUBSTANCES CHIEFLY NONMEDICINAL AS TO SOURCE
C0161679|T037|AB|980.0|ICD9CM|Toxic eff ethyl alcohol|Toxic eff ethyl alcohol
C0161679|T037|PT|980.0|ICD9CM|Toxic effect of ethyl alcohol|Toxic effect of ethyl alcohol
C0161680|T037|AB|980.1|ICD9CM|Toxic eff methyl alcohol|Toxic eff methyl alcohol
C0161680|T037|PT|980.1|ICD9CM|Toxic effect of methyl alcohol|Toxic effect of methyl alcohol
C0161681|T037|AB|980.2|ICD9CM|Toxic eff isopropyl alc|Toxic eff isopropyl alc
C0161681|T037|PT|980.2|ICD9CM|Toxic effect of isopropyl alcohol|Toxic effect of isopropyl alcohol
C0161682|T037|AB|980.3|ICD9CM|Toxic effect fusel oil|Toxic effect fusel oil
C0161682|T037|PT|980.3|ICD9CM|Toxic effect of fusel oil|Toxic effect of fusel oil
C0161683|T037|AB|980.8|ICD9CM|Toxic effect alcohol NEC|Toxic effect alcohol NEC
C0161683|T037|PT|980.8|ICD9CM|Toxic effect of other specified alcohols|Toxic effect of other specified alcohols
C0161678|T037|AB|980.9|ICD9CM|Toxic effect alcohol NOS|Toxic effect alcohol NOS
C0161678|T037|PT|980.9|ICD9CM|Toxic effect of unspecified alcohol|Toxic effect of unspecified alcohol
C0161685|T037|AB|981|ICD9CM|Toxic eff petroleum prod|Toxic eff petroleum prod
C0161685|T037|PT|981|ICD9CM|Toxic effect of petroleum products|Toxic effect of petroleum products
C0274842|T037|HT|982|ICD9CM|Toxic effect of solvents other than petroleum based|Toxic effect of solvents other than petroleum based
C0161687|T037|AB|982.0|ICD9CM|Toxic effect benzene|Toxic effect benzene
C0161687|T037|PT|982.0|ICD9CM|Toxic effect of benzene and homologues|Toxic effect of benzene and homologues
C0392622|T037|AB|982.1|ICD9CM|Toxic eff carbon tetrach|Toxic eff carbon tetrach
C0392622|T037|PT|982.1|ICD9CM|Toxic effect of carbon tetrachloride|Toxic effect of carbon tetrachloride
C0161689|T037|AB|982.2|ICD9CM|Toxic eff carbon disulfi|Toxic eff carbon disulfi
C0161689|T037|PT|982.2|ICD9CM|Toxic effect of carbon disulfide|Toxic effect of carbon disulfide
C0412954|T037|PT|982.3|ICD9CM|Toxic effect of other chlorinated hydrocarbon solvents|Toxic effect of other chlorinated hydrocarbon solvents
C0412954|T037|AB|982.3|ICD9CM|Tx ef cl-hydcarb slv NEC|Tx ef cl-hydcarb slv NEC
C0161691|T037|AB|982.4|ICD9CM|Toxic effect nitroglycol|Toxic effect nitroglycol
C0161691|T037|PT|982.4|ICD9CM|Toxic effect of nitroglycol|Toxic effect of nitroglycol
C0161692|T037|AB|982.8|ICD9CM|Toxic eff nonpetrol solv|Toxic eff nonpetrol solv
C0161692|T037|PT|982.8|ICD9CM|Toxic effect of other nonpetroleum-based solvents|Toxic effect of other nonpetroleum-based solvents
C0161693|T037|HT|983|ICD9CM|Toxic effect of corrosive aromatics, acids, and caustic alkalis|Toxic effect of corrosive aromatics, acids, and caustic alkalis
C0161694|T037|AB|983.0|ICD9CM|Tox eff corrosive aromat|Tox eff corrosive aromat
C0161694|T037|PT|983.0|ICD9CM|Toxic effect of corrosive aromatics|Toxic effect of corrosive aromatics
C0161695|T037|AB|983.1|ICD9CM|Toxic effect acids|Toxic effect acids
C0161695|T037|PT|983.1|ICD9CM|Toxic effect of acids|Toxic effect of acids
C0161696|T037|AB|983.2|ICD9CM|Toxic eff caustic alkali|Toxic eff caustic alkali
C0161696|T037|PT|983.2|ICD9CM|Toxic effect of caustic alkalis|Toxic effect of caustic alkalis
C0375691|T037|AB|983.9|ICD9CM|Toxic effect caustic NOS|Toxic effect caustic NOS
C0375691|T037|PT|983.9|ICD9CM|Toxic effect of caustic, unspecified|Toxic effect of caustic, unspecified
C0023176|T037|HT|984|ICD9CM|Toxic effect of lead and its compounds (including fumes)|Toxic effect of lead and its compounds (including fumes)
C0161699|T037|PT|984.0|ICD9CM|Toxic effect of inorganic lead compounds|Toxic effect of inorganic lead compounds
C0161699|T037|AB|984.0|ICD9CM|Tx eff inorg lead compnd|Tx eff inorg lead compnd
C0161700|T037|AB|984.1|ICD9CM|Tox eff org lead compnd|Tox eff org lead compnd
C0161700|T037|PT|984.1|ICD9CM|Toxic effect of organic lead compounds|Toxic effect of organic lead compounds
C0161701|T037|AB|984.8|ICD9CM|Tox eff lead compnd NEC|Tox eff lead compnd NEC
C0161701|T037|PT|984.8|ICD9CM|Toxic effect of other lead compounds|Toxic effect of other lead compounds
C0023176|T037|AB|984.9|ICD9CM|Tox eff lead compnd NOS|Tox eff lead compnd NOS
C0023176|T037|PT|984.9|ICD9CM|Toxic effect of unspecified lead compound|Toxic effect of unspecified lead compound
C0274869|T037|HT|985|ICD9CM|Toxic effect of other metals|Toxic effect of other metals
C0025427|T037|AB|985.0|ICD9CM|Toxic effect mercury|Toxic effect mercury
C0025427|T037|PT|985.0|ICD9CM|Toxic effect of mercury and its compounds|Toxic effect of mercury and its compounds
C0311375|T037|AB|985.1|ICD9CM|Toxic effect arsenic|Toxic effect arsenic
C0311375|T037|PT|985.1|ICD9CM|Toxic effect of arsenic and its compounds|Toxic effect of arsenic and its compounds
C0412991|T037|AB|985.2|ICD9CM|Toxic effect manganese|Toxic effect manganese
C0412991|T037|PT|985.2|ICD9CM|Toxic effect of manganese and its compounds|Toxic effect of manganese and its compounds
C0412992|T037|AB|985.3|ICD9CM|Toxic effect beryllium|Toxic effect beryllium
C0412992|T037|PT|985.3|ICD9CM|Toxic effect of beryllium and its compounds|Toxic effect of beryllium and its compounds
C0412993|T037|AB|985.4|ICD9CM|Toxic effect antimony|Toxic effect antimony
C0412993|T037|PT|985.4|ICD9CM|Toxic effect of antimony and its compounds|Toxic effect of antimony and its compounds
C0412994|T037|AB|985.5|ICD9CM|Toxic effect cadmium|Toxic effect cadmium
C0412994|T037|PT|985.5|ICD9CM|Toxic effect of cadmium and its compounds|Toxic effect of cadmium and its compounds
C0161708|T037|AB|985.6|ICD9CM|Toxic effect chromium|Toxic effect chromium
C0161708|T037|PT|985.6|ICD9CM|Toxic effect of chromium|Toxic effect of chromium
C0040531|T037|AB|985.8|ICD9CM|Toxic effect metals NEC|Toxic effect metals NEC
C0040531|T037|PT|985.8|ICD9CM|Toxic effect of other specified metals|Toxic effect of other specified metals
C0161709|T037|AB|985.9|ICD9CM|Toxic effect metal NOS|Toxic effect metal NOS
C0161709|T037|PT|985.9|ICD9CM|Toxic effect of unspecified metal|Toxic effect of unspecified metal
C1370867|T037|AB|986|ICD9CM|Tox eff carbon monoxide|Tox eff carbon monoxide
C1370867|T037|PT|986|ICD9CM|Toxic effect of carbon monoxide|Toxic effect of carbon monoxide
C0413000|T037|HT|987|ICD9CM|Toxic effect of other gases, fumes, or vapors|Toxic effect of other gases, fumes, or vapors
C0413005|T037|AB|987.0|ICD9CM|Toxic eff liq petrol gas|Toxic eff liq petrol gas
C0413005|T037|PT|987.0|ICD9CM|Toxic effect of liquefied petroleum gases|Toxic effect of liquefied petroleum gases
C0413004|T037|AB|987.1|ICD9CM|Tox ef hydrocarb gas NEC|Tox ef hydrocarb gas NEC
C0413004|T037|PT|987.1|ICD9CM|Toxic effect of other hydrocarbon gas|Toxic effect of other hydrocarbon gas
C0161713|T037|AB|987.2|ICD9CM|Toxic eff nitrogen oxide|Toxic eff nitrogen oxide
C0161713|T037|PT|987.2|ICD9CM|Toxic effect of nitrogen oxides|Toxic effect of nitrogen oxides
C0161714|T037|AB|987.3|ICD9CM|Toxic eff sulfur dioxide|Toxic eff sulfur dioxide
C0161714|T037|PT|987.3|ICD9CM|Toxic effect of sulfur dioxide|Toxic effect of sulfur dioxide
C0161715|T037|AB|987.4|ICD9CM|Toxic effect freon|Toxic effect freon
C0161715|T037|PT|987.4|ICD9CM|Toxic effect of freon|Toxic effect of freon
C0161716|T037|AB|987.5|ICD9CM|Tox eff lacrimogenic gas|Tox eff lacrimogenic gas
C0161716|T037|PT|987.5|ICD9CM|Toxic effect of lacrimogenic gas|Toxic effect of lacrimogenic gas
C0161717|T037|AB|987.6|ICD9CM|Toxic eff chlorine gas|Toxic eff chlorine gas
C0161717|T037|PT|987.6|ICD9CM|Toxic effect of chlorine gas|Toxic effect of chlorine gas
C0161718|T037|AB|987.7|ICD9CM|Tox eff hydrocyan acd gs|Tox eff hydrocyan acd gs
C0161718|T037|PT|987.7|ICD9CM|Toxic effect of hydrocyanic acid gas|Toxic effect of hydrocyanic acid gas
C0161719|T037|AB|987.8|ICD9CM|Toxic eff gas/vapor NEC|Toxic eff gas/vapor NEC
C0161719|T037|PT|987.8|ICD9CM|Toxic effect of other specified gases, fumes, or vapors|Toxic effect of other specified gases, fumes, or vapors
C0274870|T037|AB|987.9|ICD9CM|Toxic eff gas/vapor NOS|Toxic eff gas/vapor NOS
C0274870|T037|PT|987.9|ICD9CM|Toxic effect of unspecified gas, fume, or vapor|Toxic effect of unspecified gas, fume, or vapor
C0161721|T037|HT|988|ICD9CM|Toxic effect of noxious substances eaten as food|Toxic effect of noxious substances eaten as food
C0161722|T037|AB|988.0|ICD9CM|Toxic eff fish/shellfish|Toxic eff fish/shellfish
C0161722|T037|PT|988.0|ICD9CM|Toxic effect of fish and shellfish eaten as food|Toxic effect of fish and shellfish eaten as food
C0497026|T037|AB|988.1|ICD9CM|Toxic effect mushrooms|Toxic effect mushrooms
C0497026|T037|PT|988.1|ICD9CM|Toxic effect of mushrooms eaten as food|Toxic effect of mushrooms eaten as food
C0040528|T037|AB|988.2|ICD9CM|Tox eff berry/plant NEC|Tox eff berry/plant NEC
C0040528|T037|PT|988.2|ICD9CM|Toxic effect of berries and other plants eaten as food|Toxic effect of berries and other plants eaten as food
C0161723|T037|AB|988.8|ICD9CM|Tox eff noxious food NEC|Tox eff noxious food NEC
C0161723|T037|PT|988.8|ICD9CM|Toxic effect of other specified noxious substances eaten as food|Toxic effect of other specified noxious substances eaten as food
C0161721|T037|AB|988.9|ICD9CM|Tox eff noxious food NOS|Tox eff noxious food NOS
C0161721|T037|PT|988.9|ICD9CM|Toxic effect of unspecified noxious substance eaten as food|Toxic effect of unspecified noxious substance eaten as food
C0161725|T037|HT|989|ICD9CM|Toxic effect of other substances, chiefly nonmedicinal as to source|Toxic effect of other substances, chiefly nonmedicinal as to source
C0161726|T037|AB|989.0|ICD9CM|Toxic effect cyanides|Toxic effect cyanides
C0161726|T037|PT|989.0|ICD9CM|Toxic effect of hydrocyanic acid and cyanides|Toxic effect of hydrocyanic acid and cyanides
C0161727|T037|PT|989.1|ICD9CM|Toxic effect of strychnine and salts|Toxic effect of strychnine and salts
C0161727|T037|AB|989.1|ICD9CM|Toxic effect strychnine|Toxic effect strychnine
C0275016|T037|AB|989.2|ICD9CM|Tox eff chlor hydrocarb|Tox eff chlor hydrocarb
C0275016|T037|PT|989.2|ICD9CM|Toxic effect of chlorinated hydrocarbons|Toxic effect of chlorinated hydrocarbons
C0413040|T037|AB|989.3|ICD9CM|Tox eff organphos/carbam|Tox eff organphos/carbam
C0413040|T037|PT|989.3|ICD9CM|Toxic effect of organophosphate and carbamate|Toxic effect of organophosphate and carbamate
C0302408|T037|AB|989.4|ICD9CM|Toxic eff pesticides NEC|Toxic eff pesticides NEC
C0302408|T037|PT|989.4|ICD9CM|Toxic effect of other pesticides, not elsewhere classified|Toxic effect of other pesticides, not elsewhere classified
C0040533|T037|PT|989.5|ICD9CM|Toxic effect of venom|Toxic effect of venom
C0040533|T037|AB|989.5|ICD9CM|Toxic effect venom|Toxic effect venom
C0274908|T037|AB|989.6|ICD9CM|Toxic eff soap/detergent|Toxic eff soap/detergent
C0274908|T037|PT|989.6|ICD9CM|Toxic effect of soaps and detergents|Toxic effect of soaps and detergents
C0161732|T037|AB|989.7|ICD9CM|Tox eff aflatox/mycotox|Tox eff aflatox/mycotox
C0161732|T037|PT|989.7|ICD9CM|Toxic effect of aflatoxin and other mycotoxin (food contaminants)|Toxic effect of aflatoxin and other mycotoxin (food contaminants)
C0161725|T037|HT|989.8|ICD9CM|Toxic effect of other substances, chiefly nonmedicinal as to source|Toxic effect of other substances, chiefly nonmedicinal as to source
C0375692|T037|AB|989.81|ICD9CM|Toxic effect of asbestos|Toxic effect of asbestos
C0375692|T037|PT|989.81|ICD9CM|Toxic effect of asbestos|Toxic effect of asbestos
C0375693|T037|AB|989.82|ICD9CM|Toxic effect of latex|Toxic effect of latex
C0375693|T037|PT|989.82|ICD9CM|Toxic effect of latex|Toxic effect of latex
C0375694|T037|AB|989.83|ICD9CM|Toxic effect of silicone|Toxic effect of silicone
C0375694|T037|PT|989.83|ICD9CM|Toxic effect of silicone|Toxic effect of silicone
C0375695|T037|AB|989.84|ICD9CM|Toxic effect of tobacco|Toxic effect of tobacco
C0375695|T037|PT|989.84|ICD9CM|Toxic effect of tobacco|Toxic effect of tobacco
C0161725|T037|AB|989.89|ICD9CM|Tox eff nonmed subst NEC|Tox eff nonmed subst NEC
C0161725|T037|PT|989.89|ICD9CM|Toxic effect of other substance, chiefly nonmedicinal as to source, not elsewhere classified|Toxic effect of other substance, chiefly nonmedicinal as to source, not elsewhere classified
C0274829|T037|AB|989.9|ICD9CM|Tox eff nonmed subst NOS|Tox eff nonmed subst NOS
C0274829|T037|PT|989.9|ICD9CM|Toxic effect of unspecified substance, chiefly nonmedicinal as to source|Toxic effect of unspecified substance, chiefly nonmedicinal as to source
C0013679|T037|HT|990-995.99|ICD9CM|OTHER AND UNSPECIFIED EFFECTS OF EXTERNAL CAUSES|OTHER AND UNSPECIFIED EFFECTS OF EXTERNAL CAUSES
C0161734|T037|HT|991|ICD9CM|Effects of reduced temperature|Effects of reduced temperature
C0161735|T037|AB|991.0|ICD9CM|Frostbite of face|Frostbite of face
C0161735|T037|PT|991.0|ICD9CM|Frostbite of face|Frostbite of face
C0161736|T037|AB|991.1|ICD9CM|Frostbite of hand|Frostbite of hand
C0161736|T037|PT|991.1|ICD9CM|Frostbite of hand|Frostbite of hand
C0161737|T037|AB|991.2|ICD9CM|Frostbite of foot|Frostbite of foot
C0161737|T037|PT|991.2|ICD9CM|Frostbite of foot|Frostbite of foot
C0016737|T037|AB|991.3|ICD9CM|Frostbite NEC/NOS|Frostbite NEC/NOS
C0016737|T037|PT|991.3|ICD9CM|Frostbite of other and unspecified sites|Frostbite of other and unspecified sites
C0020941|T037|AB|991.4|ICD9CM|Immersion foot|Immersion foot
C0020941|T037|PT|991.4|ICD9CM|Immersion foot|Immersion foot
C0008058|T047|AB|991.5|ICD9CM|Chilblains|Chilblains
C0008058|T047|PT|991.5|ICD9CM|Chilblains|Chilblains
C0413252|T037|AB|991.6|ICD9CM|Hypothermia|Hypothermia
C0413252|T037|PT|991.6|ICD9CM|Hypothermia|Hypothermia
C0161738|T037|AB|991.8|ICD9CM|Effect reduced temp NEC|Effect reduced temp NEC
C0161738|T037|PT|991.8|ICD9CM|Other specified effects of reduced temperature|Other specified effects of reduced temperature
C0161734|T037|AB|991.9|ICD9CM|Effect reduced temp NOS|Effect reduced temp NOS
C0161734|T037|PT|991.9|ICD9CM|Unspecified effect of reduced temperature|Unspecified effect of reduced temperature
C0274287|T037|HT|992|ICD9CM|Effects of heat and light|Effects of heat and light
C0018844|T037|AB|992.0|ICD9CM|Heat stroke & sunstroke|Heat stroke & sunstroke
C0018844|T037|PT|992.0|ICD9CM|Heat stroke and sunstroke|Heat stroke and sunstroke
C0018845|T037|AB|992.1|ICD9CM|Heat syncope|Heat syncope
C0018845|T037|PT|992.1|ICD9CM|Heat syncope|Heat syncope
C0085592|T037|AB|992.2|ICD9CM|Heat cramps|Heat cramps
C0085592|T037|PT|992.2|ICD9CM|Heat cramps|Heat cramps
C0274288|T037|AB|992.3|ICD9CM|Heat exhaust-anhydrotic|Heat exhaust-anhydrotic
C0274288|T037|PT|992.3|ICD9CM|Heat exhaustion, anhydrotic|Heat exhaustion, anhydrotic
C0152144|T037|AB|992.4|ICD9CM|Heat exhaust-salt deple|Heat exhaust-salt deple
C0152144|T037|PT|992.4|ICD9CM|Heat exhaustion due to salt depletion|Heat exhaustion due to salt depletion
C0018839|T037|AB|992.5|ICD9CM|Heat exhaustion NOS|Heat exhaustion NOS
C0018839|T037|PT|992.5|ICD9CM|Heat exhaustion, unspecified|Heat exhaustion, unspecified
C0152145|T037|AB|992.6|ICD9CM|Heat fatigue, transient|Heat fatigue, transient
C0152145|T037|PT|992.6|ICD9CM|Heat fatigue, transient|Heat fatigue, transient
C0161741|T046|AB|992.7|ICD9CM|Heat edema|Heat edema
C0161741|T046|PT|992.7|ICD9CM|Heat edema|Heat edema
C0161742|T037|AB|992.8|ICD9CM|Heat effect NEC|Heat effect NEC
C0161742|T037|PT|992.8|ICD9CM|Other specified heat effects|Other specified heat effects
C0274287|T037|AB|992.9|ICD9CM|Heat effect NOS|Heat effect NOS
C0274287|T037|PT|992.9|ICD9CM|Unspecified effects of heat and light|Unspecified effects of heat and light
C1306873|T037|HT|993|ICD9CM|Effects of air pressure|Effects of air pressure
C0161744|T037|AB|993.0|ICD9CM|Barotrauma, otitic|Barotrauma, otitic
C0161744|T037|PT|993.0|ICD9CM|Barotrauma, otitic|Barotrauma, otitic
C0161745|T037|AB|993.1|ICD9CM|Barotrauma, sinus|Barotrauma, sinus
C0161745|T037|PT|993.1|ICD9CM|Barotrauma, sinus|Barotrauma, sinus
C0029499|T037|AB|993.2|ICD9CM|Eff high altitud NEC/NOS|Eff high altitud NEC/NOS
C0029499|T037|PT|993.2|ICD9CM|Other and unspecified effects of high altitude|Other and unspecified effects of high altitude
C0011119|T047|AB|993.3|ICD9CM|Caisson disease|Caisson disease
C0011119|T047|PT|993.3|ICD9CM|Caisson disease|Caisson disease
C0005700|T037|AB|993.4|ICD9CM|Eff air press by explos|Eff air press by explos
C0005700|T037|PT|993.4|ICD9CM|Effects of air pressure caused by explosion|Effects of air pressure caused by explosion
C0161747|T037|AB|993.8|ICD9CM|Effect air pressure NEC|Effect air pressure NEC
C0161747|T037|PT|993.8|ICD9CM|Other specified effects of air pressure|Other specified effects of air pressure
C0161748|T037|AB|993.9|ICD9CM|Effect air pressure NOS|Effect air pressure NOS
C0161748|T037|PT|993.9|ICD9CM|Unspecified effect of air pressure|Unspecified effect of air pressure
C0013679|T037|HT|994|ICD9CM|Effects of other external causes|Effects of other external causes
C0023702|T037|AB|994.0|ICD9CM|Effects of lightning|Effects of lightning
C0023702|T037|PT|994.0|ICD9CM|Effects of lightning|Effects of lightning
C0013143|T037|PT|994.1|ICD9CM|Drowning and nonfatal submersion|Drowning and nonfatal submersion
C0013143|T037|AB|994.1|ICD9CM|Drowning/nonfatal submer|Drowning/nonfatal submer
C0311274|T037|AB|994.2|ICD9CM|Effects of hunger|Effects of hunger
C0311274|T037|PT|994.2|ICD9CM|Effects of hunger|Effects of hunger
C0013680|T047|AB|994.3|ICD9CM|Effects of thirst|Effects of thirst
C0013680|T047|PT|994.3|ICD9CM|Effects of thirst|Effects of thirst
C0161749|T037|PT|994.4|ICD9CM|Exhaustion due to exposure|Exhaustion due to exposure
C0161749|T037|AB|994.4|ICD9CM|Exhaustion-exposure|Exhaustion-exposure
C0161750|T037|PT|994.5|ICD9CM|Exhaustion due to excessive exertion|Exhaustion due to excessive exertion
C0161750|T037|AB|994.5|ICD9CM|Exhaustion-excess exert|Exhaustion-excess exert
C0026603|T047|AB|994.6|ICD9CM|Motion sickness|Motion sickness
C0026603|T047|PT|994.6|ICD9CM|Motion sickness|Motion sickness
C0161751|T037|PT|994.7|ICD9CM|Asphyxiation and strangulation|Asphyxiation and strangulation
C0161751|T037|AB|994.7|ICD9CM|Asphyxiation/strangulat|Asphyxiation/strangulat
C0161752|T037|AB|994.8|ICD9CM|Effects electric current|Effects electric current
C0161752|T037|PT|994.8|ICD9CM|Electrocution and nonfatal effects of electric current|Electrocution and nonfatal effects of electric current
C2240397|T037|AB|994.9|ICD9CM|Effect external caus NEC|Effect external caus NEC
C2240397|T037|PT|994.9|ICD9CM|Other effects of external causes|Other effects of external causes
C0302409|T037|HT|995|ICD9CM|Certain adverse effects not elsewhere classified|Certain adverse effects not elsewhere classified
C3161335|T037|AB|995.0|ICD9CM|Other anaphylactic react|Other anaphylactic react
C3161335|T037|PT|995.0|ICD9CM|Other anaphylactic reaction|Other anaphylactic reaction
C0877771|T046|AB|995.1|ICD9CM|Angioneurotic edema|Angioneurotic edema
C0877771|T046|PT|995.1|ICD9CM|Angioneurotic edema, not elsewhere classified|Angioneurotic edema, not elsewhere classified
C2921193|T037|HT|995.2|ICD9CM|Other and unspecified adverse effect of drug, medicinal and biological substance|Other and unspecified adverse effect of drug, medicinal and biological substance
C1719666|T046|AB|995.20|ICD9CM|Adv eff med/biol sub NOS|Adv eff med/biol sub NOS
C1719666|T046|PT|995.20|ICD9CM|Unspecified adverse effect of unspecified drug, medicinal and biological substance|Unspecified adverse effect of unspecified drug, medicinal and biological substance
C0003907|T047|PT|995.21|ICD9CM|Arthus phenomenon|Arthus phenomenon
C0003907|T047|AB|995.21|ICD9CM|Arthus phenomenon|Arthus phenomenon
C1719667|T046|AB|995.22|ICD9CM|Adv eff anesthesia NOS|Adv eff anesthesia NOS
C1719667|T046|PT|995.22|ICD9CM|Unspecified adverse effect of anesthesia|Unspecified adverse effect of anesthesia
C1719668|T046|AB|995.23|ICD9CM|Adverse eff insulin NOS|Adverse eff insulin NOS
C1719668|T046|PT|995.23|ICD9CM|Unspecified adverse effect of insulin|Unspecified adverse effect of insulin
C2712382|T037|AB|995.24|ICD9CM|Fail mod sedate dur proc|Fail mod sedate dur proc
C2712382|T037|PT|995.24|ICD9CM|Failed moderate sedation during procedure|Failed moderate sedation during procedure
C1719669|T047|AB|995.27|ICD9CM|Drug allergy NEC|Drug allergy NEC
C1719669|T047|PT|995.27|ICD9CM|Other drug allergy|Other drug allergy
C1719670|T046|AB|995.29|ICD9CM|Adv eff med/biol NEC/NOS|Adv eff med/biol NEC/NOS
C1719670|T046|PT|995.29|ICD9CM|Unspecified adverse effect of other drug, medicinal and biological substance|Unspecified adverse effect of other drug, medicinal and biological substance
C0700625|T047|AB|995.3|ICD9CM|Allergy, unspecified|Allergy, unspecified
C0700625|T047|PT|995.3|ICD9CM|Allergy, unspecified, not elsewhere classified|Allergy, unspecified, not elsewhere classified
C0812420|T037|AB|995.4|ICD9CM|Shock due to anesthesia|Shock due to anesthesia
C0812420|T037|PT|995.4|ICD9CM|Shock due to anesthesia, not elsewhere classified|Shock due to anesthesia, not elsewhere classified
C0008060|T048|HT|995.5|ICD9CM|Child maltreatment syndrome|Child maltreatment syndrome
C0008060|T048|AB|995.50|ICD9CM|Child abuse NOS|Child abuse NOS
C0008060|T048|PT|995.50|ICD9CM|Child abuse, unspecified|Child abuse, unspecified
C0375699|T048|PT|995.51|ICD9CM|Child emotional/psychological abuse|Child emotional/psychological abuse
C0375699|T048|AB|995.51|ICD9CM|Child emotnl/psych abuse|Child emotnl/psych abuse
C0375700|T033|PT|995.52|ICD9CM|Child neglect (nutritional)|Child neglect (nutritional)
C0375700|T033|AB|995.52|ICD9CM|Child neglect-nutrition|Child neglect-nutrition
C0008062|T048|AB|995.53|ICD9CM|Child sexual abuse|Child sexual abuse
C0008062|T048|PT|995.53|ICD9CM|Child sexual abuse|Child sexual abuse
C0236861|T033|AB|995.54|ICD9CM|Child physical abuse|Child physical abuse
C0236861|T033|PT|995.54|ICD9CM|Child physical abuse|Child physical abuse
C0686721|T037|PT|995.55|ICD9CM|Shaken baby syndrome|Shaken baby syndrome
C0686721|T037|AB|995.55|ICD9CM|Shaken infant syndrome|Shaken infant syndrome
C0375702|T037|AB|995.59|ICD9CM|Child abuse/neglect NEC|Child abuse/neglect NEC
C0375702|T037|PT|995.59|ICD9CM|Other child abuse and neglect|Other child abuse and neglect
C0685898|T047|HT|995.6|ICD9CM|Anaphylactic reaction due to food|Anaphylactic reaction due to food
C0375703|T037|PT|995.60|ICD9CM|Anaphylactic reaction due to unspecified food|Anaphylactic reaction due to unspecified food
C0375703|T037|AB|995.60|ICD9CM|Anphylct react food NOS|Anphylct react food NOS
C0859855|T046|PT|995.61|ICD9CM|Anaphylactic reaction due to peanuts|Anaphylactic reaction due to peanuts
C0859855|T046|AB|995.61|ICD9CM|Anphylct react peanuts|Anphylct react peanuts
C0859856|T046|PT|995.62|ICD9CM|Anaphylactic reaction due to crustaceans|Anaphylactic reaction due to crustaceans
C0859856|T046|AB|995.62|ICD9CM|Anphylct react crstacns|Anphylct react crstacns
C0859857|T046|PT|995.63|ICD9CM|Anaphylactic reaction due to fruits and vegetables|Anaphylactic reaction due to fruits and vegetables
C0859857|T046|AB|995.63|ICD9CM|Anphylct react frts veg|Anphylct react frts veg
C0375707|T046|PT|995.64|ICD9CM|Anaphylactic reaction due to tree nuts and seeds|Anaphylactic reaction due to tree nuts and seeds
C0375707|T046|AB|995.64|ICD9CM|Anphyl react tr nts seed|Anphyl react tr nts seed
C0859858|T046|PT|995.65|ICD9CM|Anaphylactic reaction due to fish|Anaphylactic reaction due to fish
C0859858|T046|AB|995.65|ICD9CM|Anphylct reaction fish|Anphylct reaction fish
C0859859|T046|PT|995.66|ICD9CM|Anaphylactic reaction due to food additives|Anaphylactic reaction due to food additives
C0859859|T046|AB|995.66|ICD9CM|Anphylct react food addv|Anphylct react food addv
C0859860|T046|PT|995.67|ICD9CM|Anaphylactic reaction due to milk products|Anaphylactic reaction due to milk products
C0859860|T046|AB|995.67|ICD9CM|Anphylct react milk prod|Anphylct react milk prod
C0859861|T046|PT|995.68|ICD9CM|Anaphylactic reaction due to eggs|Anaphylactic reaction due to eggs
C0859861|T046|AB|995.68|ICD9CM|Anphylct reaction eggs|Anphylct reaction eggs
C3161345|T046|PT|995.69|ICD9CM|Anaphylactic reaction due to other specified food|Anaphylactic reaction due to other specified food
C3161345|T046|AB|995.69|ICD9CM|Anphyl react oth sp food|Anphyl react oth sp food
C0869098|T037|AB|995.7|ICD9CM|Adverse food react NEC|Adverse food react NEC
C0869098|T037|PT|995.7|ICD9CM|Other adverse food reactions, not elsewhere classified|Other adverse food reactions, not elsewhere classified
C1561653|T037|HT|995.8|ICD9CM|Other specified adverse effects, not elsewhere classified|Other specified adverse effects, not elsewhere classified
C0375714|T037|AB|995.80|ICD9CM|Adult maltreatment NOS|Adult maltreatment NOS
C0375714|T037|PT|995.80|ICD9CM|Adult maltreatment, unspecified|Adult maltreatment, unspecified
C0236859|T037|AB|995.81|ICD9CM|Adult physical abuse|Adult physical abuse
C0236859|T037|PT|995.81|ICD9CM|Adult physical abuse|Adult physical abuse
C0375715|T048|PT|995.82|ICD9CM|Adult emotional/psychological abuse|Adult emotional/psychological abuse
C0375715|T048|AB|995.82|ICD9CM|Adult emotnl/psych abuse|Adult emotnl/psych abuse
C0236860|T048|AB|995.83|ICD9CM|Adult sexual abuse|Adult sexual abuse
C0236860|T048|PT|995.83|ICD9CM|Adult sexual abuse|Adult sexual abuse
C0375716|T033|PT|995.84|ICD9CM|Adult neglect (nutritional)|Adult neglect (nutritional)
C0375716|T033|AB|995.84|ICD9CM|Adult neglect-nutrition|Adult neglect-nutrition
C0375717|T048|AB|995.85|ICD9CM|Oth adult abuse/neglect|Oth adult abuse/neglect
C0375717|T048|PT|995.85|ICD9CM|Other adult abuse and neglect|Other adult abuse and neglect
C0024591|T047|AB|995.86|ICD9CM|Malignant hyperthermia|Malignant hyperthermia
C0024591|T047|PT|995.86|ICD9CM|Malignant hyperthermia|Malignant hyperthermia
C1561653|T037|AB|995.89|ICD9CM|Adverse effect NEC|Adverse effect NEC
C1561653|T037|PT|995.89|ICD9CM|Other specified adverse effects, not elsewhere classified|Other specified adverse effects, not elsewhere classified
C0242966|T047|HT|995.9|ICD9CM|Systemic inflammatory response syndrome (SIRS)|Systemic inflammatory response syndrome (SIRS)
C0242966|T047|AB|995.90|ICD9CM|SIRS, NOS|SIRS, NOS
C0242966|T047|PT|995.90|ICD9CM|Systemic inflammatory response syndrome, unspecified|Systemic inflammatory response syndrome, unspecified
C0243026|T047|PT|995.91|ICD9CM|Sepsis|Sepsis
C0243026|T047|AB|995.91|ICD9CM|Sepsis|Sepsis
C1719672|T047|PT|995.92|ICD9CM|Severe sepsis|Severe sepsis
C1719672|T047|AB|995.92|ICD9CM|Severe sepsis|Severe sepsis
C1719676|T047|AB|995.93|ICD9CM|SIRS-noninf w/o ac or ds|SIRS-noninf w/o ac or ds
C1719676|T047|PT|995.93|ICD9CM|Systemic inflammatory response syndrome due to noninfectious process without acute organ dysfunction|Systemic inflammatory response syndrome due to noninfectious process without acute organ dysfunction
C1719677|T037|AB|995.94|ICD9CM|SIRS-noninf w ac org dys|SIRS-noninf w ac org dys
C1719677|T037|PT|995.94|ICD9CM|Systemic inflammatory response syndrome due to noninfectious process with acute organ dysfunction|Systemic inflammatory response syndrome due to noninfectious process with acute organ dysfunction
C0496137|T046|HT|996|ICD9CM|Complications peculiar to certain specified procedures|Complications peculiar to certain specified procedures
C0869272|T046|HT|996-999.99|ICD9CM|COMPLICATIONS OF SURGICAL AND MEDICAL CARE, NOT ELSEWHERE CLASSIFIED|COMPLICATIONS OF SURGICAL AND MEDICAL CARE, NOT ELSEWHERE CLASSIFIED
C0274323|T046|HT|996.0|ICD9CM|Mechanical complication of cardiac device, implant, and graft|Mechanical complication of cardiac device, implant, and graft
C0274323|T046|AB|996.00|ICD9CM|Malfunc card dev/grf NOS|Malfunc card dev/grf NOS
C0274323|T046|PT|996.00|ICD9CM|Mechanical complication of unspecified cardiac device, implant, and graft|Mechanical complication of unspecified cardiac device, implant, and graft
C0161759|T037|AB|996.01|ICD9CM|Malfunc cardiac pacemake|Malfunc cardiac pacemake
C0161759|T037|PT|996.01|ICD9CM|Mechanical complication due to cardiac pacemaker (electrode)|Mechanical complication due to cardiac pacemaker (electrode)
C0161760|T046|AB|996.02|ICD9CM|Malfunc prosth hrt valve|Malfunc prosth hrt valve
C0161760|T046|PT|996.02|ICD9CM|Mechanical complication due to heart valve prosthesis|Mechanical complication due to heart valve prosthesis
C0161761|T037|AB|996.03|ICD9CM|Malfunc coron bypass grf|Malfunc coron bypass grf
C0161761|T037|PT|996.03|ICD9CM|Mechanical complication due to coronary bypass graft|Mechanical complication due to coronary bypass graft
C0375718|T046|AB|996.04|ICD9CM|Mch cmp autm mplnt dfbrl|Mch cmp autm mplnt dfbrl
C0375718|T046|PT|996.04|ICD9CM|Mechanical complication of automatic implantable cardiac defibrillator|Mechanical complication of automatic implantable cardiac defibrillator
C0161762|T046|AB|996.09|ICD9CM|Malfunc card dev/grf NEC|Malfunc card dev/grf NEC
C0161762|T046|PT|996.09|ICD9CM|Other mechanical complication of cardiac device, implant, and graft|Other mechanical complication of cardiac device, implant, and graft
C0161763|T046|AB|996.1|ICD9CM|Malfunc vasc device/graf|Malfunc vasc device/graf
C0161763|T046|PT|996.1|ICD9CM|Mechanical complication of other vascular device, implant, and graft|Mechanical complication of other vascular device, implant, and graft
C0274338|T037|AB|996.2|ICD9CM|Malfun neuro device/graf|Malfun neuro device/graf
C0274338|T037|PT|996.2|ICD9CM|Mechanical complication of nervous system device, implant, and graft|Mechanical complication of nervous system device, implant, and graft
C0274344|T046|HT|996.3|ICD9CM|Mechanical complication of genitourinary device, implant, and graft|Mechanical complication of genitourinary device, implant, and graft
C0274344|T046|AB|996.30|ICD9CM|Malfunc gu dev/graft NOS|Malfunc gu dev/graft NOS
C0274344|T046|PT|996.30|ICD9CM|Mechanical complication of unspecified genitourinary device, implant, and graft|Mechanical complication of unspecified genitourinary device, implant, and graft
C0161767|T046|AB|996.31|ICD9CM|Malfunc urethral cath|Malfunc urethral cath
C0161767|T046|PT|996.31|ICD9CM|Mechanical complication due to urethral (indwelling) catheter|Mechanical complication due to urethral (indwelling) catheter
C0161768|T046|AB|996.32|ICD9CM|Malfunction iud|Malfunction iud
C0161768|T046|PT|996.32|ICD9CM|Mechanical complication due to intrauterine contraceptive device|Mechanical complication due to intrauterine contraceptive device
C0161769|T037|AB|996.39|ICD9CM|Malfunc gu dev/graft NEC|Malfunc gu dev/graft NEC
C0161769|T037|PT|996.39|ICD9CM|Other mechanical complication of genitourinary device, implant, and graft|Other mechanical complication of genitourinary device, implant, and graft
C0161770|T046|HT|996.4|ICD9CM|Mechanical complication of internal orthopedic device, implant, and graft|Mechanical complication of internal orthopedic device, implant, and graft
C1561654|T046|AB|996.40|ICD9CM|Cmp int orth dev/gft NOS|Cmp int orth dev/gft NOS
C1561654|T046|PT|996.40|ICD9CM|Unspecified mechanical complication of internal orthopedic device, implant, and graft|Unspecified mechanical complication of internal orthopedic device, implant, and graft
C1561655|T046|AB|996.41|ICD9CM|Mech loosening pros jt|Mech loosening pros jt
C1561655|T046|PT|996.41|ICD9CM|Mechanical loosening of prosthetic joint|Mechanical loosening of prosthetic joint
C0410807|T033|AB|996.42|ICD9CM|Dislocate prosthetic jt|Dislocate prosthetic jt
C0410807|T033|PT|996.42|ICD9CM|Dislocation of prosthetic joint|Dislocation of prosthetic joint
C2712383|T037|AB|996.43|ICD9CM|Broke prosthtc jt implnt|Broke prosthtc jt implnt
C2712383|T037|PT|996.43|ICD9CM|Broken prosthetic joint implant|Broken prosthetic joint implant
C1561661|T046|PT|996.44|ICD9CM|Peri-prosthetic fracture around prosthetic joint|Peri-prosthetic fracture around prosthetic joint
C1561661|T046|AB|996.44|ICD9CM|Periprosthetc fx-pros jt|Periprosthetc fx-pros jt
C0948364|T046|PT|996.45|ICD9CM|Peri-prosthetic osteolysis|Peri-prosthetic osteolysis
C0948364|T046|AB|996.45|ICD9CM|Periprosthetc osteolysis|Periprosthetc osteolysis
C2711887|T046|PT|996.46|ICD9CM|Articular bearing surface wear of prosthetic joint|Articular bearing surface wear of prosthetic joint
C2711887|T046|AB|996.46|ICD9CM|Articular wear prosth jt|Articular wear prosth jt
C1561664|T046|AB|996.47|ICD9CM|Mech com pros jt implant|Mech com pros jt implant
C1561664|T046|PT|996.47|ICD9CM|Other mechanical complication of prosthetic joint implant|Other mechanical complication of prosthetic joint implant
C1561666|T046|AB|996.49|ICD9CM|Mech com orth dev NEC|Mech com orth dev NEC
C1561666|T046|PT|996.49|ICD9CM|Other mechanical complication of other internal orthopedic device, implant, and graft|Other mechanical complication of other internal orthopedic device, implant, and graft
C0161771|T037|HT|996.5|ICD9CM|Mechanical complication of other specified prosthetic device, implant, and graft|Mechanical complication of other specified prosthetic device, implant, and graft
C0274354|T046|AB|996.51|ICD9CM|Corneal grft malfunction|Corneal grft malfunction
C0274354|T046|PT|996.51|ICD9CM|Mechanical complication due to corneal graft|Mechanical complication due to corneal graft
C0302411|T046|PT|996.52|ICD9CM|Mechanical complication due to graft of other tissue, not elsewhere classified|Mechanical complication due to graft of other tissue, not elsewhere classified
C0302411|T046|AB|996.52|ICD9CM|Oth tissue graft malfunc|Oth tissue graft malfunc
C0274356|T046|AB|996.53|ICD9CM|Lens prosthesis malfunc|Lens prosthesis malfunc
C0274356|T046|PT|996.53|ICD9CM|Mechanical complication due to ocular lens prosthesis|Mechanical complication due to ocular lens prosthesis
C0274357|T046|AB|996.54|ICD9CM|Breast prosth malfunc|Breast prosth malfunc
C0274357|T046|PT|996.54|ICD9CM|Mechanical complication due to breast prosthesis|Mechanical complication due to breast prosthesis
C0695254|T046|AB|996.55|ICD9CM|Comp-artificial skin grf|Comp-artificial skin grf
C0695254|T046|PT|996.55|ICD9CM|Mechanical complication due to artificial skin graft and decellularized allodermis|Mechanical complication due to artificial skin graft and decellularized allodermis
C0695255|T046|AB|996.56|ICD9CM|Comp-periton dialys cath|Comp-periton dialys cath
C0695255|T046|PT|996.56|ICD9CM|Mechanical complication due to peritoneal dialysis catheter|Mechanical complication due to peritoneal dialysis catheter
C2228890|T037|AB|996.57|ICD9CM|Complcation-insulin pump|Complcation-insulin pump
C2228890|T037|PT|996.57|ICD9CM|Mechanical complication due to insulin pump|Mechanical complication due to insulin pump
C0302412|T046|AB|996.59|ICD9CM|Malfunc oth device/graft|Malfunc oth device/graft
C0302412|T046|PT|996.59|ICD9CM|Mechanical complication due to other implant and internal device, not elsewhere classified|Mechanical complication due to other implant and internal device, not elsewhere classified
C0161777|T047|HT|996.6|ICD9CM|Infection and inflammatory reaction due to internal prosthetic device, implant, and graft|Infection and inflammatory reaction due to internal prosthetic device, implant, and graft
C0161778|T047|PT|996.60|ICD9CM|Infection and inflammatory reaction due to unspecified device, implant, and graft|Infection and inflammatory reaction due to unspecified device, implant, and graft
C0161778|T047|AB|996.60|ICD9CM|Reaction-unsp devic/grft|Reaction-unsp devic/grft
C0161779|T047|PT|996.61|ICD9CM|Infection and inflammatory reaction due to cardiac device, implant, and graft|Infection and inflammatory reaction due to cardiac device, implant, and graft
C0161779|T047|AB|996.61|ICD9CM|React-cardiac dev/graft|React-cardiac dev/graft
C0161780|T047|PT|996.62|ICD9CM|Infection and inflammatory reaction due to other vascular device, implant, and graft|Infection and inflammatory reaction due to other vascular device, implant, and graft
C0161780|T047|AB|996.62|ICD9CM|React-oth vasc dev/graft|React-oth vasc dev/graft
C0161781|T046|PT|996.63|ICD9CM|Infection and inflammatory reaction due to nervous system device, implant, and graft|Infection and inflammatory reaction due to nervous system device, implant, and graft
C0161781|T046|AB|996.63|ICD9CM|React-nerv sys dev/graft|React-nerv sys dev/graft
C0161782|T047|PT|996.64|ICD9CM|Infection and inflammatory reaction due to indwelling urinary catheter|Infection and inflammatory reaction due to indwelling urinary catheter
C0161782|T047|AB|996.64|ICD9CM|React-indwell urin cath|React-indwell urin cath
C0161783|T047|PT|996.65|ICD9CM|Infection and inflammatory reaction due to other genitourinary device, implant, and graft|Infection and inflammatory reaction due to other genitourinary device, implant, and graft
C0161783|T047|AB|996.65|ICD9CM|React-oth genitourin dev|React-oth genitourin dev
C0161784|T047|PT|996.66|ICD9CM|Infection and inflammatory reaction due to internal joint prosthesis|Infection and inflammatory reaction due to internal joint prosthesis
C0161784|T047|AB|996.66|ICD9CM|React-inter joint prost|React-inter joint prost
C0161785|T047|PT|996.67|ICD9CM|Infection and inflammatory reaction due to other internal orthopedic device, implant, and graft|Infection and inflammatory reaction due to other internal orthopedic device, implant, and graft
C0161785|T047|AB|996.67|ICD9CM|React-oth int ortho dev|React-oth int ortho dev
C0695256|T046|PT|996.68|ICD9CM|Infection and inflammatory reaction due to peritoneal dialysis catheter|Infection and inflammatory reaction due to peritoneal dialysis catheter
C0695256|T046|AB|996.68|ICD9CM|React-periton dialy cath|React-periton dialy cath
C0161786|T046|PT|996.69|ICD9CM|Infection and inflammatory reaction due to other internal prosthetic device, implant, and graft|Infection and inflammatory reaction due to other internal prosthetic device, implant, and graft
C0161786|T046|AB|996.69|ICD9CM|React-int pros devic NEC|React-int pros devic NEC
C0161787|T046|HT|996.7|ICD9CM|Other complications of internal (biological) (synthetic) prosthetic device, implant, and graft|Other complications of internal (biological) (synthetic) prosthetic device, implant, and graft
C0161788|T047|AB|996.70|ICD9CM|Comp-unsp device/graft|Comp-unsp device/graft
C0161788|T047|PT|996.70|ICD9CM|Other complications due to unspecified device, implant, and graft|Other complications due to unspecified device, implant, and graft
C0161789|T047|AB|996.71|ICD9CM|Comp-heart valve prosth|Comp-heart valve prosth
C0161789|T047|PT|996.71|ICD9CM|Other complications due to heart valve prosthesis|Other complications due to heart valve prosthesis
C0161790|T047|AB|996.72|ICD9CM|Comp-oth cardiac device|Comp-oth cardiac device
C0161790|T047|PT|996.72|ICD9CM|Other complications due to other cardiac device, implant, and graft|Other complications due to other cardiac device, implant, and graft
C0161791|T047|AB|996.73|ICD9CM|Comp-ren dialys dev/grft|Comp-ren dialys dev/grft
C0161791|T047|PT|996.73|ICD9CM|Other complications due to renal dialysis device, implant, and graft|Other complications due to renal dialysis device, implant, and graft
C0161792|T047|AB|996.74|ICD9CM|Comp-oth vasc dev/graft|Comp-oth vasc dev/graft
C0161792|T047|PT|996.74|ICD9CM|Other complications due to other vascular device, implant, and graft|Other complications due to other vascular device, implant, and graft
C0840880|T046|AB|996.75|ICD9CM|Comp-nerv sys dev/graft|Comp-nerv sys dev/graft
C0840880|T046|PT|996.75|ICD9CM|Other complications due to nervous system device, implant, and graft|Other complications due to nervous system device, implant, and graft
C0161794|T047|AB|996.76|ICD9CM|Comp-genitourin dev/grft|Comp-genitourin dev/grft
C0161794|T047|PT|996.76|ICD9CM|Other complications due to genitourinary device, implant, and graft|Other complications due to genitourinary device, implant, and graft
C0161795|T047|AB|996.77|ICD9CM|Comp-internal joint pros|Comp-internal joint pros
C0161795|T047|PT|996.77|ICD9CM|Other complications due to internal joint prosthesis|Other complications due to internal joint prosthesis
C0161796|T047|AB|996.78|ICD9CM|Comp-oth int ortho devic|Comp-oth int ortho devic
C0161796|T047|PT|996.78|ICD9CM|Other complications due to other internal orthopedic device, implant, and graft|Other complications due to other internal orthopedic device, implant, and graft
C0161797|T047|AB|996.79|ICD9CM|Comp-int prost devic NEC|Comp-int prost devic NEC
C0161797|T047|PT|996.79|ICD9CM|Other complications due to other internal prosthetic device, implant, and graft|Other complications due to other internal prosthetic device, implant, and graft
C0009568|T046|HT|996.8|ICD9CM|Complications of transplanted organ|Complications of transplanted organ
C0375720|T046|AB|996.80|ICD9CM|Comp organ transplnt NOS|Comp organ transplnt NOS
C0375720|T046|PT|996.80|ICD9CM|Complications of transplanted organ, unspecified|Complications of transplanted organ, unspecified
C1261281|T046|AB|996.81|ICD9CM|Compl kidney transplant|Compl kidney transplant
C1261281|T046|PT|996.81|ICD9CM|Complications of transplanted kidney|Complications of transplanted kidney
C1261282|T046|AB|996.82|ICD9CM|Compl liver transplant|Compl liver transplant
C1261282|T046|PT|996.82|ICD9CM|Complications of transplanted liver|Complications of transplanted liver
C0340529|T046|AB|996.83|ICD9CM|Compl heart transplant|Compl heart transplant
C0340529|T046|PT|996.83|ICD9CM|Complications of transplanted heart|Complications of transplanted heart
C0161801|T046|AB|996.84|ICD9CM|Compl lung transplant|Compl lung transplant
C0161801|T046|PT|996.84|ICD9CM|Complications of transplanted lung|Complications of transplanted lung
C0161802|T046|AB|996.85|ICD9CM|Compl marrow transplant|Compl marrow transplant
C0161802|T046|PT|996.85|ICD9CM|Complications of transplanted bone marrow|Complications of transplanted bone marrow
C0161803|T046|AB|996.86|ICD9CM|Compl pancreas transplnt|Compl pancreas transplnt
C0161803|T046|PT|996.86|ICD9CM|Complications of transplanted pancreas|Complications of transplanted pancreas
C0274370|T046|AB|996.87|ICD9CM|Comp intestine transplnt|Comp intestine transplnt
C0274370|T046|PT|996.87|ICD9CM|Complications of transplanted intestine|Complications of transplanted intestine
C3251587|T046|AB|996.88|ICD9CM|Comp tp organ-stem cell|Comp tp organ-stem cell
C3251587|T046|PT|996.88|ICD9CM|Complications of transplanted organ, stem cell|Complications of transplanted organ, stem cell
C0161804|T046|AB|996.89|ICD9CM|Comp oth organ transplnt|Comp oth organ transplnt
C0161804|T046|PT|996.89|ICD9CM|Complications of other specified transplanted organ|Complications of other specified transplanted organ
C0161805|T047|HT|996.9|ICD9CM|Complications of reattached extremity or body part|Complications of reattached extremity or body part
C1439344|T037|AB|996.90|ICD9CM|Comp reattach extrem NOS|Comp reattach extrem NOS
C1439344|T037|PT|996.90|ICD9CM|Complications of unspecified reattached extremity|Complications of unspecified reattached extremity
C0161807|T047|AB|996.91|ICD9CM|Compl reattached forearm|Compl reattached forearm
C0161807|T047|PT|996.91|ICD9CM|Complications of reattached forearm|Complications of reattached forearm
C0161808|T046|AB|996.92|ICD9CM|Compl reattached hand|Compl reattached hand
C0161808|T046|PT|996.92|ICD9CM|Complications of reattached hand|Complications of reattached hand
C0274372|T046|AB|996.93|ICD9CM|Compl reattached finger|Compl reattached finger
C0274372|T046|PT|996.93|ICD9CM|Complications of reattached finger(s)|Complications of reattached finger(s)
C0489974|T037|AB|996.94|ICD9CM|Compl reattached arm NEC|Compl reattached arm NEC
C0489974|T037|PT|996.94|ICD9CM|Complications of reattached upper extremity, other and unspecified|Complications of reattached upper extremity, other and unspecified
C0274373|T046|AB|996.95|ICD9CM|Compl reattached foot|Compl reattached foot
C0274373|T046|PT|996.95|ICD9CM|Complication of reattached foot and toe(s)|Complication of reattached foot and toe(s)
C2240398|T046|AB|996.96|ICD9CM|Compl reattached leg NEC|Compl reattached leg NEC
C2240398|T046|PT|996.96|ICD9CM|Complication of reattached lower extremity, other and unspecified|Complication of reattached lower extremity, other and unspecified
C0161813|T037|AB|996.99|ICD9CM|Compl reattach part NEC|Compl reattach part NEC
C0161813|T037|PT|996.99|ICD9CM|Complication of other specified reattached body part|Complication of other specified reattached body part
C0868769|T037|HT|997|ICD9CM|Complications affecting specified body systems, not elsewhere classified|Complications affecting specified body systems, not elsewhere classified
C0302414|T037|HT|997.0|ICD9CM|Central nervous system complications, not elsewhere classified|Central nervous system complications, not elsewhere classified
C0235029|T046|AB|997.00|ICD9CM|Nervous syst complc NOS|Nervous syst complc NOS
C0235029|T046|PT|997.00|ICD9CM|Nervous system complication, unspecified|Nervous system complication, unspecified
C0161815|T046|PT|997.01|ICD9CM|Central nervous system complication|Central nervous system complication
C0161815|T046|AB|997.01|ICD9CM|Surg complication - cns|Surg complication - cns
C0375722|T047|AB|997.02|ICD9CM|Iatrogen CV infarc/hmrhg|Iatrogen CV infarc/hmrhg
C0375722|T047|PT|997.02|ICD9CM|Iatrogenic cerebrovascular infarction or hemorrhage|Iatrogenic cerebrovascular infarction or hemorrhage
C0375723|T046|PT|997.09|ICD9CM|Other nervous system complications|Other nervous system complications
C0375723|T046|AB|997.09|ICD9CM|Surg comp nerv systm NEC|Surg comp nerv systm NEC
C0549147|T046|PT|997.1|ICD9CM|Cardiac complications, not elsewhere classified|Cardiac complications, not elsewhere classified
C0549147|T046|AB|997.1|ICD9CM|Surg compl-heart|Surg compl-heart
C0877738|T046|PT|997.2|ICD9CM|Peripheral vascular complications, not elsewhere classified|Peripheral vascular complications, not elsewhere classified
C0877738|T046|AB|997.2|ICD9CM|Surg comp-peri vasc syst|Surg comp-peri vasc syst
C0729250|T037|HT|997.3|ICD9CM|Respiratory complications, not elsewhere classified|Respiratory complications, not elsewhere classified
C1701940|T047|PT|997.31|ICD9CM|Ventilator associated pneumonia|Ventilator associated pneumonia
C1701940|T047|AB|997.31|ICD9CM|Ventltr assoc pneumonia|Ventltr assoc pneumonia
C3161132|T047|AB|997.32|ICD9CM|Postproc aspiration pneu|Postproc aspiration pneu
C3161132|T047|PT|997.32|ICD9CM|Postprocedural aspiration pneumonia|Postprocedural aspiration pneumonia
C2349769|T047|PT|997.39|ICD9CM|Other respiratory complications|Other respiratory complications
C2349769|T047|AB|997.39|ICD9CM|Respiratory comp NEC|Respiratory comp NEC
C0161819|T046|HT|997.4|ICD9CM|Digestive system complications|Digestive system complications
C3161133|T046|AB|997.41|ICD9CM|Ret cholelh fol cholecys|Ret cholelh fol cholecys
C3161133|T046|PT|997.41|ICD9CM|Retained cholelithiasis following cholecystectomy|Retained cholelithiasis following cholecystectomy
C3161134|T046|AB|997.49|ICD9CM|Oth digestv system comp|Oth digestv system comp
C3161134|T046|PT|997.49|ICD9CM|Other digestive system complications|Other digestive system complications
C0595943|T046|AB|997.5|ICD9CM|Surg compl-urinary tract|Surg compl-urinary tract
C0595943|T046|PT|997.5|ICD9CM|Urinary complications, not elsewhere classified|Urinary complications, not elsewhere classified
C0302473|T046|HT|997.6|ICD9CM|Amputation stump complication|Amputation stump complication
C0161821|T037|AB|997.60|ICD9CM|Amputat stump compl NOS|Amputat stump compl NOS
C0161821|T037|PT|997.60|ICD9CM|Unspecified complication of amputation stump|Unspecified complication of amputation stump
C0392617|T047|AB|997.61|ICD9CM|Neuroma amputation stump|Neuroma amputation stump
C0392617|T047|PT|997.61|ICD9CM|Neuroma of amputation stump|Neuroma of amputation stump
C0161824|T046|PT|997.62|ICD9CM|Infection (chronic) of amputation stump|Infection (chronic) of amputation stump
C0161824|T046|AB|997.62|ICD9CM|Infection amputat stump|Infection amputat stump
C2891341|T046|AB|997.69|ICD9CM|Amputat stump compl NEC|Amputat stump compl NEC
C2891341|T046|PT|997.69|ICD9CM|Other amputation stump complication|Other amputation stump complication
C0949152|T047|HT|997.7|ICD9CM|Vascular complications of other vessels|Vascular complications of other vessels
C0949150|T047|AB|997.71|ICD9CM|Vasc comp mesenteric art|Vasc comp mesenteric art
C0949150|T047|PT|997.71|ICD9CM|Vascular complications of mesenteric artery|Vascular complications of mesenteric artery
C0949151|T047|AB|997.72|ICD9CM|Vasc comp renal artery|Vasc comp renal artery
C0949151|T047|PT|997.72|ICD9CM|Vascular complications of renal artery|Vascular complications of renal artery
C0949152|T047|AB|997.79|ICD9CM|Vascular comp vessel NEC|Vascular comp vessel NEC
C0949152|T047|PT|997.79|ICD9CM|Vascular complications of other vessels|Vascular complications of other vessels
C0302415|T037|HT|997.9|ICD9CM|Complications affecting other specified body systems, not elsewhere classified|Complications affecting other specified body systems, not elsewhere classified
C0020538|T047|PT|997.91|ICD9CM|Complications affecting other specified body systems, not elsewhere classified, hypertension|Complications affecting other specified body systems, not elsewhere classified, hypertension
C0020538|T047|AB|997.91|ICD9CM|Surg comp - hypertension|Surg comp - hypertension
C0375724|T037|PT|997.99|ICD9CM|Complications affecting other specified body systems, not elsewhere classified|Complications affecting other specified body systems, not elsewhere classified
C0375724|T037|AB|997.99|ICD9CM|Surg compl-body syst NEC|Surg compl-body syst NEC
C0869286|T037|HT|998|ICD9CM|Other complications of procedures, NEC|Other complications of procedures, NEC
C0032792|T046|HT|998.0|ICD9CM|Postoperative shock|Postoperative shock
C0032792|T046|AB|998.00|ICD9CM|Postoperative shock, NOS|Postoperative shock, NOS
C0032792|T046|PT|998.00|ICD9CM|Postoperative shock, unspecified|Postoperative shock, unspecified
C3161135|T047|AB|998.01|ICD9CM|Postop shock,cardiogenic|Postop shock,cardiogenic
C3161135|T047|PT|998.01|ICD9CM|Postoperative shock, cardiogenic|Postoperative shock, cardiogenic
C0342957|T047|AB|998.02|ICD9CM|Postop shock, septic|Postop shock, septic
C0342957|T047|PT|998.02|ICD9CM|Postoperative shock, septic|Postoperative shock, septic
C3161136|T046|AB|998.09|ICD9CM|Postop shock, other|Postop shock, other
C3161136|T046|PT|998.09|ICD9CM|Postoperative shock, other|Postoperative shock, other
C0274397|T047|HT|998.1|ICD9CM|Hemorrhage or hematoma complicating a procedure|Hemorrhage or hematoma complicating a procedure
C0375725|T046|AB|998.11|ICD9CM|Hemorrhage complic proc|Hemorrhage complic proc
C0375725|T046|PT|998.11|ICD9CM|Hemorrhage complicating a procedure|Hemorrhage complicating a procedure
C0375726|T046|AB|998.12|ICD9CM|Hematoma complic proc|Hematoma complic proc
C0375726|T046|PT|998.12|ICD9CM|Hematoma complicating a procedure|Hematoma complicating a procedure
C0375727|T046|PT|998.13|ICD9CM|Seroma complicating a procedure|Seroma complicating a procedure
C0375727|T046|AB|998.13|ICD9CM|Seroma complicting proc|Seroma complicting proc
C0161829|T037|AB|998.2|ICD9CM|Accidental op laceration|Accidental op laceration
C0161829|T037|PT|998.2|ICD9CM|Accidental puncture or laceration during a procedure, not elsewhere classified|Accidental puncture or laceration during a procedure, not elsewhere classified
C0259768|T046|HT|998.3|ICD9CM|Disruption of wound|Disruption of wound
C0259768|T046|PT|998.30|ICD9CM|Disruption of wound, unspecified|Disruption of wound, unspecified
C0259768|T046|AB|998.30|ICD9CM|Wound disruption NOS|Wound disruption NOS
C1135269|T047|AB|998.31|ICD9CM|Disrup internal op wound|Disrup internal op wound
C1135269|T047|PT|998.31|ICD9CM|Disruption of internal operation (surgical) wound|Disruption of internal operation (surgical) wound
C1135270|T047|AB|998.32|ICD9CM|Disrup-external op wound|Disrup-external op wound
C1135270|T047|PT|998.32|ICD9CM|Disruption of external operation (surgical) wound|Disruption of external operation (surgical) wound
C2349787|T046|AB|998.33|ICD9CM|Disrpt trauma wound repr|Disrpt trauma wound repr
C2349787|T046|PT|998.33|ICD9CM|Disruption of traumatic injury wound repair|Disruption of traumatic injury wound repair
C0161831|T037|AB|998.4|ICD9CM|FB left during procedure|FB left during procedure
C0161831|T037|PT|998.4|ICD9CM|Foreign body accidentally left during a procedure|Foreign body accidentally left during a procedure
C0392618|T046|HT|998.5|ICD9CM|Postoperative infection|Postoperative infection
C0375728|T047|AB|998.51|ICD9CM|Infected postop seroma|Infected postop seroma
C0375728|T047|PT|998.51|ICD9CM|Infected postoperative seroma|Infected postoperative seroma
C0375729|T047|AB|998.59|ICD9CM|Other postop infection|Other postop infection
C0375729|T047|PT|998.59|ICD9CM|Other postoperative infection|Other postoperative infection
C0161832|T020|AB|998.6|ICD9CM|Persist postop fistula|Persist postop fistula
C0161832|T020|PT|998.6|ICD9CM|Persistent postoperative fistula|Persistent postoperative fistula
C0161833|T047|PT|998.7|ICD9CM|Acute reaction to foreign substance accidentally left during a procedure|Acute reaction to foreign substance accidentally left during a procedure
C0161833|T047|AB|998.7|ICD9CM|Postop forgn subst react|Postop forgn subst react
C0302422|T037|HT|998.8|ICD9CM|Other specified complications of procedures, not elsewhere classified|Other specified complications of procedures, not elsewhere classified
C0274411|T046|PT|998.81|ICD9CM|Emphysema (subcutaneous) (surgical) resulting from procedure|Emphysema (subcutaneous) (surgical) resulting from procedure
C0274411|T046|AB|998.81|ICD9CM|Emphysema rsult frm proc|Emphysema rsult frm proc
C0375731|T020|PT|998.82|ICD9CM|Cataract fragments in eye following cataract surgery|Cataract fragments in eye following cataract surgery
C0375731|T020|AB|998.82|ICD9CM|Ctrct frgmt frm ctr surg|Ctrct frgmt frm ctr surg
C0375732|T046|AB|998.83|ICD9CM|Non-healing surgcl wound|Non-healing surgcl wound
C0375732|T046|PT|998.83|ICD9CM|Non-healing surgical wound|Non-healing surgical wound
C0161834|T046|AB|998.89|ICD9CM|Oth spcf cmplc procd NEC|Oth spcf cmplc procd NEC
C0161834|T046|PT|998.89|ICD9CM|Other specified complications of procedures not elsewhere classified|Other specified complications of procedures not elsewhere classified
C0869442|T046|AB|998.9|ICD9CM|Surgical complicat NOS|Surgical complicat NOS
C0869442|T046|PT|998.9|ICD9CM|Unspecified complication of procedure, not elsewhere classified|Unspecified complication of procedure, not elsewhere classified
C0546949|T037|HT|999|ICD9CM|Complications of medical care, not elsewhere classified|Complications of medical care, not elsewhere classified
C0302424|T047|AB|999.0|ICD9CM|Generalized vaccinia|Generalized vaccinia
C0302424|T047|PT|999.0|ICD9CM|Generalized vaccinia as a complication of medical care, not elsewhere classified|Generalized vaccinia as a complication of medical care, not elsewhere classified
C0302425|T046|AB|999.1|ICD9CM|Air embol comp med care|Air embol comp med care
C0302425|T046|PT|999.1|ICD9CM|Air embolism as a complication of medical care, not elsewhere classified|Air embolism as a complication of medical care, not elsewhere classified
C0302426|T046|PT|999.2|ICD9CM|Other vascular complications of medical care, not elsewhere classified|Other vascular complications of medical care, not elsewhere classified
C0302426|T046|AB|999.2|ICD9CM|Vasc comp med care NEC|Vasc comp med care NEC
C0302427|T037|HT|999.3|ICD9CM|Other infection due to medical care, not elsewhere classified|Other infection due to medical care, not elsewhere classified
C1955545|T046|AB|999.31|ICD9CM|Oth/uns inf-cen ven cath|Oth/uns inf-cen ven cath
C1955545|T046|PT|999.31|ICD9CM|Other and unspecified infection due to central venous catheter|Other and unspecified infection due to central venous catheter
C3161137|T046|AB|999.32|ICD9CM|Blood inf dt cen ven cth|Blood inf dt cen ven cth
C3161137|T046|PT|999.32|ICD9CM|Bloodstream infection due to central venous catheter|Bloodstream infection due to central venous catheter
C3161138|T046|AB|999.33|ICD9CM|Lcl inf dt cen ven cth|Lcl inf dt cen ven cth
C3161138|T046|PT|999.33|ICD9CM|Local infection due to central venous catheter|Local infection due to central venous catheter
C3161139|T046|AB|999.34|ICD9CM|Ac inf fol trans,inf bld|Ac inf fol trans,inf bld
C3161139|T046|PT|999.34|ICD9CM|Acute infection following transfusion, infusion, or injection of blood and blood products|Acute infection following transfusion, infusion, or injection of blood and blood products
C1955550|T047|AB|999.39|ICD9CM|Infect fol infus/inj/vac|Infect fol infus/inj/vac
C1955550|T047|PT|999.39|ICD9CM|Infection following other infusion, injection, transfusion, or vaccination|Infection following other infusion, injection, transfusion, or vaccination
C3161458|T046|HT|999.4|ICD9CM|Anaphylactic reaction due to serum, not elsewhere classified|Anaphylactic reaction due to serum, not elsewhere classified
C3161140|T046|AB|999.41|ICD9CM|Anaphyl d/t adm bld/prod|Anaphyl d/t adm bld/prod
C3161140|T046|PT|999.41|ICD9CM|Anaphylactic reaction due to administration of blood and blood products|Anaphylactic reaction due to administration of blood and blood products
C3161141|T046|AB|999.42|ICD9CM|Anaphyl react d/t vaccin|Anaphyl react d/t vaccin
C3161141|T046|PT|999.42|ICD9CM|Anaphylactic reaction due to vaccination|Anaphylactic reaction due to vaccination
C3161142|T046|AB|999.49|ICD9CM|Anaph react d/t ot serum|Anaph react d/t ot serum
C3161142|T046|PT|999.49|ICD9CM|Anaphylactic reaction due to other serum|Anaphylactic reaction due to other serum
C0302428|T046|HT|999.5|ICD9CM|Other serum reaction, not elsewhere classified|Other serum reaction, not elsewhere classified
C3161143|T046|AB|999.51|ICD9CM|Ot serum react d/t blood|Ot serum react d/t blood
C3161143|T046|PT|999.51|ICD9CM|Other serum reaction due to administration of blood and blood products|Other serum reaction due to administration of blood and blood products
C3161144|T046|AB|999.52|ICD9CM|Ot serum react d/t vacc|Ot serum react d/t vacc
C3161144|T046|PT|999.52|ICD9CM|Other serum reaction due to vaccination|Other serum reaction due to vaccination
C0478483|T046|AB|999.59|ICD9CM|Other serum reaction|Other serum reaction
C0478483|T046|PT|999.59|ICD9CM|Other serum reaction|Other serum reaction
C2886803|T046|HT|999.6|ICD9CM|ABO incompatibility reaction due to transfusion of blood or blood products|ABO incompatibility reaction due to transfusion of blood or blood products
C2921199|T046|AB|999.60|ICD9CM|Abo incompat react NOS|Abo incompat react NOS
C2921199|T046|PT|999.60|ICD9CM|ABO incompatibility reaction, unspecified|ABO incompatibility reaction, unspecified
C2921202|T046|AB|999.61|ICD9CM|Abo incomp/HTR NEC|Abo incomp/HTR NEC
C2921202|T046|PT|999.61|ICD9CM|ABO incompatibility with hemolytic transfusion reaction not specified as acute or delayed|ABO incompatibility with hemolytic transfusion reaction not specified as acute or delayed
C2921204|T046|AB|999.62|ICD9CM|Abo incompat/acute HTR|Abo incompat/acute HTR
C2921204|T046|PT|999.62|ICD9CM|ABO incompatibility with acute hemolytic transfusion reaction|ABO incompatibility with acute hemolytic transfusion reaction
C2921207|T046|AB|999.63|ICD9CM|Abo incompat/delay HTR|Abo incompat/delay HTR
C2921207|T046|PT|999.63|ICD9CM|ABO incompatibility with delayed hemolytic transfusion reaction|ABO incompatibility with delayed hemolytic transfusion reaction
C2921211|T046|AB|999.69|ICD9CM|Abo incompat reactn NEC|Abo incompat reactn NEC
C2921211|T046|PT|999.69|ICD9CM|Other ABO incompatibility reaction|Other ABO incompatibility reaction
C2921214|T046|HT|999.7|ICD9CM|Rh and other non-ABO incompatibility reaction due to transfusion of blood or blood products|Rh and other non-ABO incompatibility reaction due to transfusion of blood or blood products
C2921216|T046|AB|999.70|ICD9CM|Rh incompat reaction NOS|Rh incompat reaction NOS
C2921216|T046|PT|999.70|ICD9CM|Rh incompatibility reaction, unspecified|Rh incompatibility reaction, unspecified
C2921222|T046|AB|999.71|ICD9CM|Rh incomp/HTR NEC|Rh incomp/HTR NEC
C2921222|T046|PT|999.71|ICD9CM|Rh incompatibility with hemolytic transfusion reaction not specified as acute or delayed|Rh incompatibility with hemolytic transfusion reaction not specified as acute or delayed
C2921225|T046|AB|999.72|ICD9CM|Rh incompat/acute HTR|Rh incompat/acute HTR
C2921225|T046|PT|999.72|ICD9CM|Rh incompatibility with acute hemolytic transfusion reaction|Rh incompatibility with acute hemolytic transfusion reaction
C2921229|T046|AB|999.73|ICD9CM|Rh incompat/delay HTR|Rh incompat/delay HTR
C2921229|T046|PT|999.73|ICD9CM|Rh incompatibility with delayed hemolytic transfusion reaction|Rh incompatibility with delayed hemolytic transfusion reaction
C2921232|T047|PT|999.74|ICD9CM|Other Rh incompatibility reaction|Other Rh incompatibility reaction
C2921232|T047|AB|999.74|ICD9CM|Rh incompat reaction NEC|Rh incompat reaction NEC
C2921235|T047|AB|999.75|ICD9CM|Non-abo incomp react NOS|Non-abo incomp react NOS
C2921235|T047|PT|999.75|ICD9CM|Non-ABO incompatibility reaction, unspecified|Non-ABO incompatibility reaction, unspecified
C2921242|T047|AB|999.76|ICD9CM|Non-abo incomp/HTR NEC|Non-abo incomp/HTR NEC
C2921242|T047|PT|999.76|ICD9CM|Non-ABO incompatibility with hemolytic transfusion reaction not specified as acute or delayed|Non-ABO incompatibility with hemolytic transfusion reaction not specified as acute or delayed
C2921245|T046|AB|999.77|ICD9CM|Non-abo incomp/acute HTR|Non-abo incomp/acute HTR
C2921245|T046|PT|999.77|ICD9CM|Non-ABO incompatibility with acute hemolytic transfusion reaction|Non-ABO incompatibility with acute hemolytic transfusion reaction
C2921249|T046|AB|999.78|ICD9CM|Non-abo incomp/delay HTR|Non-abo incomp/delay HTR
C2921249|T046|PT|999.78|ICD9CM|Non-ABO incompatibility with delayed hemolytic transfusion reaction|Non-ABO incompatibility with delayed hemolytic transfusion reaction
C2921252|T047|AB|999.79|ICD9CM|Non-abo incomp react NEC|Non-abo incomp react NEC
C2921252|T047|PT|999.79|ICD9CM|Other non-ABO incompatibility reaction|Other non-ABO incompatibility reaction
C2349800|T037|HT|999.8|ICD9CM|Other infusion and transfusion reaction, not elsewhere classified|Other infusion and transfusion reaction, not elsewhere classified
C0274435|T046|AB|999.80|ICD9CM|Transfusion reaction NOS|Transfusion reaction NOS
C0274435|T046|PT|999.80|ICD9CM|Transfusion reaction, unspecified|Transfusion reaction, unspecified
C2349794|T037|PT|999.81|ICD9CM|Extravasation of vesicant chemotherapy|Extravasation of vesicant chemotherapy
C2349794|T037|AB|999.81|ICD9CM|Extravstn vesicant chemo|Extravstn vesicant chemo
C2349796|T037|PT|999.82|ICD9CM|Extravasation of other vesicant agent|Extravasation of other vesicant agent
C2349796|T037|AB|999.82|ICD9CM|Extravasn vesicant NEC|Extravasn vesicant NEC
C2921258|T046|AB|999.83|ICD9CM|Hemolytc trans react NOS|Hemolytc trans react NOS
C2921258|T046|PT|999.83|ICD9CM|Hemolytic transfusion reaction, incompatibility unspecified|Hemolytic transfusion reaction, incompatibility unspecified
C2921260|T046|PT|999.84|ICD9CM|Acute hemolytic transfusion reaction, incompatibility unspecified|Acute hemolytic transfusion reaction, incompatibility unspecified
C2921260|T046|AB|999.84|ICD9CM|Acute HTR NOS|Acute HTR NOS
C2921262|T046|PT|999.85|ICD9CM|Delayed hemolytic transfusion reaction, incompatibility unspecified|Delayed hemolytic transfusion reaction, incompatibility unspecified
C2921262|T046|AB|999.85|ICD9CM|Delayed HTR NOS|Delayed HTR NOS
C2349798|T047|AB|999.88|ICD9CM|Infusion reaction NEC|Infusion reaction NEC
C2349798|T047|PT|999.88|ICD9CM|Other infusion reaction|Other infusion reaction
C2349799|T046|PT|999.89|ICD9CM|Other transfusion reaction|Other transfusion reaction
C2349799|T046|AB|999.89|ICD9CM|Transfusion reaction NEC|Transfusion reaction NEC
C0302430|T037|AB|999.9|ICD9CM|Complic med care NEC/NOS|Complic med care NEC/NOS
C0302430|T037|PT|999.9|ICD9CM|Other and unspecified complications of medical care, not elsewhere classified|Other and unspecified complications of medical care, not elsewhere classified
C2712898|T033|HT|E000|ICD9CM|External cause status|External cause status
C2712898|T033|HT|E000-E000.9|ICD9CM|EXTERNAL CAUSE STATUS|EXTERNAL CAUSE STATUS
C2712384|T037|PT|E000.0|ICD9CM|Civilian activity done for income or pay|Civilian activity done for income or pay
C2712384|T037|AB|E000.0|ICD9CM|Civilian activity-income|Civilian activity-income
C2712385|T037|PT|E000.1|ICD9CM|Military activity|Military activity
C2712385|T037|AB|E000.1|ICD9CM|Military activity|Military activity
C2712386|T033|AB|E000.8|ICD9CM|Externl cause status NEC|Externl cause status NEC
C2712386|T033|PT|E000.8|ICD9CM|Other external cause status|Other external cause status
C2712387|T037|AB|E000.9|ICD9CM|Externl cause status NOS|Externl cause status NOS
C2712387|T037|PT|E000.9|ICD9CM|Unspecified external cause status|Unspecified external cause status
C0260969|T037|HT|E800|ICD9CM|Railway accident involving collision with rolling stock|Railway accident involving collision with rolling stock
C0414085|T037|HT|E800-E807.9|ICD9CM|RAILWAY ACCIDENTS|RAILWAY ACCIDENTS
C0362049|T037|HT|E800-E848.9|ICD9CM|TRANSPORT ACCIDENTS|TRANSPORT ACCIDENTS
C0260970|T037|PT|E800.0|ICD9CM|Railway accident involving collision with rolling stock and injuring railway employee|Railway accident involving collision with rolling stock and injuring railway employee
C0260970|T037|AB|E800.0|ICD9CM|RR collision NOS-employ|RR collision NOS-employ
C0260971|T037|PT|E800.1|ICD9CM|Railway accident involving collision with rolling stock and injuring passenger on railway|Railway accident involving collision with rolling stock and injuring passenger on railway
C0260971|T037|AB|E800.1|ICD9CM|RR coll NOS-passenger|RR coll NOS-passenger
C0260972|T037|PT|E800.2|ICD9CM|Railway accident involving collision with rolling stock and injuring pedestrian|Railway accident involving collision with rolling stock and injuring pedestrian
C0260972|T037|AB|E800.2|ICD9CM|RR coll NOS-pedestrian|RR coll NOS-pedestrian
C0260973|T037|PT|E800.3|ICD9CM|Railway accident involving collision with rolling stock and injuring pedal cyclist|Railway accident involving collision with rolling stock and injuring pedal cyclist
C0260973|T037|AB|E800.3|ICD9CM|RR coll NOS-ped cyclist|RR coll NOS-ped cyclist
C0260974|T037|PT|E800.8|ICD9CM|Railway accident involving collision with rolling stock and injuring other specified person|Railway accident involving collision with rolling stock and injuring other specified person
C0260974|T037|AB|E800.8|ICD9CM|RR coll NOS-person NEC|RR coll NOS-person NEC
C0260975|T037|PT|E800.9|ICD9CM|Railway accident involving collision with rolling stock and injuring unspecified person|Railway accident involving collision with rolling stock and injuring unspecified person
C0260975|T037|AB|E800.9|ICD9CM|RR coll NOS-person NOS|RR coll NOS-person NOS
C0260976|T037|HT|E801|ICD9CM|Railway accident involving collision with other object|Railway accident involving collision with other object
C0414276|T037|HT|E804|ICD9CM|Fall in, on, or from railway train|Fall in, on, or from railway train
C0414302|T037|HT|E805|ICD9CM|Hit by rolling stock|Hit by rolling stock
C0261012|T037|PT|E806.0|ICD9CM|Other specified railway accident injuring railway employee|Other specified railway accident injuring railway employee
C0261012|T037|AB|E806.0|ICD9CM|RR acc NEC-employee|RR acc NEC-employee
C0261016|T037|PT|E806.8|ICD9CM|Other specified railway accident injuring other specified person|Other specified railway accident injuring other specified person
C0261016|T037|AB|E806.8|ICD9CM|RR acc NEC-person NEC|RR acc NEC-person NEC
C0261017|T037|PT|E806.9|ICD9CM|Other specified railway accident injuring unspecified person|Other specified railway accident injuring unspecified person
C0261017|T037|AB|E806.9|ICD9CM|RR acc NEC-person NOS|RR acc NEC-person NOS
C0414085|T037|HT|E807|ICD9CM|Railway accident of unspecified nature|Railway accident of unspecified nature
C0414438|T037|HT|E810|ICD9CM|Motor vehicle traffic accident involving collision with train|Motor vehicle traffic accident involving collision with train
C4760746|T037|HT|E810-E819.9|ICD9CM|MOTOR VEHICLE TRAFFIC ACCIDENTS|MOTOR VEHICLE TRAFFIC ACCIDENTS
C0261028|T037|PT|E810.2|ICD9CM|Motor vehicle traffic accident involving collision with train injuring motorcyclist|Motor vehicle traffic accident involving collision with train injuring motorcyclist
C0261028|T037|AB|E810.2|ICD9CM|Mv-train coll-motorcycl|Mv-train coll-motorcycl
C0261029|T037|PT|E810.3|ICD9CM|Motor vehicle traffic accident involving collision with train injuring passenger on motorcycle|Motor vehicle traffic accident involving collision with train injuring passenger on motorcycle
C0261029|T037|AB|E810.3|ICD9CM|Mv-train coll-mcycl psgr|Mv-train coll-mcycl psgr
C0261030|T037|PT|E810.4|ICD9CM|Motor vehicle traffic accident involving collision with train injuring occupant of streetcar|Motor vehicle traffic accident involving collision with train injuring occupant of streetcar
C0261030|T037|AB|E810.4|ICD9CM|Mv-train coll-st car|Mv-train coll-st car
C0414441|T037|PT|E810.6|ICD9CM|Motor vehicle traffic accident involving collision with train injuring pedal cyclist|Motor vehicle traffic accident involving collision with train injuring pedal cyclist
C0414441|T037|AB|E810.6|ICD9CM|Mv-train coll-ped cycl|Mv-train coll-ped cycl
C0414440|T037|PT|E810.7|ICD9CM|Motor vehicle traffic accident involving collision with train injuring pedestrian|Motor vehicle traffic accident involving collision with train injuring pedestrian
C0414440|T037|AB|E810.7|ICD9CM|Mv-train coll-pedest|Mv-train coll-pedest
C0414439|T037|PT|E810.8|ICD9CM|Motor vehicle traffic accident involving collision with train injuring other specified person|Motor vehicle traffic accident involving collision with train injuring other specified person
C0414439|T037|AB|E810.8|ICD9CM|Mv-train coll-pers NEC|Mv-train coll-pers NEC
C0414438|T037|PT|E810.9|ICD9CM|Motor vehicle traffic accident involving collision with train injuring unspecified person|Motor vehicle traffic accident involving collision with train injuring unspecified person
C0414438|T037|AB|E810.9|ICD9CM|Mv-train coll-pers NOS|Mv-train coll-pers NOS
C0261036|T037|HT|E811|ICD9CM|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle
C0261039|T037|AB|E811.2|ICD9CM|Reentrant coll-motcycl|Reentrant coll-motcycl
C0261040|T037|AB|E811.3|ICD9CM|Reentrant coll-mcyc psgr|Reentrant coll-mcyc psgr
C0261041|T037|AB|E811.4|ICD9CM|Reentrant coll-st car|Reentrant coll-st car
C0261043|T037|AB|E811.6|ICD9CM|Reentrant coll-ped cycl|Reentrant coll-ped cycl
C0261045|T037|AB|E811.8|ICD9CM|Reentrant coll-pers NEC|Reentrant coll-pers NEC
C0261046|T037|AB|E811.9|ICD9CM|Reentrant coll-pers NOS|Reentrant coll-pers NOS
C0261061|T037|PT|E813.2|ICD9CM|Motor vehicle traffic accident involving collision with other vehicle injuring motorcyclist|Motor vehicle traffic accident involving collision with other vehicle injuring motorcyclist
C0261061|T037|AB|E813.2|ICD9CM|Mv-oth veh coll-motcycl|Mv-oth veh coll-motcycl
C0261062|T037|AB|E813.3|ICD9CM|Mv-oth veh coll-mcyc psg|Mv-oth veh coll-mcyc psg
C0261063|T037|PT|E813.4|ICD9CM|Motor vehicle traffic accident involving collision with other vehicle injuring occupant of streetcar|Motor vehicle traffic accident involving collision with other vehicle injuring occupant of streetcar
C0261063|T037|AB|E813.4|ICD9CM|Mv-oth veh coll-st car|Mv-oth veh coll-st car
C0414471|T037|PT|E813.9|ICD9CM|Motor vehicle traffic accident involving collision with other vehicle injuring unspecified person|Motor vehicle traffic accident involving collision with other vehicle injuring unspecified person
C0414471|T037|AB|E813.9|ICD9CM|Mv-oth veh coll-pers NOS|Mv-oth veh coll-pers NOS
C0261069|T037|HT|E814|ICD9CM|Motor vehicle traffic accident involving collision with pedestrian|Motor vehicle traffic accident involving collision with pedestrian
C0261080|T037|HT|E815|ICD9CM|Other motor vehicle traffic accident involving collision on the highway|Other motor vehicle traffic accident involving collision on the highway
C0261091|T037|HT|E816|ICD9CM|Motor vehicle traffic accident due to loss of control, without collision on the highway|Motor vehicle traffic accident due to loss of control, without collision on the highway
C0414740|T037|AB|E816.2|ICD9CM|Loss control mv-mocycl|Loss control mv-mocycl
C0261095|T037|AB|E816.3|ICD9CM|Loss control mv-mcyc psg|Loss control mv-mcyc psg
C0261096|T037|AB|E816.4|ICD9CM|Loss cont mv acc-st car|Loss cont mv acc-st car
C0414736|T037|AB|E816.6|ICD9CM|Loss control mv-ped cycl|Loss control mv-ped cycl
C0414735|T037|AB|E816.7|ICD9CM|Loss control mv-pedest|Loss control mv-pedest
C0414734|T037|AB|E816.8|ICD9CM|Loss control mv-pers NEC|Loss control mv-pers NEC
C0414733|T037|AB|E816.9|ICD9CM|Loss control mv-pers NOS|Loss control mv-pers NOS
C0261102|T037|HT|E817|ICD9CM|Noncollision motor vehicle traffic accident while boarding or alighting|Noncollision motor vehicle traffic accident while boarding or alighting
C0026614|T037|HT|E819|ICD9CM|Motor vehicle traffic accident of unspecified nature|Motor vehicle traffic accident of unspecified nature
C0415270|T037|HT|E820|ICD9CM|Nontraffic accident involving motor-driven snow vehicle|Nontraffic accident involving motor-driven snow vehicle
C0178348|T037|HT|E820-E825.9|ICD9CM|MOTOR VEHICLE NONTRAFFIC ACCIDENTS|MOTOR VEHICLE NONTRAFFIC ACCIDENTS
C0261141|T037|PT|E820.6|ICD9CM|Nontraffic accident involving motor-driven snow vehicle injuring pedal cyclist|Nontraffic accident involving motor-driven snow vehicle injuring pedal cyclist
C0261141|T037|AB|E820.6|ICD9CM|Snow veh acc-ped cycl|Snow veh acc-ped cycl
C0261142|T037|PT|E820.7|ICD9CM|Nontraffic accident involving motor-driven snow vehicle injuring pedestrian|Nontraffic accident involving motor-driven snow vehicle injuring pedestrian
C0261142|T037|AB|E820.7|ICD9CM|Snow veh acc-pedest|Snow veh acc-pedest
C0261143|T037|PT|E820.8|ICD9CM|Nontraffic accident involving motor-driven snow vehicle injuring other specified person|Nontraffic accident involving motor-driven snow vehicle injuring other specified person
C0261143|T037|AB|E820.8|ICD9CM|Snow veh acc-pers NEC|Snow veh acc-pers NEC
C0261144|T037|PT|E820.9|ICD9CM|Nontraffic accident involving motor-driven snow vehicle injuring unspecified person|Nontraffic accident involving motor-driven snow vehicle injuring unspecified person
C0261144|T037|AB|E820.9|ICD9CM|Snow veh acc-pers NOS|Snow veh acc-pers NOS
C0261156|T037|HT|E822|ICD9CM|Other motor vehicle nontraffic accident involving collision with moving object|Other motor vehicle nontraffic accident involving collision with moving object
C0261167|T037|HT|E823|ICD9CM|Other motor vehicle nontraffic accident involving collision with stationary object|Other motor vehicle nontraffic accident involving collision with stationary object
C0261178|T037|HT|E824|ICD9CM|Other motor vehicle nontraffic accident while boarding and alighting|Other motor vehicle nontraffic accident while boarding and alighting
C0261189|T037|HT|E825|ICD9CM|Other motor vehicle nontraffic accident of other and unspecified nature|Other motor vehicle nontraffic accident of other and unspecified nature
C0261200|T037|HT|E826|ICD9CM|Pedal cycle accident|Pedal cycle accident
C0176004|T037|HT|E826-E829.9|ICD9CM|OTHER ROAD VEHICLE ACCIDENTS|OTHER ROAD VEHICLE ACCIDENTS
C0261201|T037|AB|E826.0|ICD9CM|Pedal cycle acc-pedest|Pedal cycle acc-pedest
C0261201|T037|PT|E826.0|ICD9CM|Pedal cycle accident injuring pedestrian|Pedal cycle accident injuring pedestrian
C0261202|T037|AB|E826.1|ICD9CM|Ped cycl acc-ped cyclist|Ped cycl acc-ped cyclist
C0261202|T037|PT|E826.1|ICD9CM|Pedal cycle accident injuring pedal cyclist|Pedal cycle accident injuring pedal cyclist
C0261203|T037|AB|E826.2|ICD9CM|Ped cycle acc-anim rider|Ped cycle acc-anim rider
C0261203|T037|PT|E826.2|ICD9CM|Pedal cycle accident injuring rider of animal|Pedal cycle accident injuring rider of animal
C0415505|T037|AB|E826.3|ICD9CM|Ped cyc acc-occ anim veh|Ped cyc acc-occ anim veh
C0415505|T037|PT|E826.3|ICD9CM|Pedal cycle accident injuring occupant of animal-drawn vehicle|Pedal cycle accident injuring occupant of animal-drawn vehicle
C0261205|T037|AB|E826.4|ICD9CM|Ped cycle acc-occ st car|Ped cycle acc-occ st car
C0261205|T037|PT|E826.4|ICD9CM|Pedal cycle accident injuring occupant of streetcar|Pedal cycle accident injuring occupant of streetcar
C0261206|T037|AB|E826.8|ICD9CM|Ped cycle acc-pers NEC|Ped cycle acc-pers NEC
C0261206|T037|PT|E826.8|ICD9CM|Pedal cycle accident injuring other specified person|Pedal cycle accident injuring other specified person
C0261207|T037|AB|E826.9|ICD9CM|Ped cycle acc-pers NOS|Ped cycle acc-pers NOS
C0261207|T037|PT|E826.9|ICD9CM|Pedal cycle accident injuring unspecified person|Pedal cycle accident injuring unspecified person
C0261208|T037|HT|E827|ICD9CM|Animal-drawn vehicle accident|Animal-drawn vehicle accident
C0261209|T037|AB|E827.0|ICD9CM|Animal drawn veh-pedest|Animal drawn veh-pedest
C0261209|T037|PT|E827.0|ICD9CM|Animal-drawn vehicle accident injuring pedestrian|Animal-drawn vehicle accident injuring pedestrian
C0261210|T037|AB|E827.2|ICD9CM|Anim drawn veh-anim rid|Anim drawn veh-anim rid
C0261210|T037|PT|E827.2|ICD9CM|Animal-drawn vehicle accident injuring rider of animal|Animal-drawn vehicle accident injuring rider of animal
C0261211|T037|AB|E827.3|ICD9CM|Animal drawn veh-occupan|Animal drawn veh-occupan
C0261211|T037|PT|E827.3|ICD9CM|Animal-drawn vehicle accident injuring occupant of animal drawn vehicle|Animal-drawn vehicle accident injuring occupant of animal drawn vehicle
C0261212|T037|AB|E827.4|ICD9CM|Anim drawn-occ st car|Anim drawn-occ st car
C0261212|T037|PT|E827.4|ICD9CM|Animal-drawn vehicle accident injuring occupant of streetcar|Animal-drawn vehicle accident injuring occupant of streetcar
C0261213|T037|AB|E827.8|ICD9CM|Anim drawn veh-pers NEC|Anim drawn veh-pers NEC
C0261213|T037|PT|E827.8|ICD9CM|Animal-drawn vehicle accident injuring other specified person|Animal-drawn vehicle accident injuring other specified person
C0261214|T037|AB|E827.9|ICD9CM|Anim drawn veh-pers NOS|Anim drawn veh-pers NOS
C0261214|T037|PT|E827.9|ICD9CM|Animal-drawn vehicle accident injuring unspecified person|Animal-drawn vehicle accident injuring unspecified person
C0261215|T037|HT|E828|ICD9CM|Accident involving animal being ridden|Accident involving animal being ridden
C0415659|T037|PT|E828.0|ICD9CM|Accident involving animal being ridden injuring pedestrian|Accident involving animal being ridden injuring pedestrian
C0415659|T037|AB|E828.0|ICD9CM|Ridden animal acc-pedest|Ridden animal acc-pedest
C0415658|T037|PT|E828.2|ICD9CM|Accident involving animal being ridden injuring rider of animal|Accident involving animal being ridden injuring rider of animal
C0415658|T037|AB|E828.2|ICD9CM|Ridden animal acc-rider|Ridden animal acc-rider
C0261218|T037|PT|E828.4|ICD9CM|Accident involving animal being ridden injuring occupant of streetcar|Accident involving animal being ridden injuring occupant of streetcar
C0261218|T037|AB|E828.4|ICD9CM|Ridden animal acc-st car|Ridden animal acc-st car
C0176004|T037|HT|E829|ICD9CM|Other road vehicle accidents|Other road vehicle accidents
C0261221|T037|AB|E829.0|ICD9CM|Oth road veh acc-pedest|Oth road veh acc-pedest
C0261221|T037|PT|E829.0|ICD9CM|Other road vehicle accidents injuring pedestrian|Other road vehicle accidents injuring pedestrian
C0414364|T037|AB|E829.8|ICD9CM|Oth rd veh acc-pers NEC|Oth rd veh acc-pers NEC
C0414364|T037|PT|E829.8|ICD9CM|Other road vehicle accidents injuring other specified person|Other road vehicle accidents injuring other specified person
C0261225|T037|HT|E830|ICD9CM|Accident to watercraft causing submersion|Accident to watercraft causing submersion
C2712469|T037|PT|E830.7|ICD9CM|Accident to watercraft causing submersion, occupant of military watercraft, any type|Accident to watercraft causing submersion, occupant of military watercraft, any type
C2712469|T037|AB|E830.7|ICD9CM|Boat submers-military|Boat submers-military
C0261235|T037|HT|E831|ICD9CM|Accident to watercraft causing other injury|Accident to watercraft causing other injury
C2712470|T037|PT|E831.7|ICD9CM|Accident to watercraft causing other injury, occupant of military watercraft, any type|Accident to watercraft causing other injury, occupant of military watercraft, any type
C2712470|T037|AB|E831.7|ICD9CM|Boat acc inj NEC-militry|Boat acc inj NEC-militry
C0261245|T037|HT|E832|ICD9CM|Other accidental submersion or drowning in water transport accident|Other accidental submersion or drowning in water transport accident
C2712471|T037|AB|E832.7|ICD9CM|Submersion NEC-military|Submersion NEC-military
C0261255|T037|HT|E833|ICD9CM|Fall on stairs or ladders in water transport|Fall on stairs or ladders in water transport
C0261256|T037|PT|E833.0|ICD9CM|Fall on stairs or ladders in water transport injuring occupant of small boat, unpowered|Fall on stairs or ladders in water transport injuring occupant of small boat, unpowered
C0261256|T037|AB|E833.0|ICD9CM|W/craft stair fall-unpow|W/craft stair fall-unpow
C0261257|T037|PT|E833.1|ICD9CM|Fall on stairs or ladders in water transport injuring occupant of small boat, powered|Fall on stairs or ladders in water transport injuring occupant of small boat, powered
C0261257|T037|AB|E833.1|ICD9CM|W/craft stair fall-power|W/craft stair fall-power
C0261258|T037|PT|E833.2|ICD9CM|Fall on stairs or ladders in water transport injuring occupant of other watercraft -- crew|Fall on stairs or ladders in water transport injuring occupant of other watercraft -- crew
C0261258|T037|AB|E833.2|ICD9CM|Wtrcraft stair fall-crew|Wtrcraft stair fall-crew
C0261259|T037|AB|E833.3|ICD9CM|Wtrcraft stair fall-psgr|Wtrcraft stair fall-psgr
C0261260|T037|PT|E833.4|ICD9CM|Fall on stairs or ladders in water transport injuring water skier|Fall on stairs or ladders in water transport injuring water skier
C0261260|T037|AB|E833.4|ICD9CM|W/craft stair fall-skier|W/craft stair fall-skier
C0261261|T037|PT|E833.5|ICD9CM|Fall on stairs or ladders in water transport injuring swimmer|Fall on stairs or ladders in water transport injuring swimmer
C0261261|T037|AB|E833.5|ICD9CM|W/craft stair fall-swim|W/craft stair fall-swim
C0261262|T037|PT|E833.6|ICD9CM|Fall on stairs or ladders in water transport injuring dockers, stevedores|Fall on stairs or ladders in water transport injuring dockers, stevedores
C0261262|T037|AB|E833.6|ICD9CM|W/crf stair fall-docker|W/crf stair fall-docker
C2712472|T037|PT|E833.7|ICD9CM|Fall on stairs or ladders in water transport, occupant of military watercraft, any type|Fall on stairs or ladders in water transport, occupant of military watercraft, any type
C2712472|T037|AB|E833.7|ICD9CM|W/crf stair fall-militry|W/crf stair fall-militry
C0261263|T037|PT|E833.8|ICD9CM|Fall on stairs or ladders in water transport injuring other specified person|Fall on stairs or ladders in water transport injuring other specified person
C0261263|T037|AB|E833.8|ICD9CM|W/crf stair fall-per NEC|W/crf stair fall-per NEC
C0261264|T037|PT|E833.9|ICD9CM|Fall on stairs or ladders in water transport injuring unspecified person|Fall on stairs or ladders in water transport injuring unspecified person
C0261264|T037|AB|E833.9|ICD9CM|W/crf stair fall-per NOS|W/crf stair fall-per NOS
C2712473|T037|PT|E834.7|ICD9CM|Other fall from one level to another in water transport, occupant of military watercraft, any type|Other fall from one level to another in water transport, occupant of military watercraft, any type
C2712473|T037|AB|E834.7|ICD9CM|W/crft fall NEC-military|W/crft fall NEC-military
C0261273|T037|PT|E834.8|ICD9CM|Other fall from one level to another in water transport injuring other specified person|Other fall from one level to another in water transport injuring other specified person
C0261273|T037|AB|E834.8|ICD9CM|W/crft fall NEC-pers NEC|W/crft fall NEC-pers NEC
C2712474|T037|PT|E835.7|ICD9CM|Other and unspecified fall in water transport, occupant of military watercraft, any type|Other and unspecified fall in water transport, occupant of military watercraft, any type
C2712474|T037|AB|E835.7|ICD9CM|W/crft fall NEC/NOS-mil|W/crft fall NEC/NOS-mil
C0261285|T037|HT|E836|ICD9CM|Machinery accident in water transport|Machinery accident in water transport
C0261286|T037|AB|E836.0|ICD9CM|Machine acc-unpow boat|Machine acc-unpow boat
C0261286|T037|PT|E836.0|ICD9CM|Machinery accident in water transport injuring occupant of small boat, unpowered|Machinery accident in water transport injuring occupant of small boat, unpowered
C0261287|T037|AB|E836.1|ICD9CM|Mach acc-occ power boat|Mach acc-occ power boat
C0261287|T037|PT|E836.1|ICD9CM|Machinery accident in water transport injuring occupant of small boat, powered|Machinery accident in water transport injuring occupant of small boat, powered
C0261288|T037|PT|E836.2|ICD9CM|Machinery accident in water transport injuring occupant of other watercraft -- crew|Machinery accident in water transport injuring occupant of other watercraft -- crew
C0261288|T037|AB|E836.2|ICD9CM|Machinery accident-crew|Machinery accident-crew
C0261289|T037|AB|E836.3|ICD9CM|Machinery acc-pasngr|Machinery acc-pasngr
C0261289|T037|PT|E836.3|ICD9CM|Machinery accident in water transport injuring occupant of other watercraft -- other than crew|Machinery accident in water transport injuring occupant of other watercraft -- other than crew
C0261290|T037|AB|E836.4|ICD9CM|Machine accident-skier|Machine accident-skier
C0261290|T037|PT|E836.4|ICD9CM|Machinery accident in water transport injuring water skier|Machinery accident in water transport injuring water skier
C0261291|T037|AB|E836.5|ICD9CM|Machine accident-swim|Machine accident-swim
C0261291|T037|PT|E836.5|ICD9CM|Machinery accident in water transport injuring swimmer|Machinery accident in water transport injuring swimmer
C0261292|T037|AB|E836.6|ICD9CM|Machinery acc-docker|Machinery acc-docker
C0261292|T037|PT|E836.6|ICD9CM|Machinery accident in water transport injuring dockers, stevedores|Machinery accident in water transport injuring dockers, stevedores
C2712475|T037|PT|E836.7|ICD9CM|Machinery accident in water transport, occupant of military watercraft, any type|Machinery accident in water transport, occupant of military watercraft, any type
C2712475|T037|AB|E836.7|ICD9CM|W/crft machine-military|W/crft machine-military
C0261293|T037|AB|E836.8|ICD9CM|Machinery acc-pers NEC|Machinery acc-pers NEC
C0261293|T037|PT|E836.8|ICD9CM|Machinery accident in water transport injuring other specified person|Machinery accident in water transport injuring other specified person
C0261294|T037|AB|E836.9|ICD9CM|Machinery acc-pers NOS|Machinery acc-pers NOS
C0261294|T037|PT|E836.9|ICD9CM|Machinery accident in water transport injuring unspecified person|Machinery accident in water transport injuring unspecified person
C0261295|T037|HT|E837|ICD9CM|Explosion, fire, or burning in watercraft|Explosion, fire, or burning in watercraft
C2712476|T037|PT|E837.7|ICD9CM|Explosion, fire, or burning in watercraft, occupant of military watercraft, any type|Explosion, fire, or burning in watercraft, occupant of military watercraft, any type
C2712476|T037|AB|E837.7|ICD9CM|W/crft explosn-military|W/crft explosn-military
C0261314|T037|HT|E838|ICD9CM|Other and unspecified water transport accident|Other and unspecified water transport accident
C0261306|T037|PT|E838.0|ICD9CM|Other and unspecified water transport accident injuring occupant of small boat, unpowered|Other and unspecified water transport accident injuring occupant of small boat, unpowered
C0261306|T037|AB|E838.0|ICD9CM|Watercraft acc NEC-unpow|Watercraft acc NEC-unpow
C0261307|T037|PT|E838.1|ICD9CM|Other and unspecified water transport accident injuring occupant of small boat, powered|Other and unspecified water transport accident injuring occupant of small boat, powered
C0261307|T037|AB|E838.1|ICD9CM|Watercraft acc NEC-power|Watercraft acc NEC-power
C0261308|T037|PT|E838.2|ICD9CM|Other and unspecified water transport accident injuring occupant of other watercraft -- crew|Other and unspecified water transport accident injuring occupant of other watercraft -- crew
C0261308|T037|AB|E838.2|ICD9CM|Watercraft acc NEC-crew|Watercraft acc NEC-crew
C0261309|T037|AB|E838.3|ICD9CM|Watercrft acc NEC-pasngr|Watercrft acc NEC-pasngr
C2712477|T037|PT|E838.7|ICD9CM|Other and unspecified water transport accident, occupant of military watercraft, any type|Other and unspecified water transport accident, occupant of military watercraft, any type
C2712477|T037|AB|E838.7|ICD9CM|W/crft-military NEC/NOS|W/crft-military NEC/NOS
C0261313|T037|PT|E838.8|ICD9CM|Other and unspecified water transport accident injuring other specified person|Other and unspecified water transport accident injuring other specified person
C0261313|T037|AB|E838.8|ICD9CM|Wtrcrft acc NEC-pers NEC|Wtrcrft acc NEC-pers NEC
C0261314|T037|PT|E838.9|ICD9CM|Other and unspecified water transport accident injuring unspecified person|Other and unspecified water transport accident injuring unspecified person
C0261314|T037|AB|E838.9|ICD9CM|Wtrcrft acc NEC-pers NOS|Wtrcrft acc NEC-pers NOS
C0261315|T037|HT|E840|ICD9CM|Accident to powered aircraft at takeoff or landing|Accident to powered aircraft at takeoff or landing
C0178350|T037|HT|E840-E845.9|ICD9CM|AIR AND SPACE TRANSPORT ACCIDENTS|AIR AND SPACE TRANSPORT ACCIDENTS
C0416143|T037|HT|E841|ICD9CM|Accident to powered aircraft, other and unspecified|Accident to powered aircraft, other and unspecified
C0261337|T037|HT|E842|ICD9CM|Accident to unpowered aircraft|Accident to unpowered aircraft
C0261342|T037|HT|E843|ICD9CM|Fall in, on, or from aircraft|Fall in, on, or from aircraft
C0261351|T037|AB|E843.8|ICD9CM|Aircrft fall-ground crew|Aircrft fall-ground crew
C0261351|T037|PT|E843.8|ICD9CM|Fall in, on, or from aircraft injuring ground crew, airline employee|Fall in, on, or from aircraft injuring ground crew, airline employee
C0261353|T037|HT|E844|ICD9CM|Other specified air transport accidents|Other specified air transport accidents
C0261371|T033|HT|E849-E849.9|ICD9CM|PLACE OF OCCURRENCE|PLACE OF OCCURRENCE
C0261377|T037|AB|E849.6|ICD9CM|Accident in public bldg|Accident in public bldg
C0261377|T037|PT|E849.6|ICD9CM|Accidents occurring in public building|Accidents occurring in public building
C0261378|T033|AB|E849.7|ICD9CM|Accid in resident instit|Accid in resident instit
C0261378|T033|PT|E849.7|ICD9CM|Accidents occurring in residential institution|Accidents occurring in residential institution
C0261381|T037|HT|E850|ICD9CM|Accidental poisoning by analgesics, antipyretics, and antirheumatics|Accidental poisoning by analgesics, antipyretics, and antirheumatics
C0178352|T037|HT|E850-E858.9|ICD9CM|ACCIDENTAL POISONING BY DRUGS, MEDICINAL SUBSTANCES, AND BIOLOGICALS|ACCIDENTAL POISONING BY DRUGS, MEDICINAL SUBSTANCES, AND BIOLOGICALS
C0261382|T037|AB|E850.0|ICD9CM|Acc poison-heroin|Acc poison-heroin
C0261382|T037|PT|E850.0|ICD9CM|Accidental poisoning by heroin|Accidental poisoning by heroin
C0261383|T037|AB|E850.1|ICD9CM|Acc poison-methadone|Acc poison-methadone
C0261383|T037|PT|E850.1|ICD9CM|Accidental poisoning by methadone|Accidental poisoning by methadone
C0261384|T037|AB|E850.2|ICD9CM|Acc poison-opiates NEC|Acc poison-opiates NEC
C0261384|T037|PT|E850.2|ICD9CM|Accidental poisoning by other opiates and related narcotics|Accidental poisoning by other opiates and related narcotics
C0261385|T037|AB|E850.3|ICD9CM|Acc poison-salicylates|Acc poison-salicylates
C0261385|T037|PT|E850.3|ICD9CM|Accidental poisoning by salicylates|Accidental poisoning by salicylates
C0869513|T037|AB|E850.4|ICD9CM|Acc poison-arom analgesc|Acc poison-arom analgesc
C0869513|T037|PT|E850.4|ICD9CM|Accidental poisoning by aromatic analgesics, not elsewhere classified|Accidental poisoning by aromatic analgesics, not elsewhere classified
C0261387|T037|AB|E850.5|ICD9CM|Acc poison-pyrazole derv|Acc poison-pyrazole derv
C0261387|T037|PT|E850.5|ICD9CM|Accidental poisoning by pyrazole derivatives|Accidental poisoning by pyrazole derivatives
C0416598|T037|AB|E850.6|ICD9CM|Acc poison-antirheumatic|Acc poison-antirheumatic
C0416598|T037|PT|E850.6|ICD9CM|Accidental poisoning by antirheumatics (antiphlogistics)|Accidental poisoning by antirheumatics (antiphlogistics)
C0261389|T037|AB|E850.7|ICD9CM|Acc poison-nonnarc analg|Acc poison-nonnarc analg
C0261389|T037|PT|E850.7|ICD9CM|Accidental poisoning by other non-narcotic analgesics|Accidental poisoning by other non-narcotic analgesics
C0261390|T037|AB|E850.8|ICD9CM|Acc poison-analgesic NEC|Acc poison-analgesic NEC
C0261390|T037|PT|E850.8|ICD9CM|Accidental poisoning by other specified analgesics and antipyretics|Accidental poisoning by other specified analgesics and antipyretics
C0261391|T037|AB|E850.9|ICD9CM|Acc poison-analgesic NOS|Acc poison-analgesic NOS
C0261391|T037|PT|E850.9|ICD9CM|Accidental poisoning by unspecified analgesic or antipyretic|Accidental poisoning by unspecified analgesic or antipyretic
C0261392|T037|AB|E851|ICD9CM|Acc poison-barbiturates|Acc poison-barbiturates
C0261392|T037|PT|E851|ICD9CM|Accidental poisoning by barbiturates|Accidental poisoning by barbiturates
C0261393|T037|HT|E852|ICD9CM|Accidental poisoning by other sedatives and hypnotics|Accidental poisoning by other sedatives and hypnotics
C0261394|T037|AB|E852.0|ICD9CM|Acc poisn-chlorl hydrate|Acc poisn-chlorl hydrate
C0261394|T037|PT|E852.0|ICD9CM|Accidental poisoning by chloral hydrate group|Accidental poisoning by chloral hydrate group
C0261395|T037|AB|E852.1|ICD9CM|Acc poison-paraldehyde|Acc poison-paraldehyde
C0261395|T037|PT|E852.1|ICD9CM|Accidental poisoning by paraldehyde|Accidental poisoning by paraldehyde
C0261396|T037|AB|E852.2|ICD9CM|Acc poison-bromine cmpnd|Acc poison-bromine cmpnd
C0261396|T037|PT|E852.2|ICD9CM|Accidental poisoning by bromine compounds|Accidental poisoning by bromine compounds
C0261397|T037|AB|E852.3|ICD9CM|Acc poison-methaqualone|Acc poison-methaqualone
C0261397|T037|PT|E852.3|ICD9CM|Accidental poisoning by methaqualone compounds|Accidental poisoning by methaqualone compounds
C0261398|T037|AB|E852.4|ICD9CM|Acc poison-glutethimide|Acc poison-glutethimide
C0261398|T037|PT|E852.4|ICD9CM|Accidental poisoning by glutethimide group|Accidental poisoning by glutethimide group
C0869445|T037|AB|E852.5|ICD9CM|Acc poison-mix sedtv NEC|Acc poison-mix sedtv NEC
C0869445|T037|PT|E852.5|ICD9CM|Accidental poisoning by mixed sedatives, not elsewhere classified|Accidental poisoning by mixed sedatives, not elsewhere classified
C0261400|T037|AB|E852.8|ICD9CM|Acc poison-sedatives NEC|Acc poison-sedatives NEC
C0261400|T037|PT|E852.8|ICD9CM|Accidental poisoning by other specified sedatives and hypnotics|Accidental poisoning by other specified sedatives and hypnotics
C0261401|T037|AB|E852.9|ICD9CM|Acc poison-sedatives NOS|Acc poison-sedatives NOS
C0261401|T037|PT|E852.9|ICD9CM|Accidental poisoning by unspecified sedative or hypnotic|Accidental poisoning by unspecified sedative or hypnotic
C0261402|T037|HT|E853|ICD9CM|Accidental poisoning by tranquilizers|Accidental poisoning by tranquilizers
C0261403|T037|AB|E853.0|ICD9CM|Acc pois-phenthiaz tranq|Acc pois-phenthiaz tranq
C0261403|T037|PT|E853.0|ICD9CM|Accidental poisoning by phenothiazine-based tranquilizers|Accidental poisoning by phenothiazine-based tranquilizers
C0261404|T037|AB|E853.1|ICD9CM|Acc pois-butyrphen tranq|Acc pois-butyrphen tranq
C0261404|T037|PT|E853.1|ICD9CM|Accidental poisoning by butyrophenone-based tranquilizers|Accidental poisoning by butyrophenone-based tranquilizers
C0261405|T037|AB|E853.2|ICD9CM|Acc poisn-benzdiaz tranq|Acc poisn-benzdiaz tranq
C0261405|T037|PT|E853.2|ICD9CM|Accidental poisoning by benzodiazepine-based tranquilizers|Accidental poisoning by benzodiazepine-based tranquilizers
C0261406|T037|AB|E853.8|ICD9CM|Acc poisn-tranquilzr NEC|Acc poisn-tranquilzr NEC
C0261406|T037|PT|E853.8|ICD9CM|Accidental poisoning by other specified tranquilizers|Accidental poisoning by other specified tranquilizers
C0261407|T037|AB|E853.9|ICD9CM|Acc poisn-tranquilzr NOS|Acc poisn-tranquilzr NOS
C0261407|T037|PT|E853.9|ICD9CM|Accidental poisoning by unspecified tranquilizer|Accidental poisoning by unspecified tranquilizer
C0261408|T037|HT|E854|ICD9CM|Accidental poisoning by other psychotropic agents|Accidental poisoning by other psychotropic agents
C0261409|T037|AB|E854.0|ICD9CM|Acc poison-antidepressnt|Acc poison-antidepressnt
C0261409|T037|PT|E854.0|ICD9CM|Accidental poisoning by antidepressants|Accidental poisoning by antidepressants
C0480040|T037|AB|E854.1|ICD9CM|Acc poison-hallucinogens|Acc poison-hallucinogens
C0480040|T037|PT|E854.1|ICD9CM|Accidental poisoning by psychodysleptics [hallucinogens]|Accidental poisoning by psychodysleptics [hallucinogens]
C0261411|T037|AB|E854.2|ICD9CM|Acc poisn-psychstimulant|Acc poisn-psychstimulant
C0261411|T037|PT|E854.2|ICD9CM|Accidental poisoning by psychostimulants|Accidental poisoning by psychostimulants
C0261412|T037|AB|E854.3|ICD9CM|Acc poison-cns stimulant|Acc poison-cns stimulant
C0261412|T037|PT|E854.3|ICD9CM|Accidental poisoning by central nervous system stimulants|Accidental poisoning by central nervous system stimulants
C0261408|T037|AB|E854.8|ICD9CM|Acc poisn psychotrop NEC|Acc poisn psychotrop NEC
C0261408|T037|PT|E854.8|ICD9CM|Accidental poisoning by other psychotropic agents|Accidental poisoning by other psychotropic agents
C0261413|T037|HT|E855|ICD9CM|Accidental poisoning by other drugs acting on central and autonomic nervous system|Accidental poisoning by other drugs acting on central and autonomic nervous system
C0261414|T037|AB|E855.0|ICD9CM|Acc poisn-anticonvulsant|Acc poisn-anticonvulsant
C0261414|T037|PT|E855.0|ICD9CM|Accidental poisoning by anticonvulsant and anti-parkinsonism drugs|Accidental poisoning by anticonvulsant and anti-parkinsonism drugs
C0261415|T037|AB|E855.1|ICD9CM|Acc poisn-cns depres NEC|Acc poisn-cns depres NEC
C0261415|T037|PT|E855.1|ICD9CM|Accidental poisoning by other central nervous system depressants|Accidental poisoning by other central nervous system depressants
C0261416|T037|AB|E855.2|ICD9CM|Acc poisn-local anesthet|Acc poisn-local anesthet
C0261416|T037|PT|E855.2|ICD9CM|Accidental poisoning by local anesthetics|Accidental poisoning by local anesthetics
C0416665|T037|AB|E855.3|ICD9CM|Acc poison-cholinergics|Acc poison-cholinergics
C0416665|T037|PT|E855.3|ICD9CM|Accidental poisoning by parasympathomimetics [cholinergics]|Accidental poisoning by parasympathomimetics [cholinergics]
C0261418|T037|AB|E855.4|ICD9CM|Acc poisn-anticholinerg|Acc poisn-anticholinerg
C0261418|T037|PT|E855.4|ICD9CM|Accidental poisoning by parasympatholytics [anticholinergics and antimuscarinics] and spasmolytics|Accidental poisoning by parasympatholytics [anticholinergics and antimuscarinics] and spasmolytics
C0416674|T037|AB|E855.5|ICD9CM|Acc poison-adrenergics|Acc poison-adrenergics
C0416674|T037|PT|E855.5|ICD9CM|Accidental poisoning by sympathomimetics [adrenergics]|Accidental poisoning by sympathomimetics [adrenergics]
C0416678|T037|AB|E855.6|ICD9CM|Acc poisn-sympatholytics|Acc poisn-sympatholytics
C0416678|T037|PT|E855.6|ICD9CM|Accidental poisoning by sympatholytics [antiadrenergics]|Accidental poisoning by sympatholytics [antiadrenergics]
C0261421|T037|AB|E855.8|ICD9CM|Acc poison-cns drug NEC|Acc poison-cns drug NEC
C0261421|T037|PT|E855.8|ICD9CM|Accidental poisoning by other specified drugs acting on central and autonomic nervous systems|Accidental poisoning by other specified drugs acting on central and autonomic nervous systems
C0261422|T037|AB|E855.9|ICD9CM|Acc poison-cns drug NOS|Acc poison-cns drug NOS
C0261422|T037|PT|E855.9|ICD9CM|Accidental poisoning by unspecified drug acting on central and autonomic nervous systems|Accidental poisoning by unspecified drug acting on central and autonomic nervous systems
C0261423|T037|AB|E856|ICD9CM|Acc poison-antibiotics|Acc poison-antibiotics
C0261423|T037|PT|E856|ICD9CM|Accidental poisoning by antibiotics|Accidental poisoning by antibiotics
C0261424|T037|AB|E857|ICD9CM|Acc pois-oth anti-infect|Acc pois-oth anti-infect
C0261424|T037|PT|E857|ICD9CM|Accidental poisoning by other anti-infectives|Accidental poisoning by other anti-infectives
C0261425|T037|HT|E858|ICD9CM|Accidental poisoning by other drugs|Accidental poisoning by other drugs
C0261426|T037|AB|E858.0|ICD9CM|Acc poison-hormones|Acc poison-hormones
C0261426|T037|PT|E858.0|ICD9CM|Accidental poisoning by hormones and synthetic substitutes|Accidental poisoning by hormones and synthetic substitutes
C0261427|T037|AB|E858.1|ICD9CM|Acc poisn-systemic agent|Acc poisn-systemic agent
C0261427|T037|PT|E858.1|ICD9CM|Accidental poisoning by primarily systemic agents|Accidental poisoning by primarily systemic agents
C0261428|T037|AB|E858.2|ICD9CM|Acc poison-blood agent|Acc poison-blood agent
C0261428|T037|PT|E858.2|ICD9CM|Accidental poisoning by agents primarily affecting blood constituents|Accidental poisoning by agents primarily affecting blood constituents
C0261429|T037|AB|E858.3|ICD9CM|Acc poisn-cardiovasc agt|Acc poisn-cardiovasc agt
C0261429|T037|PT|E858.3|ICD9CM|Accidental poisoning by agents primarily affecting cardiovascular system|Accidental poisoning by agents primarily affecting cardiovascular system
C0261430|T037|AB|E858.4|ICD9CM|Acc poison-gi agent|Acc poison-gi agent
C0261430|T037|PT|E858.4|ICD9CM|Accidental poisoning by agents primarily affecting gastrointestinal system|Accidental poisoning by agents primarily affecting gastrointestinal system
C0261431|T037|AB|E858.5|ICD9CM|Acc poisn-metabol agnt|Acc poisn-metabol agnt
C0261431|T037|PT|E858.5|ICD9CM|Accidental poisoning by water, mineral, and uric acid metabolism drugs|Accidental poisoning by water, mineral, and uric acid metabolism drugs
C0261432|T037|AB|E858.6|ICD9CM|Acc poisn-muscl/resp agt|Acc poisn-muscl/resp agt
C1384500|T033|AB|E858.7|ICD9CM|Acc poisn-skin/eent agnt|Acc poisn-skin/eent agnt
C0261434|T037|AB|E858.8|ICD9CM|Acc poisoning-drug NEC|Acc poisoning-drug NEC
C0261434|T037|PT|E858.8|ICD9CM|Accidental poisoning by other specified drugs|Accidental poisoning by other specified drugs
C0261435|T037|AB|E858.9|ICD9CM|Acc poisoning-drug NOS|Acc poisoning-drug NOS
C0261435|T037|PT|E858.9|ICD9CM|Accidental poisoning by unspecified drug|Accidental poisoning by unspecified drug
C0868867|T037|HT|E860|ICD9CM|Accidental poisoning by alcohol, not elsewhere classified|Accidental poisoning by alcohol, not elsewhere classified
C0178353|T037|HT|E860-E869.9|ICD9CM|ACCIDENTAL POISONING BY OTHER SOLID AND LIQUID SUBSTANCES, GASES, AND VAPORS|ACCIDENTAL POISONING BY OTHER SOLID AND LIQUID SUBSTANCES, GASES, AND VAPORS
C0261437|T037|AB|E860.0|ICD9CM|Acc poisn-alcohol bevrag|Acc poisn-alcohol bevrag
C0261437|T037|PT|E860.0|ICD9CM|Accidental poisoning by alcoholic beverages|Accidental poisoning by alcoholic beverages
C0261438|T037|AB|E860.1|ICD9CM|Acc poison-ethyl alcohol|Acc poison-ethyl alcohol
C0261438|T037|PT|E860.1|ICD9CM|Accidental poisoning by other and unspecified ethyl alcohol and its products|Accidental poisoning by other and unspecified ethyl alcohol and its products
C0261439|T037|AB|E860.2|ICD9CM|Acc poisn-methyl alcohol|Acc poisn-methyl alcohol
C0261439|T037|PT|E860.2|ICD9CM|Accidental poisoning by methyl alcohol|Accidental poisoning by methyl alcohol
C0261440|T037|AB|E860.3|ICD9CM|Acc poisn-isopropyl alc|Acc poisn-isopropyl alc
C0261440|T037|PT|E860.3|ICD9CM|Accidental poisoning by isopropyl alcohol|Accidental poisoning by isopropyl alcohol
C0261441|T037|AB|E860.4|ICD9CM|Acc poison-fusel oil|Acc poison-fusel oil
C0261441|T037|PT|E860.4|ICD9CM|Accidental poisoning by fusel oil|Accidental poisoning by fusel oil
C0261442|T037|AB|E860.8|ICD9CM|Acc poison-alcohol NEC|Acc poison-alcohol NEC
C0261442|T037|PT|E860.8|ICD9CM|Accidental poisoning by other specified alcohols|Accidental poisoning by other specified alcohols
C0480073|T037|AB|E860.9|ICD9CM|Acc poison-alcohol NOS|Acc poison-alcohol NOS
C0480073|T037|PT|E860.9|ICD9CM|Accidental poisoning by unspecified alcohol|Accidental poisoning by unspecified alcohol
C0261444|T037|HT|E861|ICD9CM|Accidental poisoning by cleansing and polishing agents, disinfectants, paints, and varnishes|Accidental poisoning by cleansing and polishing agents, disinfectants, paints, and varnishes
C0261445|T037|AB|E861.0|ICD9CM|Acc pois-synth detergent|Acc pois-synth detergent
C0261445|T037|PT|E861.0|ICD9CM|Accidental poisoning by synthetic detergents and shampoos|Accidental poisoning by synthetic detergents and shampoos
C0261446|T037|AB|E861.1|ICD9CM|Acc poison-soap products|Acc poison-soap products
C0261446|T037|PT|E861.1|ICD9CM|Accidental poisoning by soap products|Accidental poisoning by soap products
C0261447|T037|AB|E861.2|ICD9CM|Acc poison-polishes|Acc poison-polishes
C0261447|T037|PT|E861.2|ICD9CM|Accidental poisoning by polishes|Accidental poisoning by polishes
C0416707|T037|AB|E861.3|ICD9CM|Acc poison-cleanser NEC|Acc poison-cleanser NEC
C0416707|T037|PT|E861.3|ICD9CM|Accidental poisoning by other cleansing and polishing agents|Accidental poisoning by other cleansing and polishing agents
C0261449|T037|AB|E861.4|ICD9CM|Acc poison-disinfectants|Acc poison-disinfectants
C0261449|T037|PT|E861.4|ICD9CM|Accidental poisoning by disinfectants|Accidental poisoning by disinfectants
C0261450|T037|AB|E861.5|ICD9CM|Acc poison-lead paints|Acc poison-lead paints
C0261450|T037|PT|E861.5|ICD9CM|Accidental poisoning by lead paints|Accidental poisoning by lead paints
C0261451|T037|AB|E861.6|ICD9CM|Acc poison-paints NEC|Acc poison-paints NEC
C0261451|T037|PT|E861.6|ICD9CM|Accidental poisoning by other paints and varnishes|Accidental poisoning by other paints and varnishes
C0261452|T037|AB|E861.9|ICD9CM|Acc poison-cleanser NOS|Acc poison-cleanser NOS
C0261454|T037|AB|E862.0|ICD9CM|Acc poisn-petrol solvent|Acc poisn-petrol solvent
C0261454|T037|PT|E862.0|ICD9CM|Accidental poisoning by petroleum solvents|Accidental poisoning by petroleum solvents
C0416882|T037|AB|E862.1|ICD9CM|Acc poisn-petroleum fuel|Acc poisn-petroleum fuel
C0416882|T037|PT|E862.1|ICD9CM|Accidental poisoning by petroleum fuels and cleaners|Accidental poisoning by petroleum fuels and cleaners
C0261456|T037|AB|E862.2|ICD9CM|Acc pois-lubricating oil|Acc pois-lubricating oil
C0261456|T037|PT|E862.2|ICD9CM|Accidental poisoning by lubricating oils|Accidental poisoning by lubricating oils
C0261457|T037|AB|E862.3|ICD9CM|Acc pois-petroleum solid|Acc pois-petroleum solid
C0261457|T037|PT|E862.3|ICD9CM|Accidental poisoning by petroleum solids|Accidental poisoning by petroleum solids
C0302441|T037|AB|E862.4|ICD9CM|Acc poisn-solvents NEC|Acc poisn-solvents NEC
C0302441|T037|PT|E862.4|ICD9CM|Accidental poisoning by other specified solvents, not elsewhere classified|Accidental poisoning by other specified solvents, not elsewhere classified
C0302442|T037|AB|E862.9|ICD9CM|Acc poisn-solvent NOS|Acc poisn-solvent NOS
C0302442|T037|PT|E862.9|ICD9CM|Accidental poisoning by unspecified solvent, not elsewhere classified|Accidental poisoning by unspecified solvent, not elsewhere classified
C0261461|T037|AB|E863.0|ICD9CM|Acc pois-chlorine pestic|Acc pois-chlorine pestic
C0261461|T037|PT|E863.0|ICD9CM|Accidental poisoning by insecticides of organochlorine compounds|Accidental poisoning by insecticides of organochlorine compounds
C0261462|T037|AB|E863.1|ICD9CM|Acc pois-phosph pesticid|Acc pois-phosph pesticid
C0261462|T037|PT|E863.1|ICD9CM|Accidental poisoning by insecticides of organophosphorus compounds|Accidental poisoning by insecticides of organophosphorus compounds
C0261463|T037|AB|E863.2|ICD9CM|Acc poison-carbamates|Acc poison-carbamates
C0261463|T037|PT|E863.2|ICD9CM|Accidental poisoning by carbamates|Accidental poisoning by carbamates
C0261464|T037|AB|E863.3|ICD9CM|Acc poisn-mixed pesticid|Acc poisn-mixed pesticid
C0261464|T037|PT|E863.3|ICD9CM|Accidental poisoning by mixtures of insecticides|Accidental poisoning by mixtures of insecticides
C0261465|T037|AB|E863.4|ICD9CM|Acc poison-pesticide NEC|Acc poison-pesticide NEC
C0261465|T037|PT|E863.4|ICD9CM|Accidental poisoning by other and unspecified insecticides|Accidental poisoning by other and unspecified insecticides
C0261466|T037|AB|E863.5|ICD9CM|Acc poison-herbicides|Acc poison-herbicides
C0261466|T037|PT|E863.5|ICD9CM|Accidental poisoning by herbicides|Accidental poisoning by herbicides
C0261467|T037|AB|E863.6|ICD9CM|Acc poison-fungicides|Acc poison-fungicides
C0261467|T037|PT|E863.6|ICD9CM|Accidental poisoning by fungicides|Accidental poisoning by fungicides
C0261468|T037|AB|E863.7|ICD9CM|Acc poison-rodenticides|Acc poison-rodenticides
C0261468|T037|PT|E863.7|ICD9CM|Accidental poisoning by rodenticides|Accidental poisoning by rodenticides
C0261469|T037|AB|E863.8|ICD9CM|Acc poison-fumigants|Acc poison-fumigants
C0261469|T037|PT|E863.8|ICD9CM|Accidental poisoning by fumigants|Accidental poisoning by fumigants
C0261470|T037|AB|E863.9|ICD9CM|Acc pois-agrcult NEC/NOS|Acc pois-agrcult NEC/NOS
C0869267|T037|HT|E864|ICD9CM|Accidental poisoning by corrosives and caustics, not elsewhere classified|Accidental poisoning by corrosives and caustics, not elsewhere classified
C0302444|T037|AB|E864.0|ICD9CM|Acc pois-corrosiv aromat|Acc pois-corrosiv aromat
C0302444|T037|PT|E864.0|ICD9CM|Accidental poisoning by corrosive aromatics not elsewhere classified|Accidental poisoning by corrosive aromatics not elsewhere classified
C0302445|T037|AB|E864.1|ICD9CM|Acc poison-acids|Acc poison-acids
C0302445|T037|PT|E864.1|ICD9CM|Accidental poisoning by acids not elsewhere classified|Accidental poisoning by acids not elsewhere classified
C0302446|T037|AB|E864.2|ICD9CM|Acc poisn-caustic alkali|Acc poisn-caustic alkali
C0302446|T037|PT|E864.2|ICD9CM|Accidental poisoning by caustic alkalis not elsewhere classified|Accidental poisoning by caustic alkalis not elsewhere classified
C0302447|T037|AB|E864.3|ICD9CM|Acc poison-caustic NEC|Acc poison-caustic NEC
C0302447|T037|PT|E864.3|ICD9CM|Accidental poisoning by other specified corrosives and caustics not elsewhere classified|Accidental poisoning by other specified corrosives and caustics not elsewhere classified
C0302448|T037|AB|E864.4|ICD9CM|Acc poison-caustic NOS|Acc poison-caustic NOS
C0302448|T037|PT|E864.4|ICD9CM|Accidental poisoning by unspecified corrosives and caustics not elsewhere classified|Accidental poisoning by unspecified corrosives and caustics not elsewhere classified
C0375733|T037|HT|E865|ICD9CM|Accidental poisoning from poisonous foodstuffs and poisonous plants|Accidental poisoning from poisonous foodstuffs and poisonous plants
C0416786|T037|AB|E865.0|ICD9CM|Acc poison-meat|Acc poison-meat
C0416786|T037|PT|E865.0|ICD9CM|Accidental poisoning by meat|Accidental poisoning by meat
C0261479|T037|AB|E865.1|ICD9CM|Acc poison-shellfish|Acc poison-shellfish
C0261479|T037|PT|E865.1|ICD9CM|Accidental poisoning by shellfish|Accidental poisoning by shellfish
C0000923|T037|AB|E865.2|ICD9CM|Acc poison-fish NEC|Acc poison-fish NEC
C0000923|T037|PT|E865.2|ICD9CM|Accidental poisoning from other fish|Accidental poisoning from other fish
C1535481|T037|AB|E865.3|ICD9CM|Acc poison-berries/seeds|Acc poison-berries/seeds
C1535481|T037|PT|E865.3|ICD9CM|Accidental poisoning from berries and seeds|Accidental poisoning from berries and seeds
C0261481|T037|AB|E865.4|ICD9CM|Acc poison-plants NEC|Acc poison-plants NEC
C0261481|T037|PT|E865.4|ICD9CM|Accidental poisoning from other specified plants|Accidental poisoning from other specified plants
C0261482|T037|AB|E865.5|ICD9CM|Acc poison-mushrooms|Acc poison-mushrooms
C0261482|T037|PT|E865.5|ICD9CM|Accidental poisoning from mushrooms and other fungi|Accidental poisoning from mushrooms and other fungi
C0261483|T037|AB|E865.8|ICD9CM|Acc poison-food NEC|Acc poison-food NEC
C0261483|T037|PT|E865.8|ICD9CM|Accidental poisoning from other specified foods|Accidental poisoning from other specified foods
C0261484|T037|AB|E865.9|ICD9CM|Acc poisn-food/plant NOS|Acc poisn-food/plant NOS
C0261484|T037|PT|E865.9|ICD9CM|Accidental poisoning from unspecified foodstuff or poisonous plant|Accidental poisoning from unspecified foodstuff or poisonous plant
C0261485|T037|HT|E866|ICD9CM|Accidental poisoning by other and unspecified solid and liquid substances|Accidental poisoning by other and unspecified solid and liquid substances
C0261486|T037|AB|E866.0|ICD9CM|Acc poisoning-lead|Acc poisoning-lead
C0261486|T037|PT|E866.0|ICD9CM|Accidental poisoning by lead and its compounds and fumes|Accidental poisoning by lead and its compounds and fumes
C0261487|T037|AB|E866.1|ICD9CM|Acc poisoning-mercury|Acc poisoning-mercury
C0261487|T037|PT|E866.1|ICD9CM|Accidental poisoning by mercury and its compounds and fumes|Accidental poisoning by mercury and its compounds and fumes
C0261488|T037|AB|E866.2|ICD9CM|Acc poisoning-antimony|Acc poisoning-antimony
C0261488|T037|PT|E866.2|ICD9CM|Accidental poisoning by antimony and its compounds and fumes|Accidental poisoning by antimony and its compounds and fumes
C0261489|T037|AB|E866.3|ICD9CM|Acc poisoning-arsenic|Acc poisoning-arsenic
C0261489|T037|PT|E866.3|ICD9CM|Accidental poisoning by arsenic and its compounds and fumes|Accidental poisoning by arsenic and its compounds and fumes
C0261490|T037|AB|E866.4|ICD9CM|Acc poison-metals NEC|Acc poison-metals NEC
C0261490|T037|PT|E866.4|ICD9CM|Accidental poisoning by other metals and their compounds and fumes|Accidental poisoning by other metals and their compounds and fumes
C0261491|T037|AB|E866.5|ICD9CM|Acc poison-plant food|Acc poison-plant food
C0261491|T037|PT|E866.5|ICD9CM|Accidental poisoning by plant foods and fertilizers|Accidental poisoning by plant foods and fertilizers
C0261492|T037|AB|E866.6|ICD9CM|Acc poison-glues|Acc poison-glues
C0261492|T037|PT|E866.6|ICD9CM|Accidental poisoning by glues and adhesives|Accidental poisoning by glues and adhesives
C0261493|T037|AB|E866.7|ICD9CM|Acc poison-cosmetics|Acc poison-cosmetics
C0261493|T037|PT|E866.7|ICD9CM|Accidental poisoning by cosmetics|Accidental poisoning by cosmetics
C0261494|T037|AB|E866.8|ICD9CM|Acc pois-solid/liq NEC|Acc pois-solid/liq NEC
C0261494|T037|PT|E866.8|ICD9CM|Accidental poisoning by other specified solid or liquid substances|Accidental poisoning by other specified solid or liquid substances
C0261495|T037|AB|E866.9|ICD9CM|Acc pois-solid/liq NOS|Acc pois-solid/liq NOS
C0261495|T037|PT|E866.9|ICD9CM|Accidental poisoning by unspecified solid or liquid substance|Accidental poisoning by unspecified solid or liquid substance
C0261496|T037|AB|E867|ICD9CM|Acc poison-piped gas|Acc poison-piped gas
C0261496|T037|PT|E867|ICD9CM|Accidental poisoning by gas distributed by pipeline|Accidental poisoning by gas distributed by pipeline
C0261497|T037|HT|E868|ICD9CM|Accidental poisoning by other utility gas and other carbon monoxide|Accidental poisoning by other utility gas and other carbon monoxide
C0261498|T037|AB|E868.0|ICD9CM|Acc pois-liq petrol gas|Acc pois-liq petrol gas
C0261498|T037|PT|E868.0|ICD9CM|Accidental poisoning by liquefied petroleum gas distributed in mobile containers|Accidental poisoning by liquefied petroleum gas distributed in mobile containers
C0261499|T037|AB|E868.1|ICD9CM|Acc pois-utl gas NEC/NOS|Acc pois-utl gas NEC/NOS
C0261499|T037|PT|E868.1|ICD9CM|Accidental poisoning by other and unspecified utility gas|Accidental poisoning by other and unspecified utility gas
C0261500|T037|AB|E868.2|ICD9CM|Acc poison-exhaust gas|Acc poison-exhaust gas
C0261500|T037|PT|E868.2|ICD9CM|Accidental poisoning by motor vehicle exhaust gas|Accidental poisoning by motor vehicle exhaust gas
C0261501|T037|AB|E868.3|ICD9CM|Acc pois-co/domestc fuel|Acc pois-co/domestc fuel
C0261501|T037|PT|E868.3|ICD9CM|Accidental poisoning by carbon monoxide from incomplete combustion of other domestic fuels|Accidental poisoning by carbon monoxide from incomplete combustion of other domestic fuels
C0261502|T037|AB|E868.8|ICD9CM|Acc pois-carbn monox NEC|Acc pois-carbn monox NEC
C0261502|T037|PT|E868.8|ICD9CM|Accidental poisoning by carbon monoxide from other sources|Accidental poisoning by carbon monoxide from other sources
C0261503|T037|AB|E868.9|ICD9CM|Acc pois-carbn monox NOS|Acc pois-carbn monox NOS
C0261503|T037|PT|E868.9|ICD9CM|Accidental poisoning by unspecified carbon monoxide|Accidental poisoning by unspecified carbon monoxide
C0261504|T037|HT|E869|ICD9CM|Accidental poisoning by other gases and vapors|Accidental poisoning by other gases and vapors
C0261505|T037|AB|E869.0|ICD9CM|Acc poisn-nitrogen oxide|Acc poisn-nitrogen oxide
C0261505|T037|PT|E869.0|ICD9CM|Accidental poisoning by nitrogen oxides|Accidental poisoning by nitrogen oxides
C0261506|T037|AB|E869.1|ICD9CM|Acc poisn-sulfur dioxide|Acc poisn-sulfur dioxide
C0261506|T037|PT|E869.1|ICD9CM|Accidental poisoning by sulfur dioxide|Accidental poisoning by sulfur dioxide
C0261507|T037|AB|E869.2|ICD9CM|Acc poison-freon|Acc poison-freon
C0261507|T037|PT|E869.2|ICD9CM|Accidental poisoning by freon|Accidental poisoning by freon
C0416973|T037|AB|E869.3|ICD9CM|Acc poison-tear gas|Acc poison-tear gas
C0416973|T037|PT|E869.3|ICD9CM|Accidental poisoning by lacrimogenic gas [tear gas]|Accidental poisoning by lacrimogenic gas [tear gas]
C0375734|T037|AB|E869.4|ICD9CM|Scndhnd tbcco smoke|Scndhnd tbcco smoke
C0375734|T037|PT|E869.4|ICD9CM|Second hand tobacco smoke|Second hand tobacco smoke
C0261509|T037|AB|E869.8|ICD9CM|Acc poison-gas/vapor NEC|Acc poison-gas/vapor NEC
C0261509|T037|PT|E869.8|ICD9CM|Accidental poisoning by other specified gases and vapors|Accidental poisoning by other specified gases and vapors
C0261510|T037|AB|E869.9|ICD9CM|Acc poison-gas/vapor NOS|Acc poison-gas/vapor NOS
C0261510|T037|PT|E869.9|ICD9CM|Accidental poisoning by unspecified gases and vapors|Accidental poisoning by unspecified gases and vapors
C0261513|T037|HT|E870|ICD9CM|Accidental cut, puncture, perforation, or hemorrhage during medical care|Accidental cut, puncture, perforation, or hemorrhage during medical care
C0481263|T037|HT|E870-E876.9|ICD9CM|MISADVENTURES TO PATIENTS DURING SURGICAL AND MEDICAL CARE|MISADVENTURES TO PATIENTS DURING SURGICAL AND MEDICAL CARE
C0481222|T037|AB|E870.0|ICD9CM|Acc cut/hem in surgery|Acc cut/hem in surgery
C0481222|T037|PT|E870.0|ICD9CM|Accidental cut, puncture, perforation or hemorrhage during surgical operation|Accidental cut, puncture, perforation or hemorrhage during surgical operation
C2939422|T037|AB|E870.1|ICD9CM|Acc cut/hem in infusion|Acc cut/hem in infusion
C2939422|T037|PT|E870.1|ICD9CM|Accidental cut, puncture, perforation or hemorrhage during infusion or transfusion|Accidental cut, puncture, perforation or hemorrhage during infusion or transfusion
C0261514|T037|AB|E870.2|ICD9CM|Acc cut/hem-perfusn NEC|Acc cut/hem-perfusn NEC
C0261514|T037|PT|E870.2|ICD9CM|Accidental cut, puncture, perforation or hemorrhage during kidney dialysis or other perfusion|Accidental cut, puncture, perforation or hemorrhage during kidney dialysis or other perfusion
C0261515|T037|AB|E870.3|ICD9CM|Acc cut/hem in injection|Acc cut/hem in injection
C0261515|T037|PT|E870.3|ICD9CM|Accidental cut, puncture, perforation or hemorrhage during injection or vaccination|Accidental cut, puncture, perforation or hemorrhage during injection or vaccination
C0261516|T037|AB|E870.4|ICD9CM|Acc cut/hem w scope exam|Acc cut/hem w scope exam
C0261516|T037|PT|E870.4|ICD9CM|Accidental cut, puncture, perforation or hemorrhage during endoscopic examination|Accidental cut, puncture, perforation or hemorrhage during endoscopic examination
C0261517|T037|AB|E870.5|ICD9CM|Acc cut/hem w catheteriz|Acc cut/hem w catheteriz
C0261518|T037|AB|E870.6|ICD9CM|Acc cut/hem w heart cath|Acc cut/hem w heart cath
C0261518|T037|PT|E870.6|ICD9CM|Accidental cut, puncture, perforation or hemorrhage during heart catheterization|Accidental cut, puncture, perforation or hemorrhage during heart catheterization
C0261519|T037|AB|E870.7|ICD9CM|Acc cut/hem w enema|Acc cut/hem w enema
C0261519|T037|PT|E870.7|ICD9CM|Accidental cut, puncture, perforation or hemorrhage during administration of enema|Accidental cut, puncture, perforation or hemorrhage during administration of enema
C0261520|T037|AB|E870.8|ICD9CM|Acc cut in med care NEC|Acc cut in med care NEC
C0261520|T037|PT|E870.8|ICD9CM|Accidental cut, puncture, perforation or hemorrhage during other specified medical care|Accidental cut, puncture, perforation or hemorrhage during other specified medical care
C0261513|T037|AB|E870.9|ICD9CM|Acc cut in med care NOS|Acc cut in med care NOS
C0261513|T037|PT|E870.9|ICD9CM|Accidental cut, puncture, perforation or hemorrhage during unspecified medical care|Accidental cut, puncture, perforation or hemorrhage during unspecified medical care
C0261522|T037|HT|E871|ICD9CM|Foreign object left in body during procedure|Foreign object left in body during procedure
C0702090|T037|PT|E871.0|ICD9CM|Foreign object left in body during surgical operation|Foreign object left in body during surgical operation
C0702090|T037|AB|E871.0|ICD9CM|Post-surgical forgn body|Post-surgical forgn body
C0481232|T037|PT|E871.1|ICD9CM|Foreign object left in body during infusion or transfusion|Foreign object left in body during infusion or transfusion
C0481232|T037|AB|E871.1|ICD9CM|Postinfusion foreign bdy|Postinfusion foreign bdy
C0481233|T037|PT|E871.2|ICD9CM|Foreign object left in body during kidney dialysis or other perfusion|Foreign object left in body during kidney dialysis or other perfusion
C0481233|T037|AB|E871.2|ICD9CM|Postperfusion forgn body|Postperfusion forgn body
C0481234|T037|PT|E871.3|ICD9CM|Foreign object left in body during injection or vaccination|Foreign object left in body during injection or vaccination
C0481234|T037|AB|E871.3|ICD9CM|Postinjection forgn body|Postinjection forgn body
C0481235|T037|PT|E871.4|ICD9CM|Foreign object left in body during endoscopic examination|Foreign object left in body during endoscopic examination
C0481235|T037|AB|E871.4|ICD9CM|Postendoscopy forgn body|Postendoscopy forgn body
C0481237|T037|PT|E871.5|ICD9CM|Foreign object left in body during aspiration of fluid or tissue, puncture, and catheterization|Foreign object left in body during aspiration of fluid or tissue, puncture, and catheterization
C0481237|T037|AB|E871.5|ICD9CM|Postcatheter forgn body|Postcatheter forgn body
C0481236|T037|AB|E871.6|ICD9CM|FB post heart catheter|FB post heart catheter
C0481236|T037|PT|E871.6|ICD9CM|Foreign object left in body during heart catheterization|Foreign object left in body during heart catheterization
C0496530|T037|AB|E871.7|ICD9CM|FB post-catheter removal|FB post-catheter removal
C0496530|T037|PT|E871.7|ICD9CM|Foreign object left in body during removal of catheter or packing|Foreign object left in body during removal of catheter or packing
C0261531|T037|PT|E871.8|ICD9CM|Foreign object left in body during other specified procedures|Foreign object left in body during other specified procedures
C0261531|T037|AB|E871.8|ICD9CM|Post-op foreign body NEC|Post-op foreign body NEC
C0261532|T037|PT|E871.9|ICD9CM|Foreign object left in body during unspecified procedure|Foreign object left in body during unspecified procedure
C0261532|T037|AB|E871.9|ICD9CM|Post-op foreign body NOS|Post-op foreign body NOS
C0261533|T037|HT|E872|ICD9CM|Failure of sterile precautions during procedure|Failure of sterile precautions during procedure
C0261533|T037|PT|E872.0|ICD9CM|Failure of sterile precautions during surgical operation|Failure of sterile precautions during surgical operation
C0261533|T037|AB|E872.0|ICD9CM|Failure sterile surgery|Failure sterile surgery
C0497080|T037|PT|E872.1|ICD9CM|Failure of sterile precautions during infusion or transfusion|Failure of sterile precautions during infusion or transfusion
C0497080|T037|AB|E872.1|ICD9CM|Failure sterile infusion|Failure sterile infusion
C0261536|T037|AB|E872.2|ICD9CM|Fail sterile perfusn NEC|Fail sterile perfusn NEC
C0261536|T037|PT|E872.2|ICD9CM|Failure of sterile precautions during kidney dialysis and other perfusion|Failure of sterile precautions during kidney dialysis and other perfusion
C0497081|T037|AB|E872.3|ICD9CM|Fail sterile injection|Fail sterile injection
C0497081|T037|PT|E872.3|ICD9CM|Failure of sterile precautions during injection or vaccination|Failure of sterile precautions during injection or vaccination
C0497082|T037|AB|E872.4|ICD9CM|Fail sterile endoscopy|Fail sterile endoscopy
C0497082|T037|PT|E872.4|ICD9CM|Failure of sterile precautions during endoscopic examination|Failure of sterile precautions during endoscopic examination
C0261539|T037|AB|E872.5|ICD9CM|Fail sterile catheter|Fail sterile catheter
C0261539|T037|PT|E872.5|ICD9CM|Failure of sterile precautions during aspiration of fluid or tissue, puncture, and catheterization|Failure of sterile precautions during aspiration of fluid or tissue, puncture, and catheterization
C0497083|T037|AB|E872.6|ICD9CM|Fail sterile heart cath|Fail sterile heart cath
C0497083|T037|PT|E872.6|ICD9CM|Failure of sterile precautions during heart catheterization|Failure of sterile precautions during heart catheterization
C0261541|T033|AB|E872.8|ICD9CM|Fail sterile proced NEC|Fail sterile proced NEC
C0261541|T033|PT|E872.8|ICD9CM|Failure of sterile precautions during other specified procedures|Failure of sterile precautions during other specified procedures
C0261542|T033|AB|E872.9|ICD9CM|Fail sterile proced NOS|Fail sterile proced NOS
C0261542|T033|PT|E872.9|ICD9CM|Failure of sterile precautions during unspecified procedure|Failure of sterile precautions during unspecified procedure
C0261543|T033|HT|E873|ICD9CM|Failure in dosage|Failure in dosage
C0481246|T037|AB|E873.0|ICD9CM|Excess fluid in infusion|Excess fluid in infusion
C0481246|T037|PT|E873.0|ICD9CM|Excessive amount of blood or other fluid during transfusion or infusion|Excessive amount of blood or other fluid during transfusion or infusion
C0481247|T037|AB|E873.1|ICD9CM|Incor dilut infusn fluid|Incor dilut infusn fluid
C0481247|T037|PT|E873.1|ICD9CM|Incorrect dilution of fluid during infusion|Incorrect dilution of fluid during infusion
C0481248|T037|PT|E873.2|ICD9CM|Overdose of radiation in therapy|Overdose of radiation in therapy
C0481248|T037|AB|E873.2|ICD9CM|Therap radiation overdos|Therap radiation overdos
C0261547|T037|AB|E873.3|ICD9CM|Inadv radiat exp-medical|Inadv radiat exp-medical
C0261547|T037|PT|E873.3|ICD9CM|Inadvertent exposure of patient to radiation during medical care|Inadvertent exposure of patient to radiation during medical care
C0261548|T037|AB|E873.4|ICD9CM|Dosag fail-shock therapy|Dosag fail-shock therapy
C0261548|T037|PT|E873.4|ICD9CM|Failure in dosage in electroshock or insulin-shock therapy|Failure in dosage in electroshock or insulin-shock therapy
C0418626|T037|PT|E873.5|ICD9CM|Inappropriate [too hot or too cold] temperature in local application and packing|Inappropriate [too hot or too cold] temperature in local application and packing
C0418626|T037|AB|E873.5|ICD9CM|Wrng temp in applic/pack|Wrng temp in applic/pack
C0418624|T033|AB|E873.6|ICD9CM|Nonadmin necess medicine|Nonadmin necess medicine
C0418624|T033|PT|E873.6|ICD9CM|Nonadministration of necessary drug or medicinal substance|Nonadministration of necessary drug or medicinal substance
C0261551|T033|AB|E873.8|ICD9CM|Failure in dosage NEC|Failure in dosage NEC
C0261551|T033|PT|E873.8|ICD9CM|Other specified failure in dosage|Other specified failure in dosage
C0261543|T033|AB|E873.9|ICD9CM|Failure in dosage NOS|Failure in dosage NOS
C0261543|T033|PT|E873.9|ICD9CM|Unspecified failure in dosage|Unspecified failure in dosage
C0261553|T037|HT|E874|ICD9CM|Mechanical failure of instrument or apparatus during procedure|Mechanical failure of instrument or apparatus during procedure
C0261554|T037|AB|E874.0|ICD9CM|Instrmnt fail in surgery|Instrmnt fail in surgery
C0261554|T037|PT|E874.0|ICD9CM|Mechanical failure of instrument or apparatus during surgical operation|Mechanical failure of instrument or apparatus during surgical operation
C0261557|T037|AB|E874.3|ICD9CM|Instrumnt fail-endoscopy|Instrumnt fail-endoscopy
C0261557|T037|PT|E874.3|ICD9CM|Mechanical failure of instrument or apparatus during endoscopic examination|Mechanical failure of instrument or apparatus during endoscopic examination
C0261558|T037|AB|E874.4|ICD9CM|Instrmnt fail-catheteriz|Instrmnt fail-catheteriz
C0261559|T037|AB|E874.5|ICD9CM|Instrmnt fail-heart cath|Instrmnt fail-heart cath
C0261559|T037|PT|E874.5|ICD9CM|Mechanical failure of instrument or apparatus during heart catheterization|Mechanical failure of instrument or apparatus during heart catheterization
C0481253|T037|PT|E875.0|ICD9CM|Contaminated substance transfused or infused|Contaminated substance transfused or infused
C0481253|T037|AB|E875.0|ICD9CM|Contaminated transfusion|Contaminated transfusion
C0481254|T037|AB|E875.1|ICD9CM|Contaminated injection|Contaminated injection
C0481254|T037|PT|E875.1|ICD9CM|Contaminated substance injected or used for vaccination|Contaminated substance injected or used for vaccination
C0261567|T037|AB|E875.9|ICD9CM|Contamination NOS|Contamination NOS
C0261567|T037|PT|E875.9|ICD9CM|Misadventure to patient from unspecified contamination|Misadventure to patient from unspecified contamination
C0161841|T037|AB|E876.0|ICD9CM|Mismatch blood-transfusn|Mismatch blood-transfusn
C0161841|T037|PT|E876.0|ICD9CM|Mismatched blood in transfusion|Mismatched blood in transfusion
C0261570|T033|AB|E876.1|ICD9CM|Wrong fluid in infusion|Wrong fluid in infusion
C0261570|T033|PT|E876.1|ICD9CM|Wrong fluid in infusion|Wrong fluid in infusion
C0481259|T037|AB|E876.2|ICD9CM|Failure in suture|Failure in suture
C0481259|T037|PT|E876.2|ICD9CM|Failure in suture and ligature during surgical operation|Failure in suture and ligature during surgical operation
C0261572|T037|PT|E876.3|ICD9CM|Endotracheal tube wrongly placed during anesthetic procedure|Endotracheal tube wrongly placed during anesthetic procedure
C0261572|T037|AB|E876.3|ICD9CM|Misplaced endotrach tube|Misplaced endotrach tube
C0261573|T037|AB|E876.4|ICD9CM|Fail introd/remove tube|Fail introd/remove tube
C0261573|T037|PT|E876.4|ICD9CM|Failure to introduce or to remove other tube or instrument|Failure to introduce or to remove other tube or instrument
C2712478|T037|PT|E876.5|ICD9CM|Performance of wrong operation (procedure) on correct patient|Performance of wrong operation (procedure) on correct patient
C2712478|T037|AB|E876.5|ICD9CM|Perfrm wrong op/right pt|Perfrm wrong op/right pt
C2712479|T037|PT|E876.6|ICD9CM|Performance of operation (procedure) on patient not scheduled for surgery|Performance of operation (procedure) on patient not scheduled for surgery
C2712479|T037|AB|E876.6|ICD9CM|Proc-pt not sched surg|Proc-pt not sched surg
C2712480|T037|PT|E876.7|ICD9CM|Performance of correct operation (procedure) on wrong side/body part|Performance of correct operation (procedure) on wrong side/body part
C2712480|T037|AB|E876.7|ICD9CM|Rt proc-wrong side/part|Rt proc-wrong side/part
C0418593|T037|AB|E876.9|ICD9CM|Medical misadventure NOS|Medical misadventure NOS
C0418593|T037|PT|E876.9|ICD9CM|Unspecified misadventure during medical care|Unspecified misadventure during medical care
C0496542|T037|AB|E878.3|ICD9CM|Abn react-external stoma|Abn react-external stoma
C0418696|T037|AB|E878.4|ICD9CM|Abn react-plast surg NEC|Abn react-plast surg NEC
C0418697|T046|AB|E878.5|ICD9CM|Abn react-limb amputat|Abn react-limb amputat
C0261586|T037|AB|E878.9|ICD9CM|Abn react-surg proc NOS|Abn react-surg proc NOS
C0261588|T037|AB|E879.0|ICD9CM|Abn react-cardiac cath|Abn react-cardiac cath
C0261589|T037|AB|E879.1|ICD9CM|Abn react-renal dialysis|Abn react-renal dialysis
C0261590|T037|AB|E879.2|ICD9CM|Abn react-radiotherapy|Abn react-radiotherapy
C0261591|T037|AB|E879.3|ICD9CM|Abn react-shock therapy|Abn react-shock therapy
C0261592|T037|AB|E879.4|ICD9CM|Abn react-fluid aspirat|Abn react-fluid aspirat
C0481350|T037|AB|E879.5|ICD9CM|Abn react-gastric sound|Abn react-gastric sound
C0261594|T037|AB|E879.6|ICD9CM|Abn react-urinary cath|Abn react-urinary cath
C0261595|T037|AB|E879.7|ICD9CM|Abn react-blood sampling|Abn react-blood sampling
C0261596|T037|AB|E879.8|ICD9CM|Abn react-procedure NEC|Abn react-procedure NEC
C0261597|T037|AB|E879.9|ICD9CM|Abn react-procedure NOS|Abn react-procedure NOS
C0000921|T037|HT|E880-E888.9|ICD9CM|ACCIDENTAL FALLS|ACCIDENTAL FALLS
C0337212|T033|PT|E881.0|ICD9CM|Accidental fall from ladder|Accidental fall from ladder
C0337212|T033|AB|E881.0|ICD9CM|Fall from ladder|Fall from ladder
C0478874|T037|HT|E884|ICD9CM|Other accidental falls from one level to another|Other accidental falls from one level to another
C0337231|T037|PT|E884.3|ICD9CM|Accidental fall from wheelchair|Accidental fall from wheelchair
C0337231|T037|AB|E884.3|ICD9CM|Fall from wheelchair|Fall from wheelchair
C0337228|T037|PT|E884.4|ICD9CM|Accidental fall from bed|Accidental fall from bed
C0337228|T037|AB|E884.4|ICD9CM|Fall from bed|Fall from bed
C0375736|T037|PT|E884.5|ICD9CM|Accidental fall from other furniture|Accidental fall from other furniture
C0375736|T037|AB|E884.5|ICD9CM|Fall from furniture NEC|Fall from furniture NEC
C0478874|T037|AB|E884.9|ICD9CM|Fall-1 level to oth NEC|Fall-1 level to oth NEC
C0478874|T037|PT|E884.9|ICD9CM|Other accidental fall from one level to another|Other accidental fall from one level to another
C1135313|T037|PT|E885.0|ICD9CM|Fall from (nonmotorized) scooter|Fall from (nonmotorized) scooter
C1135313|T037|AB|E885.0|ICD9CM|Fall-nonmotor scooter|Fall-nonmotor scooter
C0878747|T037|AB|E885.2|ICD9CM|Fall from skateboard|Fall from skateboard
C0878747|T037|PT|E885.2|ICD9CM|Fall from skateboard|Fall from skateboard
C0878749|T037|AB|E885.4|ICD9CM|Fall from snowboard|Fall from snowboard
C0878749|T037|PT|E885.4|ICD9CM|Fall from snowboard|Fall from snowboard
C0261618|T037|AB|E886.9|ICD9CM|Fall on level NEC/NOS|Fall on level NEC/NOS
C0016658|T037|AB|E887|ICD9CM|Fracture, cause NOS|Fracture, cause NOS
C0016658|T037|PT|E887|ICD9CM|Fracture, cause unspecified|Fracture, cause unspecified
C0949159|T033|PT|E888.0|ICD9CM|Fall resulting in striking against sharp object|Fall resulting in striking against sharp object
C0949159|T033|AB|E888.0|ICD9CM|Fall striking sharp obj|Fall striking sharp obj
C0949160|T033|PT|E888.1|ICD9CM|Fall resulting in striking against other object|Fall resulting in striking against other object
C0949160|T033|AB|E888.1|ICD9CM|Fall striking object NEC|Fall striking object NEC
C0416980|T037|AB|E888.8|ICD9CM|Fall NEC|Fall NEC
C0416980|T037|PT|E888.8|ICD9CM|Other fall|Other fall
C0085639|T033|AB|E888.9|ICD9CM|Fall NOS|Fall NOS
C0085639|T033|PT|E888.9|ICD9CM|Unspecified fall|Unspecified fall
C0261620|T037|HT|E890|ICD9CM|Conflagration in private dwelling|Conflagration in private dwelling
C0417090|T037|AB|E891.8|ICD9CM|Fire in bldg-accid NEC|Fire in bldg-accid NEC
C0417090|T037|PT|E891.8|ICD9CM|Other accident resulting from conflagration in other and unspecified building or structure|Other accident resulting from conflagration in other and unspecified building or structure
C0417413|T037|PT|E893.9|ICD9CM|Accident caused by ignition of clothing by unspecified source|Accident caused by ignition of clothing by unspecified source
C0417413|T037|AB|E893.9|ICD9CM|Clothing fire NOS|Clothing fire NOS
C0261642|T037|PT|E895|ICD9CM|Accident caused by controlled fire in private dwelling|Accident caused by controlled fire in private dwelling
C0261642|T037|AB|E895|ICD9CM|Burn acc in privat dwell|Burn acc in privat dwell
C0417496|T037|PT|E898.0|ICD9CM|Accident caused by burning bedclothes|Accident caused by burning bedclothes
C0417496|T037|AB|E898.0|ICD9CM|Burning bedclothes|Burning bedclothes
C0261648|T037|HT|E900|ICD9CM|Accident caused by excessive heat|Accident caused by excessive heat
C0178357|T037|HT|E900-E909.9|ICD9CM|ACCIDENTS DUE TO NATURAL AND ENVIRONMENTAL FACTORS|ACCIDENTS DUE TO NATURAL AND ENVIRONMENTAL FACTORS
C0000909|T037|PT|E900.0|ICD9CM|Accident caused by excessive heat due to weather conditions|Accident caused by excessive heat due to weather conditions
C0000909|T037|AB|E900.0|ICD9CM|Excessive heat: weather|Excessive heat: weather
C0000926|T037|PT|E900.9|ICD9CM|Accidents due to excessive heat of unspecified origin|Accidents due to excessive heat of unspecified origin
C0000926|T037|AB|E900.9|ICD9CM|Excessive heat NOS|Excessive heat NOS
C0261650|T037|HT|E901|ICD9CM|Accidents due to excessive cold|Accidents due to excessive cold
C0161734|T037|PT|E901.9|ICD9CM|Accident due to excessive cold of unspecified origin|Accident due to excessive cold of unspecified origin
C0161734|T037|AB|E901.9|ICD9CM|Excessive cold NOS|Excessive cold NOS
C0000916|T037|PT|E902.0|ICD9CM|Accident due to residence or prolonged visit at high altitude|Accident due to residence or prolonged visit at high altitude
C0000916|T037|AB|E902.0|ICD9CM|High altitude residence|High altitude residence
C0000914|T037|PT|E902.2|ICD9CM|Accident due to changes in air pressure due to diving|Accident due to changes in air pressure due to diving
C0000914|T037|AB|E902.2|ICD9CM|Air press change: diving|Air press change: diving
C0480147|T037|PT|E903|ICD9CM|Accident caused by travel and motion|Accident caused by travel and motion
C0480147|T037|AB|E903|ICD9CM|Travel and motion|Travel and motion
C0417672|T037|PT|E904.1|ICD9CM|Accident due to lack of food|Accident due to lack of food
C0417672|T037|AB|E904.1|ICD9CM|Lack of food|Lack of food
C0417673|T033|PT|E904.2|ICD9CM|Accident due to lack of water|Accident due to lack of water
C0417673|T033|AB|E904.2|ICD9CM|Lack of water|Lack of water
C0546841|T037|PT|E904.3|ICD9CM|Accident due to exposure (to weather conditions), not elsewhere classifiable|Accident due to exposure (to weather conditions), not elsewhere classifiable
C0546841|T037|AB|E904.3|ICD9CM|Exposure NEC|Exposure NEC
C0417584|T037|PT|E904.9|ICD9CM|Accident due to privation, unqualified|Accident due to privation, unqualified
C0417584|T037|AB|E904.9|ICD9CM|Privation NOS|Privation NOS
C0261662|T037|HT|E905|ICD9CM|Venomous animals and plants as the cause of poisoning and toxic reactions|Venomous animals and plants as the cause of poisoning and toxic reactions
C0042477|T037|AB|E905.0|ICD9CM|Venomous snake bite|Venomous snake bite
C0042477|T037|PT|E905.0|ICD9CM|Venomous snakes and lizards causing poisoning and toxic reactions|Venomous snakes and lizards causing poisoning and toxic reactions
C0042478|T037|AB|E905.1|ICD9CM|Venomous spider bite|Venomous spider bite
C0042478|T037|PT|E905.1|ICD9CM|Venomous spiders causing poisoning and toxic reactions|Venomous spiders causing poisoning and toxic reactions
C0261663|T037|AB|E905.2|ICD9CM|Scorpion sting|Scorpion sting
C0261663|T037|PT|E905.2|ICD9CM|Scorpion sting causing poisoning and toxic reactions|Scorpion sting causing poisoning and toxic reactions
C0261664|T037|AB|E905.3|ICD9CM|Hornet/wasp/bee sting|Hornet/wasp/bee sting
C0261664|T037|PT|E905.3|ICD9CM|Sting of hornets, wasps, and bees causing poisoning and toxic reactions|Sting of hornets, wasps, and bees causing poisoning and toxic reactions
C0261665|T037|PT|E905.4|ICD9CM|Centipede and venomous millipede (tropical) bite causing poisoning and toxic reactions|Centipede and venomous millipede (tropical) bite causing poisoning and toxic reactions
C0261665|T037|AB|E905.4|ICD9CM|Centipede bite|Centipede bite
C0261666|T037|PT|E905.5|ICD9CM|Other venomous arthropods causing poisoning and toxic reactions|Other venomous arthropods causing poisoning and toxic reactions
C0261666|T037|AB|E905.5|ICD9CM|Venomous arthropods NEC|Venomous arthropods NEC
C0261667|T037|AB|E905.6|ICD9CM|Venom sea animals/plants|Venom sea animals/plants
C0261667|T037|PT|E905.6|ICD9CM|Venomous marine animals and plants causing poisoning and toxic reactions|Venomous marine animals and plants causing poisoning and toxic reactions
C0261668|T037|PT|E905.7|ICD9CM|Poisoning and toxic reactions caused by other plants|Poisoning and toxic reactions caused by other plants
C0261668|T037|AB|E905.7|ICD9CM|Poisoning by other plant|Poisoning by other plant
C0261669|T037|PT|E905.8|ICD9CM|Poisoning and toxic reactions caused by other specified animals and plants|Poisoning and toxic reactions caused by other specified animals and plants
C0261669|T037|AB|E905.8|ICD9CM|Venomous bite/sting NEC|Venomous bite/sting NEC
C0261670|T037|PT|E905.9|ICD9CM|Poisoning and toxic reactions caused by unspecified animals and plants|Poisoning and toxic reactions caused by unspecified animals and plants
C0261670|T037|AB|E905.9|ICD9CM|Venomous bite/sting NOS|Venomous bite/sting NOS
C0417758|T037|HT|E906|ICD9CM|Other injury caused by animals|Other injury caused by animals
C0259797|T037|AB|E906.0|ICD9CM|Dog bite|Dog bite
C0259797|T037|PT|E906.0|ICD9CM|Dog bite|Dog bite
C0479196|T037|AB|E906.1|ICD9CM|Rat bite|Rat bite
C0479196|T037|PT|E906.1|ICD9CM|Rat bite|Rat bite
C0546830|T037|PT|E906.2|ICD9CM|Bite of nonvenomous snakes and lizards|Bite of nonvenomous snakes and lizards
C0546830|T037|AB|E906.2|ICD9CM|Nonvenomous snake bite|Nonvenomous snake bite
C0005656|T037|AB|E906.3|ICD9CM|Animal bite NEC|Animal bite NEC
C0005656|T037|PT|E906.3|ICD9CM|Bite of other animal except arthropod|Bite of other animal except arthropod
C0332815|T037|PT|E906.4|ICD9CM|Bite of nonvenomous arthropod|Bite of nonvenomous arthropod
C0332815|T037|AB|E906.4|ICD9CM|Nonvenom arthropod bite|Nonvenom arthropod bite
C0003044|T037|AB|E906.5|ICD9CM|Animal bite NOS|Animal bite NOS
C0003044|T037|PT|E906.5|ICD9CM|Bite by unspecified animal|Bite by unspecified animal
C0261675|T037|AB|E906.9|ICD9CM|Inj NOS caused by animal|Inj NOS caused by animal
C0261675|T037|PT|E906.9|ICD9CM|Unspecified injury caused by animal|Unspecified injury caused by animal
C0000915|T037|AB|E907|ICD9CM|Acc due to lightning|Acc due to lightning
C0000915|T037|PT|E907|ICD9CM|Accident due to lightning|Accident due to lightning
C0375739|T037|AB|E908.0|ICD9CM|Accident d/t hurricane|Accident d/t hurricane
C0375739|T037|PT|E908.0|ICD9CM|Hurricane|Hurricane
C0375740|T037|AB|E908.1|ICD9CM|Accident d/t tornado|Accident d/t tornado
C0375740|T037|PT|E908.1|ICD9CM|Tornado|Tornado
C0375741|T037|AB|E908.2|ICD9CM|Accident d/t floods|Accident d/t floods
C0375741|T037|PT|E908.2|ICD9CM|Floods|Floods
C0375742|T037|AB|E908.3|ICD9CM|Acc d/t snow blizzard|Acc d/t snow blizzard
C0375742|T037|PT|E908.3|ICD9CM|Blizzard (snow) (ice)|Blizzard (snow) (ice)
C0375743|T037|AB|E908.4|ICD9CM|Accident d/t dust storm|Accident d/t dust storm
C0375743|T037|PT|E908.4|ICD9CM|Dust storm|Dust storm
C0375744|T037|AB|E908.8|ICD9CM|Accident d/t storm NEC|Accident d/t storm NEC
C0375744|T037|PT|E908.8|ICD9CM|Other cataclysmic storms|Other cataclysmic storms
C0417614|T037|AB|E909.0|ICD9CM|Acc d/t earthquakes|Acc d/t earthquakes
C0417614|T037|PT|E909.0|ICD9CM|Earthquakes|Earthquakes
C0375746|T037|AB|E909.1|ICD9CM|Acc d/t volcanic erupt|Acc d/t volcanic erupt
C0375746|T037|PT|E909.1|ICD9CM|Volcanic eruptions|Volcanic eruptions
C0375747|T037|AB|E909.2|ICD9CM|Acc d/t avalanche|Acc d/t avalanche
C0375747|T037|PT|E909.2|ICD9CM|Avalanche, landslide, or mudslide|Avalanche, landslide, or mudslide
C0261678|T037|HT|E910|ICD9CM|Accidental drowning and submersion|Accidental drowning and submersion
C0261679|T037|PT|E910.0|ICD9CM|Accidental drowning and submersion while water-skiing|Accidental drowning and submersion while water-skiing
C0261679|T037|AB|E910.0|ICD9CM|Water-skiing accident|Water-skiing accident
C0417794|T037|AB|E910.1|ICD9CM|Skin/scuba diving acc|Skin/scuba diving acc
C0261681|T037|AB|E910.2|ICD9CM|Swimming accident NOS|Swimming accident NOS
C0261683|T037|PT|E910.4|ICD9CM|Accidental drowning and submersion in bathtub|Accidental drowning and submersion in bathtub
C0261683|T037|AB|E910.4|ICD9CM|Drowning in bathtub|Drowning in bathtub
C0029483|T037|AB|E910.8|ICD9CM|Accidental drowning NEC|Accidental drowning NEC
C0029483|T037|PT|E910.8|ICD9CM|Other accidental drowning or submersion|Other accidental drowning or submersion
C0261684|T037|AB|E910.9|ICD9CM|Accidental drowning NOS|Accidental drowning NOS
C0261684|T037|PT|E910.9|ICD9CM|Unspecified accidental drowning or submersion|Unspecified accidental drowning or submersion
C0261685|T037|PT|E911|ICD9CM|Inhalation and ingestion of food causing obstruction of respiratory tract or suffocation|Inhalation and ingestion of food causing obstruction of respiratory tract or suffocation
C0261685|T037|AB|E911|ICD9CM|Resp obstr-food inhal|Resp obstr-food inhal
C0261686|T037|PT|E912|ICD9CM|Inhalation and ingestion of other object causing obstruction of respiratory tract or suffocation|Inhalation and ingestion of other object causing obstruction of respiratory tract or suffocation
C0261686|T037|AB|E912|ICD9CM|Resp obstr-inhal obj NEC|Resp obstr-inhal obj NEC
C0559051|T037|HT|E913|ICD9CM|Accidental mechanical suffocation|Accidental mechanical suffocation
C0261688|T037|PT|E913.0|ICD9CM|Accidental mechanical suffocation in bed or cradle|Accidental mechanical suffocation in bed or cradle
C0261688|T037|AB|E913.0|ICD9CM|Suffocat in bed/cradle|Suffocat in bed/cradle
C0261689|T037|PT|E913.1|ICD9CM|Accidental mechanical suffocation by plastic bag|Accidental mechanical suffocation by plastic bag
C0261689|T037|AB|E913.1|ICD9CM|Suffocation-plastic bag|Suffocation-plastic bag
C0261690|T037|PT|E913.2|ICD9CM|Accidental mechanical suffocation due to lack of air (in closed place)|Accidental mechanical suffocation due to lack of air (in closed place)
C0261690|T037|AB|E913.2|ICD9CM|Suffocation-lack of air|Suffocation-lack of air
C0261691|T037|PT|E913.3|ICD9CM|Accidental mechanical suffocation by falling earth or other substance|Accidental mechanical suffocation by falling earth or other substance
C0261691|T037|AB|E913.3|ICD9CM|Cave-in NOS|Cave-in NOS
C0261692|T037|PT|E913.8|ICD9CM|Accidental mechanical suffocation by other specified means|Accidental mechanical suffocation by other specified means
C0261692|T037|AB|E913.8|ICD9CM|Suffocation NEC|Suffocation NEC
C0000922|T037|PT|E913.9|ICD9CM|Accidental mechanical suffocation by unspecified means|Accidental mechanical suffocation by unspecified means
C0000922|T037|AB|E913.9|ICD9CM|Suffocation NOS|Suffocation NOS
C0261693|T037|AB|E914|ICD9CM|FB entering eye|FB entering eye
C0261693|T037|PT|E914|ICD9CM|Foreign body accidentally entering eye and adnexa|Foreign body accidentally entering eye and adnexa
C0261694|T037|AB|E915|ICD9CM|FB entering oth orifice|FB entering oth orifice
C0261694|T037|PT|E915|ICD9CM|Foreign body accidentally entering other orifice|Foreign body accidentally entering other orifice
C0261695|T037|PT|E916|ICD9CM|Struck accidentally by falling object|Struck accidentally by falling object
C0261695|T037|AB|E916|ICD9CM|Struck by falling object|Struck by falling object
C0029484|T037|HT|E916-E928.9|ICD9CM|OTHER ACCIDENTS|OTHER ACCIDENTS
C0949169|T037|AB|E917.0|ICD9CM|Sports acc w/o sub fall|Sports acc w/o sub fall
C0949169|T037|PT|E917.0|ICD9CM|Striking against or struck accidentally by objects or persons in sports|Striking against or struck accidentally by objects or persons in sports
C0949170|T037|AB|E917.1|ICD9CM|Crowd w/o sub fall|Crowd w/o sub fall
C0949170|T037|PT|E917.1|ICD9CM|Striking against or struck accidentally by a crowd, by collective fear or panic|Striking against or struck accidentally by a crowd, by collective fear or panic
C0949171|T037|AB|E917.2|ICD9CM|Run water w/o sub fall|Run water w/o sub fall
C0949171|T037|PT|E917.2|ICD9CM|Striking against or struck accidentally in running water|Striking against or struck accidentally in running water
C0949161|T037|AB|E917.3|ICD9CM|Furnit w/o sub fall|Furnit w/o sub fall
C0949161|T037|PT|E917.3|ICD9CM|Striking against or struck accidentally by furniture without subsequent fall|Striking against or struck accidentally by furniture without subsequent fall
C0949162|T037|AB|E917.4|ICD9CM|Stat ob w/o sub fall NEC|Stat ob w/o sub fall NEC
C0949162|T037|PT|E917.4|ICD9CM|Striking against or struck accidentally by other stationary object without subsequent fall|Striking against or struck accidentally by other stationary object without subsequent fall
C0949163|T037|AB|E917.5|ICD9CM|Sports acc w sub fall|Sports acc w sub fall
C0949163|T037|PT|E917.5|ICD9CM|Striking against or struck accidentally by object in sports with subsequent fall|Striking against or struck accidentally by object in sports with subsequent fall
C0949164|T037|AB|E917.6|ICD9CM|Crowd accidnt w sub fall|Crowd accidnt w sub fall
C0949165|T037|AB|E917.7|ICD9CM|Furniture acc w sub fall|Furniture acc w sub fall
C0949165|T037|PT|E917.7|ICD9CM|Striking against or struck accidentally by furniture with subsequent fall|Striking against or struck accidentally by furniture with subsequent fall
C0949166|T037|AB|E917.8|ICD9CM|Stat obj w sub fall NEC|Stat obj w sub fall NEC
C0949166|T037|PT|E917.8|ICD9CM|Striking against or struck accidentally by other stationary object with subsequent fall|Striking against or struck accidentally by other stationary object with subsequent fall
C0949172|T037|AB|E917.9|ICD9CM|Obj w-w/o sub fall NEC|Obj w-w/o sub fall NEC
C0949172|T037|PT|E917.9|ICD9CM|Other accident caused by striking against or being struck accidentally by objects or persons|Other accident caused by striking against or being struck accidentally by objects or persons
C1278558|T037|PT|E918|ICD9CM|Caught accidentally in or between objects|Caught accidentally in or between objects
C1278558|T037|AB|E918|ICD9CM|Caught between objects|Caught between objects
C0261712|T037|HT|E919|ICD9CM|Accidents caused by machinery|Accidents caused by machinery
C0261703|T037|PT|E919.0|ICD9CM|Accidents caused by agricultural machines|Accidents caused by agricultural machines
C0261703|T037|AB|E919.0|ICD9CM|Machine accid-agricult|Machine accid-agricult
C0261704|T037|PT|E919.1|ICD9CM|Accidents caused by mining and earth-drilling machinery|Accidents caused by mining and earth-drilling machinery
C0261704|T037|AB|E919.1|ICD9CM|Machine accid-mining|Machine accid-mining
C0261706|T037|PT|E919.3|ICD9CM|Accidents caused by metalworking machines|Accidents caused by metalworking machines
C0261706|T037|AB|E919.3|ICD9CM|Metalworking machine acc|Metalworking machine acc
C0261708|T037|PT|E919.5|ICD9CM|Accidents caused by prime movers, except electrical motors|Accidents caused by prime movers, except electrical motors
C0261708|T037|AB|E919.5|ICD9CM|Prime mover machine acc|Prime mover machine acc
C0261709|T037|PT|E919.6|ICD9CM|Accidents caused by transmission machinery|Accidents caused by transmission machinery
C0261709|T037|AB|E919.6|ICD9CM|Transmission machine acc|Transmission machine acc
C0261710|T037|PT|E919.7|ICD9CM|Accidents caused by earth moving, scraping, and other excavating machines|Accidents caused by earth moving, scraping, and other excavating machines
C0261710|T037|AB|E919.7|ICD9CM|Earth moving machine acc|Earth moving machine acc
C0261711|T037|PT|E919.8|ICD9CM|Accidents caused by other specified machinery|Accidents caused by other specified machinery
C0261711|T037|AB|E919.8|ICD9CM|Machinery accident NEC|Machinery accident NEC
C0261712|T037|PT|E919.9|ICD9CM|Accidents caused by unspecified machinery|Accidents caused by unspecified machinery
C0261712|T037|AB|E919.9|ICD9CM|Machinery accident NOS|Machinery accident NOS
C0261713|T037|HT|E920|ICD9CM|Accidents caused by cutting and piercing instruments or objects|Accidents caused by cutting and piercing instruments or objects
C0261714|T037|AB|E920.0|ICD9CM|Acc-powered lawn mower|Acc-powered lawn mower
C0261714|T037|PT|E920.0|ICD9CM|Accidents caused by powered lawn mower|Accidents caused by powered lawn mower
C0261715|T037|AB|E920.1|ICD9CM|Acc-power hand tool NEC|Acc-power hand tool NEC
C0261715|T037|PT|E920.1|ICD9CM|Accidents caused by other powered hand tools|Accidents caused by other powered hand tools
C0261716|T037|AB|E920.2|ICD9CM|Acc-power house applianc|Acc-power house applianc
C0261716|T037|PT|E920.2|ICD9CM|Accidents caused by powered household appliances and implements|Accidents caused by powered household appliances and implements
C0261717|T037|PT|E920.3|ICD9CM|Accidents caused by knives, swords, and daggers|Accidents caused by knives, swords, and daggers
C0261717|T037|AB|E920.3|ICD9CM|Knife/sword/dagger acc|Knife/sword/dagger acc
C0261718|T037|AB|E920.4|ICD9CM|Accid-other hand tools|Accid-other hand tools
C0261718|T037|PT|E920.4|ICD9CM|Accidents caused by other hand tools and implements|Accidents caused by other hand tools and implements
C0375752|T037|AB|E920.5|ICD9CM|Acc-hypodermic needle|Acc-hypodermic needle
C0375752|T037|PT|E920.5|ICD9CM|Accidents caused by hypodermic needle|Accidents caused by hypodermic needle
C0261719|T037|AB|E920.8|ICD9CM|Acc-cutting instrum NEC|Acc-cutting instrum NEC
C0261719|T037|PT|E920.8|ICD9CM|Accidents caused by other specified cutting and piercing instruments or objects|Accidents caused by other specified cutting and piercing instruments or objects
C0261713|T037|AB|E920.9|ICD9CM|Acc-cutting instrum NOS|Acc-cutting instrum NOS
C0261713|T037|PT|E920.9|ICD9CM|Accidents caused by unspecified cutting and piercing instrument or object|Accidents caused by unspecified cutting and piercing instrument or object
C0261724|T037|HT|E921|ICD9CM|Accident caused by explosion of pressure vessel|Accident caused by explosion of pressure vessel
C0261721|T037|PT|E921.0|ICD9CM|Accident caused by explosion of boilers|Accident caused by explosion of boilers
C0261721|T037|AB|E921.0|ICD9CM|Boiler explosion|Boiler explosion
C0261722|T037|PT|E921.1|ICD9CM|Accident caused by explosion of gas cylinders|Accident caused by explosion of gas cylinders
C0261722|T037|AB|E921.1|ICD9CM|Gas cylinder explosion|Gas cylinder explosion
C0261724|T037|PT|E921.9|ICD9CM|Accident caused by explosion of unspecified pressure vessel|Accident caused by explosion of unspecified pressure vessel
C0261724|T037|AB|E921.9|ICD9CM|Press vessel explos NOS|Press vessel explos NOS
C0490042|T037|HT|E922|ICD9CM|Accident caused by firearm, and air gun missile|Accident caused by firearm, and air gun missile
C0261726|T037|PT|E922.0|ICD9CM|Accident caused by handgun|Accident caused by handgun
C0261726|T037|AB|E922.0|ICD9CM|Handgun accident|Handgun accident
C0565898|T037|PT|E922.1|ICD9CM|Accident caused by shotgun (automatic)|Accident caused by shotgun (automatic)
C0565898|T037|AB|E922.1|ICD9CM|Shotgun accident|Shotgun accident
C0261728|T037|PT|E922.2|ICD9CM|Accident caused by hunting rifle|Accident caused by hunting rifle
C0261728|T037|AB|E922.2|ICD9CM|Hunting rifle accident|Hunting rifle accident
C0261729|T037|PT|E922.3|ICD9CM|Accident caused by military firearms|Accident caused by military firearms
C0261729|T037|AB|E922.3|ICD9CM|Military firearm accid|Military firearm accid
C0490035|T037|AB|E922.4|ICD9CM|Accident - air gun|Accident - air gun
C0490035|T037|PT|E922.4|ICD9CM|Accident caused by air gun|Accident caused by air gun
C1135314|T037|PT|E922.5|ICD9CM|Accident caused by paintball gun|Accident caused by paintball gun
C1135314|T037|AB|E922.5|ICD9CM|Accident-paintball gun|Accident-paintball gun
C0261725|T037|PT|E922.9|ICD9CM|Accident caused by unspecified firearm missile|Accident caused by unspecified firearm missile
C0261725|T037|AB|E922.9|ICD9CM|Firearm accident NOS|Firearm accident NOS
C0261731|T037|HT|E923|ICD9CM|Accident caused by explosive material|Accident caused by explosive material
C0261732|T037|PT|E923.0|ICD9CM|Accident caused by fireworks|Accident caused by fireworks
C0261732|T037|AB|E923.0|ICD9CM|Fireworks accident|Fireworks accident
C0261733|T037|PT|E923.1|ICD9CM|Accident caused by blasting materials|Accident caused by blasting materials
C0261733|T037|AB|E923.1|ICD9CM|Blasting materials accid|Blasting materials accid
C0261734|T037|PT|E923.2|ICD9CM|Accident caused by explosive gases|Accident caused by explosive gases
C0261734|T037|AB|E923.2|ICD9CM|Explosive gases accident|Explosive gases accident
C0261735|T037|PT|E923.8|ICD9CM|Accident caused by other explosive materials|Accident caused by other explosive materials
C0261735|T037|AB|E923.8|ICD9CM|Explosives accident NEC|Explosives accident NEC
C0261731|T037|PT|E923.9|ICD9CM|Accident caused by unspecified explosive material|Accident caused by unspecified explosive material
C0261731|T037|AB|E923.9|ICD9CM|Explosives accident NOS|Explosives accident NOS
C0261736|T037|HT|E924|ICD9CM|Accident caused by hot substance or object, caustic or corrosive material, and steam|Accident caused by hot substance or object, caustic or corrosive material, and steam
C0261737|T037|AB|E924.0|ICD9CM|Acc-hot liquid & steam|Acc-hot liquid & steam
C0261737|T037|PT|E924.0|ICD9CM|Accident caused by hot liquids and vapors, including steam|Accident caused by hot liquids and vapors, including steam
C0000908|T037|AB|E924.1|ICD9CM|Accid-caustic substance|Accid-caustic substance
C0000908|T037|PT|E924.1|ICD9CM|Accident caused by caustic and corrosive substances|Accident caused by caustic and corrosive substances
C0375753|T037|AB|E924.2|ICD9CM|Acc-hot tap water|Acc-hot tap water
C0375753|T037|PT|E924.2|ICD9CM|Accident caused by hot (boiling) tap water|Accident caused by hot (boiling) tap water
C0261738|T037|PT|E924.8|ICD9CM|Accident caused by other hot substance or object|Accident caused by other hot substance or object
C0261738|T037|AB|E924.8|ICD9CM|Hot substance accid NEC|Hot substance accid NEC
C0261740|T037|HT|E925|ICD9CM|Accident caused by electric current|Accident caused by electric current
C0261744|T037|PT|E925.8|ICD9CM|Accident caused by other electric current|Accident caused by other electric current
C0261744|T037|AB|E925.8|ICD9CM|Electric current acc NEC|Electric current acc NEC
C0261740|T037|PT|E925.9|ICD9CM|Accident caused by unspecified electric current|Accident caused by unspecified electric current
C0261740|T037|AB|E925.9|ICD9CM|Electric current acc NOS|Electric current acc NOS
C0015333|T037|HT|E926|ICD9CM|Exposure to radiation|Exposure to radiation
C0261746|T037|PT|E926.0|ICD9CM|Exposure to radiofrequency radiation|Exposure to radiofrequency radiation
C0261746|T037|AB|E926.0|ICD9CM|Radiofreq radiat exposur|Radiofreq radiat exposur
C0261747|T037|PT|E926.1|ICD9CM|Exposure to infra-red radiation from heaters and lamps|Exposure to infra-red radiation from heaters and lamps
C0261747|T037|AB|E926.1|ICD9CM|Infra-red appl rad exos|Infra-red appl rad exos
C0015335|T037|PT|E926.2|ICD9CM|Exposure to visible and ultraviolet light sources|Exposure to visible and ultraviolet light sources
C0015335|T037|AB|E926.2|ICD9CM|Vis/ultraviol lght expos|Vis/ultraviol lght expos
C0261748|T037|PT|E926.3|ICD9CM|Exposure to x-rays and other electromagnetic ionizing radiation|Exposure to x-rays and other electromagnetic ionizing radiation
C0261748|T037|AB|E926.3|ICD9CM|X-ray/gamma ray exposure|X-ray/gamma ray exposure
C0261749|T037|PT|E926.4|ICD9CM|Exposure to lasers|Exposure to lasers
C0261749|T037|AB|E926.4|ICD9CM|Laser exposure|Laser exposure
C0261750|T037|PT|E926.5|ICD9CM|Exposure to radioactive isotopes|Exposure to radioactive isotopes
C0261750|T037|AB|E926.5|ICD9CM|Radioact isotope exposur|Radioact isotope exposur
C0015332|T037|PT|E926.8|ICD9CM|Exposure to other specified radiation|Exposure to other specified radiation
C0015332|T037|AB|E926.8|ICD9CM|Radiation exposure NEC|Radiation exposure NEC
C0015333|T037|PT|E926.9|ICD9CM|Exposure to unspecified radiation|Exposure to unspecified radiation
C0015333|T037|AB|E926.9|ICD9CM|Radiation exposure NOS|Radiation exposure NOS
C2349815|T033|HT|E927|ICD9CM|Overexertion and strenuous and repetitive movements or loads|Overexertion and strenuous and repetitive movements or loads
C2349803|T047|PT|E927.0|ICD9CM|Overexertion from sudden strenuous movement|Overexertion from sudden strenuous movement
C2349803|T047|AB|E927.0|ICD9CM|Overxrt-sudn stren mvmt|Overxrt-sudn stren mvmt
C2349805|T047|PT|E927.1|ICD9CM|Overexertion from prolonged static position|Overexertion from prolonged static position
C2349805|T047|AB|E927.1|ICD9CM|Overxrt-prolng stc postn|Overxrt-prolng stc postn
C2349809|T037|AB|E927.2|ICD9CM|Excess physical exert|Excess physical exert
C2349809|T037|PT|E927.2|ICD9CM|Excessive physical exertion|Excessive physical exertion
C2349810|T037|AB|E927.3|ICD9CM|Cumltv trma-repetv motn|Cumltv trma-repetv motn
C2349810|T037|PT|E927.3|ICD9CM|Cumulative trauma from repetitive motion|Cumulative trauma from repetitive motion
C2349812|T037|AB|E927.4|ICD9CM|Cumltv trma-repetv impct|Cumltv trma-repetv impct
C2349812|T037|PT|E927.4|ICD9CM|Cumulative trauma from repetitive impact|Cumulative trauma from repetitive impact
C2349813|T047|PT|E927.8|ICD9CM|Other overexertion and strenuous and repetitive movements or loads|Other overexertion and strenuous and repetitive movements or loads
C2349813|T047|AB|E927.8|ICD9CM|Overexert reptv mvmt NEC|Overexert reptv mvmt NEC
C2349814|T047|AB|E927.9|ICD9CM|Overexert reptv mvmt NOS|Overexert reptv mvmt NOS
C2349814|T047|PT|E927.9|ICD9CM|Unspecified overexertion and strenuous and repetitive movements or loads|Unspecified overexertion and strenuous and repetitive movements or loads
C0261752|T037|AB|E928.0|ICD9CM|Acc d/t weightless envir|Acc d/t weightless envir
C0261752|T037|PT|E928.0|ICD9CM|Prolonged stay in weightless environment|Prolonged stay in weightless environment
C0700522|T037|AB|E928.1|ICD9CM|Exposure to noise|Exposure to noise
C0700522|T037|PT|E928.1|ICD9CM|Exposure to noise|Exposure to noise
C0677519|T037|AB|E928.2|ICD9CM|Exposure to vibration|Exposure to vibration
C0677519|T037|PT|E928.2|ICD9CM|Vibration|Vibration
C0005660|T037|PT|E928.3|ICD9CM|Human bite|Human bite
C0005660|T037|AB|E928.3|ICD9CM|Human bite - accidental|Human bite - accidental
C1260473|T037|AB|E928.4|ICD9CM|Ext constriction-hair|Ext constriction-hair
C1260473|T037|PT|E928.4|ICD9CM|External constriction caused by hair|External constriction caused by hair
C1260474|T037|AB|E928.5|ICD9CM|Ext constriction-obj NEC|Ext constriction-obj NEC
C1260474|T037|PT|E928.5|ICD9CM|External constriction caused by other object|External constriction caused by other object
C1955556|T047|AB|E928.6|ICD9CM|Envir expose algae/toxin|Envir expose algae/toxin
C1955556|T047|PT|E928.6|ICD9CM|Environmental exposure to harmful algae and toxins|Environmental exposure to harmful algae and toxins
C2712481|T037|AB|E928.7|ICD9CM|Accidnt-mech firearm/gun|Accidnt-mech firearm/gun
C2712481|T037|PT|E928.7|ICD9CM|Environmental and accidental causes, mechanism or component of firearm and air gun|Environmental and accidental causes, mechanism or component of firearm and air gun
C0029484|T037|AB|E928.8|ICD9CM|Accident NEC|Accident NEC
C0029484|T037|PT|E928.8|ICD9CM|Other accidents|Other accidents
C4759661|T037|AB|E928.9|ICD9CM|Accident NOS|Accident NOS
C4759661|T037|PT|E928.9|ICD9CM|Unspecified accident|Unspecified accident
C0176005|T033|HT|E929|ICD9CM|Late effects of accidental injury|Late effects of accidental injury
C0176005|T033|HT|E929-E929.9|ICD9CM|LATE EFFECTS OF ACCIDENTAL INJURY|LATE EFFECTS OF ACCIDENTAL INJURY
C0481354|T037|AB|E929.0|ICD9CM|Late eff motor vehic acc|Late eff motor vehic acc
C0481354|T037|PT|E929.0|ICD9CM|Late effects of motor vehicle accident|Late effects of motor vehicle accident
C0481355|T037|AB|E929.1|ICD9CM|Late eff transport acc|Late eff transport acc
C0481355|T037|PT|E929.1|ICD9CM|Late effects of other transport accident|Late effects of other transport accident
C0261755|T046|AB|E929.2|ICD9CM|Late eff acc poisoning|Late eff acc poisoning
C0261755|T046|PT|E929.2|ICD9CM|Late effects of accidental poisoning|Late effects of accidental poisoning
C0261756|T046|AB|E929.3|ICD9CM|Late eff accidental fall|Late eff accidental fall
C0261756|T046|PT|E929.3|ICD9CM|Late effects of accidental fall|Late effects of accidental fall
C0261757|T046|AB|E929.4|ICD9CM|Late eff fire acc|Late eff fire acc
C0261757|T046|PT|E929.4|ICD9CM|Late effects of accident caused by fire|Late effects of accident caused by fire
C0261758|T046|AB|E929.5|ICD9CM|Late eff environment acc|Late eff environment acc
C0261758|T046|PT|E929.5|ICD9CM|Late effects of accident due to natural and environmental factors|Late effects of accident due to natural and environmental factors
C2733645|T046|AB|E929.8|ICD9CM|Late eff accident NEC|Late eff accident NEC
C2733645|T046|PT|E929.8|ICD9CM|Late effects of other accidents|Late effects of other accidents
C0274271|T046|AB|E929.9|ICD9CM|Late eff accident NOS|Late eff accident NOS
C0274271|T046|PT|E929.9|ICD9CM|Late effects of unspecified accident|Late effects of unspecified accident
C0261771|T037|HT|E930|ICD9CM|Antibiotics causing adverse effects in therapeutic use|Antibiotics causing adverse effects in therapeutic use
C0178359|T046|HT|E930-E949.9|ICD9CM|DRUGS, MEDICINAL AND BIOLOGICAL SUBSTANCES CAUSING ADVERSE EFFECTS IN THERAPEUTIC USE|DRUGS, MEDICINAL AND BIOLOGICAL SUBSTANCES CAUSING ADVERSE EFFECTS IN THERAPEUTIC USE
C0413443|T046|AB|E930.0|ICD9CM|Adv eff penicillins|Adv eff penicillins
C0413443|T046|PT|E930.0|ICD9CM|Penicillins causing adverse effects in therapeutic use|Penicillins causing adverse effects in therapeutic use
C0481115|T037|AB|E930.1|ICD9CM|Adv eff antifung antbiot|Adv eff antifung antbiot
C0481115|T037|PT|E930.1|ICD9CM|Antifungal antibiotics causing adverse effects in therapeutic use|Antifungal antibiotics causing adverse effects in therapeutic use
C0851330|T037|AB|E930.2|ICD9CM|Adv eff chloramphenicol|Adv eff chloramphenicol
C0851330|T037|PT|E930.2|ICD9CM|Chloramphenicol group causing adverse effects in therapeutic use|Chloramphenicol group causing adverse effects in therapeutic use
C0261765|T037|AB|E930.3|ICD9CM|Adv eff erythromycin|Adv eff erythromycin
C0261765|T037|PT|E930.3|ICD9CM|Erythromycin and other macrolides causing adverse effects in therapeutic use|Erythromycin and other macrolides causing adverse effects in therapeutic use
C0261766|T037|AB|E930.4|ICD9CM|Adv eff tetracycline|Adv eff tetracycline
C0261766|T037|PT|E930.4|ICD9CM|Tetracycline group causing adverse effects in therapeutic use|Tetracycline group causing adverse effects in therapeutic use
C0261767|T037|AB|E930.5|ICD9CM|Adv eff cephalosporin|Adv eff cephalosporin
C0261767|T037|PT|E930.5|ICD9CM|Cephalosporin group causing adverse effects in therapeutic use|Cephalosporin group causing adverse effects in therapeutic use
C0261768|T037|AB|E930.6|ICD9CM|Adv eff antmycob antbiot|Adv eff antmycob antbiot
C0261768|T037|PT|E930.6|ICD9CM|Antimycobacterial antibiotics causing adverse effects in therapeutic use|Antimycobacterial antibiotics causing adverse effects in therapeutic use
C0261769|T037|AB|E930.7|ICD9CM|Adv eff antineop antbiot|Adv eff antineop antbiot
C0261769|T037|PT|E930.7|ICD9CM|Antineoplastic antibiotics causing adverse effects in therapeutic use|Antineoplastic antibiotics causing adverse effects in therapeutic use
C0261770|T037|AB|E930.8|ICD9CM|Adv eff antibiotics NEC|Adv eff antibiotics NEC
C0261770|T037|PT|E930.8|ICD9CM|Other specified antibiotics causing adverse effects in therapeutic use|Other specified antibiotics causing adverse effects in therapeutic use
C0261771|T037|AB|E930.9|ICD9CM|Adv eff antibiotic NOS|Adv eff antibiotic NOS
C0261771|T037|PT|E930.9|ICD9CM|Unspecified antibiotic causing adverse effects in therapeutic use|Unspecified antibiotic causing adverse effects in therapeutic use
C0261772|T037|HT|E931|ICD9CM|Other anti-infectives causing adverse effects in therapeutic use|Other anti-infectives causing adverse effects in therapeutic use
C0261773|T046|AB|E931.0|ICD9CM|Adv eff sulfonamides|Adv eff sulfonamides
C0261773|T046|PT|E931.0|ICD9CM|Sulfonamides causing adverse effects in therapeutic use|Sulfonamides causing adverse effects in therapeutic use
C0261774|T037|AB|E931.1|ICD9CM|Adv eff arsenic anti-inf|Adv eff arsenic anti-inf
C0261774|T037|PT|E931.1|ICD9CM|Arsenical anti-infectives causing adverse effects in therapeutic use|Arsenical anti-infectives causing adverse effects in therapeutic use
C0261775|T037|AB|E931.2|ICD9CM|Adv eff metal anti-inf|Adv eff metal anti-inf
C0261775|T037|PT|E931.2|ICD9CM|Heavy metal anti-infectives causing adverse effects in therapeutic use|Heavy metal anti-infectives causing adverse effects in therapeutic use
C0261776|T037|AB|E931.3|ICD9CM|Adv eff quinoline|Adv eff quinoline
C0261776|T037|PT|E931.3|ICD9CM|Quinoline and hydroxyquinoline derivatives causing adverse effects in therapeutic use|Quinoline and hydroxyquinoline derivatives causing adverse effects in therapeutic use
C0261777|T037|AB|E931.4|ICD9CM|Adv eff antimalarials|Adv eff antimalarials
C0261777|T037|PT|E931.4|ICD9CM|Antimalarials and drugs acting on other blood protozoa causing adverse effects in therapeutic use|Antimalarials and drugs acting on other blood protozoa causing adverse effects in therapeutic use
C0261778|T037|AB|E931.5|ICD9CM|Adv eff antprotazoal NEC|Adv eff antprotazoal NEC
C0261778|T037|PT|E931.5|ICD9CM|Other antiprotozoal drugs causing adverse effects in therapeutic use|Other antiprotozoal drugs causing adverse effects in therapeutic use
C0413512|T046|AB|E931.6|ICD9CM|Adv eff anthelmintics|Adv eff anthelmintics
C0413512|T046|PT|E931.6|ICD9CM|Anthelmintics causing adverse effects in therapeutic use|Anthelmintics causing adverse effects in therapeutic use
C0261780|T046|AB|E931.7|ICD9CM|Adv eff antiviral drugs|Adv eff antiviral drugs
C0261780|T046|PT|E931.7|ICD9CM|Antiviral drugs causing adverse effects in therapeutic use|Antiviral drugs causing adverse effects in therapeutic use
C0261781|T037|AB|E931.8|ICD9CM|Adv eff antimycobac NEC|Adv eff antimycobac NEC
C0261781|T037|PT|E931.8|ICD9CM|Other antimycobacterial drugs causing adverse effects in therapeutic use|Other antimycobacterial drugs causing adverse effects in therapeutic use
C0261782|T037|AB|E931.9|ICD9CM|Adv eff antinfct NEC/NOS|Adv eff antinfct NEC/NOS
C0261782|T037|PT|E931.9|ICD9CM|Other and unspecified anti-infectives causing adverse effects in therapeutic use|Other and unspecified anti-infectives causing adverse effects in therapeutic use
C0261783|T037|HT|E932|ICD9CM|Hormones and synthetic substitutes causing adverse effects in therapeutic use|Hormones and synthetic substitutes causing adverse effects in therapeutic use
C0261784|T037|PT|E932.0|ICD9CM|Adrenal cortical steroids causing adverse effects in therapeutic use|Adrenal cortical steroids causing adverse effects in therapeutic use
C0261784|T037|AB|E932.0|ICD9CM|Adv eff corticosteroids|Adv eff corticosteroids
C0261785|T037|AB|E932.1|ICD9CM|Adv eff androgens|Adv eff androgens
C0261785|T037|PT|E932.1|ICD9CM|Androgens and anabolic congeners causing adverse effects in therapeutic use|Androgens and anabolic congeners causing adverse effects in therapeutic use
C0261786|T037|AB|E932.2|ICD9CM|Adv eff ovarian hormones|Adv eff ovarian hormones
C0261786|T037|PT|E932.2|ICD9CM|Ovarian hormones and synthetic substitutes causing adverse effects in therapeutic use|Ovarian hormones and synthetic substitutes causing adverse effects in therapeutic use
C0261787|T037|AB|E932.3|ICD9CM|Adv eff insulin/antidiab|Adv eff insulin/antidiab
C0261787|T037|PT|E932.3|ICD9CM|Insulins and antidiabetic agents causing adverse effects in therapeutic use|Insulins and antidiabetic agents causing adverse effects in therapeutic use
C0261788|T037|AB|E932.4|ICD9CM|Adv eff ant pituitary|Adv eff ant pituitary
C0261788|T037|PT|E932.4|ICD9CM|Anterior pituitary hormones causing adverse effects in therapeutic use|Anterior pituitary hormones causing adverse effects in therapeutic use
C0261789|T037|AB|E932.5|ICD9CM|Adv eff post pituitary|Adv eff post pituitary
C0261789|T037|PT|E932.5|ICD9CM|Posterior pituitary hormones causing adverse effects in therapeutic use|Posterior pituitary hormones causing adverse effects in therapeutic use
C0261790|T037|AB|E932.6|ICD9CM|Adv eff parathyroid|Adv eff parathyroid
C0261790|T037|PT|E932.6|ICD9CM|Parathyroid and parathyroid derivatives causing adverse effects in therapeutic use|Parathyroid and parathyroid derivatives causing adverse effects in therapeutic use
C0261791|T037|AB|E932.7|ICD9CM|Adv eff thyroid & deriv|Adv eff thyroid & deriv
C0261791|T037|PT|E932.7|ICD9CM|Thyroid and thyroid derivatives causing adverse effects in therapeutic use|Thyroid and thyroid derivatives causing adverse effects in therapeutic use
C0851314|T037|AB|E932.8|ICD9CM|Adv eff antithyroid agnt|Adv eff antithyroid agnt
C0851314|T037|PT|E932.8|ICD9CM|Antithyroid agents causing adverse effects in therapeutic use|Antithyroid agents causing adverse effects in therapeutic use
C0261793|T037|AB|E932.9|ICD9CM|Adv eff hormones NEC/NOS|Adv eff hormones NEC/NOS
C0261793|T037|PT|E932.9|ICD9CM|Other and unspecified hormones and synthetic substitutes causing adverse effects in therapeutic use|Other and unspecified hormones and synthetic substitutes causing adverse effects in therapeutic use
C0261794|T046|HT|E933|ICD9CM|Primarily systemic agents causing adverse effects in therapeutic use|Primarily systemic agents causing adverse effects in therapeutic use
C0261795|T046|AB|E933.0|ICD9CM|Adv eff anallrg/antemet|Adv eff anallrg/antemet
C0261795|T046|PT|E933.0|ICD9CM|Antiallergic and antiemetic drugs causing adverse effects in therapeutic use|Antiallergic and antiemetic drugs causing adverse effects in therapeutic use
C0261796|T037|AB|E933.1|ICD9CM|Adv eff antineoplastic|Adv eff antineoplastic
C0261796|T037|PT|E933.1|ICD9CM|Antineoplastic and immunosuppressive drugs causing adverse effects in therapeutic use|Antineoplastic and immunosuppressive drugs causing adverse effects in therapeutic use
C0261797|T037|PT|E933.2|ICD9CM|Acidifying agents causing adverse effects in therapeutic use|Acidifying agents causing adverse effects in therapeutic use
C0261797|T037|AB|E933.2|ICD9CM|Adv eff acidifying agent|Adv eff acidifying agent
C0261798|T037|AB|E933.3|ICD9CM|Adv eff alkalizing agent|Adv eff alkalizing agent
C0261798|T037|PT|E933.3|ICD9CM|Alkalizing agents causing adverse effects in therapeutic use|Alkalizing agents causing adverse effects in therapeutic use
C0869502|T037|AB|E933.4|ICD9CM|Adv eff enzymes NEC|Adv eff enzymes NEC
C0869502|T037|PT|E933.4|ICD9CM|Enzymes, not elsewhere classified, causing adverse effects in therapeutic use|Enzymes, not elsewhere classified, causing adverse effects in therapeutic use
C0869504|T037|AB|E933.5|ICD9CM|Adv eff vitamins NEC|Adv eff vitamins NEC
C0869504|T037|PT|E933.5|ICD9CM|Vitamins, not elsewhere classified, causing adverse effects in therapeutic use|Vitamins, not elsewhere classified, causing adverse effects in therapeutic use
C1955565|T037|AB|E933.6|ICD9CM|Oral bisphosphonates|Oral bisphosphonates
C1955565|T037|PT|E933.6|ICD9CM|Oral bisphosphonates|Oral bisphosphonates
C1955566|T047|PT|E933.7|ICD9CM|Intravenous bisphosphonates|Intravenous bisphosphonates
C1955566|T047|AB|E933.7|ICD9CM|IV bisphosphonates|IV bisphosphonates
C0261801|T037|AB|E933.8|ICD9CM|Adv eff systemic agt NEC|Adv eff systemic agt NEC
C0261801|T037|PT|E933.8|ICD9CM|Other systemic agents, not elsewhere classified, causing adverse effects in therapeutic use|Other systemic agents, not elsewhere classified, causing adverse effects in therapeutic use
C0261802|T037|AB|E933.9|ICD9CM|Adv eff systemic agt NOS|Adv eff systemic agt NOS
C0261802|T037|PT|E933.9|ICD9CM|Unspecified systemic agent causing adverse effects in therapeutic use|Unspecified systemic agent causing adverse effects in therapeutic use
C0261803|T046|HT|E934|ICD9CM|Agents primarily affecting blood constituents causing adverse effects in therapeutic use|Agents primarily affecting blood constituents causing adverse effects in therapeutic use
C0261804|T037|AB|E934.0|ICD9CM|Adv eff iron & compounds|Adv eff iron & compounds
C0261804|T037|PT|E934.0|ICD9CM|Iron and its compounds causing adverse effects in therapeutic use|Iron and its compounds causing adverse effects in therapeutic use
C0261805|T037|AB|E934.1|ICD9CM|Adv eff liver/antianemic|Adv eff liver/antianemic
C0261805|T037|PT|E934.1|ICD9CM|Liver preparations and other antianemic agents causing adverse effects in therapeutic use|Liver preparations and other antianemic agents causing adverse effects in therapeutic use
C0261806|T037|AB|E934.2|ICD9CM|Adv eff anticoagulants|Adv eff anticoagulants
C0261806|T037|PT|E934.2|ICD9CM|Anticoagulants causing adverse effects in therapeutic use|Anticoagulants causing adverse effects in therapeutic use
C0261807|T037|AB|E934.3|ICD9CM|Adv eff vitamin k|Adv eff vitamin k
C0261807|T037|PT|E934.3|ICD9CM|Vitamin k [phytonadione] causing adverse effects in therapeutic use|Vitamin k [phytonadione] causing adverse effects in therapeutic use
C0261808|T037|AB|E934.4|ICD9CM|Adv eff fibrinolysis agt|Adv eff fibrinolysis agt
C0261808|T037|PT|E934.4|ICD9CM|Fibrinolysis-affecting drugs causing adverse effects in therapeutic use|Fibrinolysis-affecting drugs causing adverse effects in therapeutic use
C0261809|T037|AB|E934.5|ICD9CM|Adv eff coagulants|Adv eff coagulants
C0261809|T037|PT|E934.5|ICD9CM|Anticoagulant antagonists and other coagulants causing adverse effects in therapeutic use|Anticoagulant antagonists and other coagulants causing adverse effects in therapeutic use
C0261810|T037|AB|E934.6|ICD9CM|Adv eff gamma globulin|Adv eff gamma globulin
C0261810|T037|PT|E934.6|ICD9CM|Gamma globulin causing adverse effects in therapeutic use|Gamma globulin causing adverse effects in therapeutic use
C0261811|T046|AB|E934.7|ICD9CM|Adv eff blood products|Adv eff blood products
C0261811|T046|PT|E934.7|ICD9CM|Natural blood and blood products causing adverse effects in therapeutic use|Natural blood and blood products causing adverse effects in therapeutic use
C0261812|T037|AB|E934.8|ICD9CM|Adv eff blood agent NEC|Adv eff blood agent NEC
C0261812|T037|PT|E934.8|ICD9CM|Other agents affecting blood constituents causing adverse effects in therapeutic use|Other agents affecting blood constituents causing adverse effects in therapeutic use
C0261813|T037|AB|E934.9|ICD9CM|Adv eff blood agent NOS|Adv eff blood agent NOS
C0261813|T037|PT|E934.9|ICD9CM|Unspecified agent affecting blood constituents causing adverse effects in therapeutic use|Unspecified agent affecting blood constituents causing adverse effects in therapeutic use
C0261814|T037|HT|E935|ICD9CM|Analgesics, antipyretics, and antirheumatics causing adverse effects in therapeutic use|Analgesics, antipyretics, and antirheumatics causing adverse effects in therapeutic use
C0261815|T037|AB|E935.0|ICD9CM|Adv eff heroin|Adv eff heroin
C0261815|T037|PT|E935.0|ICD9CM|Heroin causing adverse effects in therapeutic use|Heroin causing adverse effects in therapeutic use
C0261816|T046|AB|E935.1|ICD9CM|Adv eff methadone|Adv eff methadone
C0261816|T046|PT|E935.1|ICD9CM|Methadone causing averse effects in therapeutic use|Methadone causing averse effects in therapeutic use
C0261817|T037|AB|E935.2|ICD9CM|Adv eff opiates|Adv eff opiates
C0261817|T037|PT|E935.2|ICD9CM|Other opiates and related narcotics causing adverse effects in therapeutic use|Other opiates and related narcotics causing adverse effects in therapeutic use
C0851323|T037|AB|E935.3|ICD9CM|Adv eff salicylates|Adv eff salicylates
C0851323|T037|PT|E935.3|ICD9CM|Salicylates causing adverse effects in therapeutic use|Salicylates causing adverse effects in therapeutic use
C0261819|T037|AB|E935.4|ICD9CM|Adv eff arom analgsc NEC|Adv eff arom analgsc NEC
C0261819|T037|PT|E935.4|ICD9CM|Aromatic analgesics, not elsewhere classified, causing adverse effects in therapeutic use|Aromatic analgesics, not elsewhere classified, causing adverse effects in therapeutic use
C0261820|T037|AB|E935.5|ICD9CM|Adv eff pyrazole deriv|Adv eff pyrazole deriv
C0261820|T037|PT|E935.5|ICD9CM|Pyrazole derivatives causing adverse effects in therapeutic use|Pyrazole derivatives causing adverse effects in therapeutic use
C0481138|T046|AB|E935.6|ICD9CM|Adv eff antirheumatics|Adv eff antirheumatics
C0481138|T046|PT|E935.6|ICD9CM|Antirheumatics [antiphlogistics] causing adverse effects in therapeutic use|Antirheumatics [antiphlogistics] causing adverse effects in therapeutic use
C0261822|T037|AB|E935.7|ICD9CM|Adv eff non-narc analgsc|Adv eff non-narc analgsc
C0261822|T037|PT|E935.7|ICD9CM|Other non-narcotic analgesics causing adverse effects in therapeutic use|Other non-narcotic analgesics causing adverse effects in therapeutic use
C0261823|T037|AB|E935.8|ICD9CM|Adv eff analgesics NEC|Adv eff analgesics NEC
C0261823|T037|PT|E935.8|ICD9CM|Other specified analgesics and antipyretics causing adverse effects in therapeutic use|Other specified analgesics and antipyretics causing adverse effects in therapeutic use
C0261824|T037|AB|E935.9|ICD9CM|Adv eff analgesic NOS|Adv eff analgesic NOS
C0261824|T037|PT|E935.9|ICD9CM|Unspecified analgesic and antipyretic causing adverse effects in therapeutic use|Unspecified analgesic and antipyretic causing adverse effects in therapeutic use
C0481142|T037|HT|E936|ICD9CM|Anticonvulsants and anti-Parkinsonism drugs causing adverse effects in therapeutic use|Anticonvulsants and anti-Parkinsonism drugs causing adverse effects in therapeutic use
C0261826|T037|AB|E936.0|ICD9CM|Adv eff oxazolidin deriv|Adv eff oxazolidin deriv
C0261826|T037|PT|E936.0|ICD9CM|Oxazolidine derivatives causing adverse effects in therapeutic use|Oxazolidine derivatives causing adverse effects in therapeutic use
C0261827|T037|AB|E936.1|ICD9CM|Adv eff hydantoin deriv|Adv eff hydantoin deriv
C0261827|T037|PT|E936.1|ICD9CM|Hydantoin derivatives causing adverse effects in therapeutic use|Hydantoin derivatives causing adverse effects in therapeutic use
C0851324|T037|AB|E936.2|ICD9CM|Adv eff succinimides|Adv eff succinimides
C0851324|T037|PT|E936.2|ICD9CM|Succinimides causing adverse effects in therapeutic use|Succinimides causing adverse effects in therapeutic use
C0261829|T037|AB|E936.3|ICD9CM|Adv eff antconvl NEC/NOS|Adv eff antconvl NEC/NOS
C0261829|T037|PT|E936.3|ICD9CM|Other and unspecified anticonvulsants causing adverse effects in therapeutic use|Other and unspecified anticonvulsants causing adverse effects in therapeutic use
C0481147|T046|AB|E936.4|ICD9CM|Adv eff anti-parkinson|Adv eff anti-parkinson
C0481147|T046|PT|E936.4|ICD9CM|Anti-parkinsonism drugs causing adverse effects in therapeutic use|Anti-parkinsonism drugs causing adverse effects in therapeutic use
C0261831|T037|HT|E937|ICD9CM|Sedatives and hypnotics causing adverse effects in therapeutic use|Sedatives and hypnotics causing adverse effects in therapeutic use
C0261832|T037|AB|E937.0|ICD9CM|Adv eff barbiturates|Adv eff barbiturates
C0261832|T037|PT|E937.0|ICD9CM|Barbiturates causing adverse effects in therapeutic use|Barbiturates causing adverse effects in therapeutic use
C0261833|T037|AB|E937.1|ICD9CM|Adv eff chloral hydrate|Adv eff chloral hydrate
C0261833|T037|PT|E937.1|ICD9CM|Chloral hydrate group causing adverse effects in therapeutic use|Chloral hydrate group causing adverse effects in therapeutic use
C0851325|T037|AB|E937.2|ICD9CM|Adv eff paraldehyde|Adv eff paraldehyde
C0851325|T037|PT|E937.2|ICD9CM|Paraldehyde causing adverse effects in therapeutic use|Paraldehyde causing adverse effects in therapeutic use
C0261835|T037|AB|E937.3|ICD9CM|Adv eff bromine compnds|Adv eff bromine compnds
C0261835|T037|PT|E937.3|ICD9CM|Bromine compounds causing adverse effects in therapeutic use|Bromine compounds causing adverse effects in therapeutic use
C0261836|T037|AB|E937.4|ICD9CM|Adv eff methaqualone|Adv eff methaqualone
C0261836|T037|PT|E937.4|ICD9CM|Methaqualone compounds causing adverse effects in therapeutic use|Methaqualone compounds causing adverse effects in therapeutic use
C0261837|T037|AB|E937.5|ICD9CM|Adv eff glutethimide|Adv eff glutethimide
C0261837|T037|PT|E937.5|ICD9CM|Glutethimide group causing adverse effects in therapeutic use|Glutethimide group causing adverse effects in therapeutic use
C0261838|T037|AB|E937.6|ICD9CM|Adv eff mix sedative|Adv eff mix sedative
C0261838|T037|PT|E937.6|ICD9CM|Mixed sedatives, not elsewhere classified, causing adverse effects in therapeutic use|Mixed sedatives, not elsewhere classified, causing adverse effects in therapeutic use
C0261839|T037|AB|E937.8|ICD9CM|Adv eff sedat/hypnot NEC|Adv eff sedat/hypnot NEC
C0261839|T037|PT|E937.8|ICD9CM|Other sedatives and hypnotics causing adverse effects in therapeutic use|Other sedatives and hypnotics causing adverse effects in therapeutic use
C0261840|T037|AB|E937.9|ICD9CM|Adv eff sedat/hypnot NOS|Adv eff sedat/hypnot NOS
C0261840|T037|PT|E937.9|ICD9CM|Unspecified sedatives and hypnotics causing adverse effects in therapeutic use|Unspecified sedatives and hypnotics causing adverse effects in therapeutic use
C0261841|T037|HT|E938|ICD9CM|Other central nervous system depressants and anesthetics causing adverse effects in therapeutic use|Other central nervous system depressants and anesthetics causing adverse effects in therapeutic use
C0261842|T037|AB|E938.0|ICD9CM|Adv eff cns muscl depres|Adv eff cns muscl depres
C0261842|T037|PT|E938.0|ICD9CM|Central nervous system muscle-tone depressants causing adverse effects in therapeutic use|Central nervous system muscle-tone depressants causing adverse effects in therapeutic use
C0261843|T037|AB|E938.1|ICD9CM|Adv eff halothane|Adv eff halothane
C0261843|T037|PT|E938.1|ICD9CM|Halothane causing adverse effects in therapeutic use|Halothane causing adverse effects in therapeutic use
C0261844|T037|AB|E938.2|ICD9CM|Adv eff gas anesthet NEC|Adv eff gas anesthet NEC
C0261844|T037|PT|E938.2|ICD9CM|Other gaseous anesthetics causing adverse effects in therapeutic use|Other gaseous anesthetics causing adverse effects in therapeutic use
C0261845|T037|AB|E938.3|ICD9CM|Adv eff intraven anesth|Adv eff intraven anesth
C0261845|T037|PT|E938.3|ICD9CM|Intravenous anesthetics causing adverse effects in therapeutic use|Intravenous anesthetics causing adverse effects in therapeutic use
C0261846|T037|AB|E938.4|ICD9CM|Adv eff gen anes NEC/NOS|Adv eff gen anes NEC/NOS
C0261846|T037|PT|E938.4|ICD9CM|Other and unspecified general anesthetics causing adverse effects in therapeutic use|Other and unspecified general anesthetics causing adverse effects in therapeutic use
C0474019|T046|AB|E938.5|ICD9CM|Adv eff topic/infil anes|Adv eff topic/infil anes
C0474019|T046|PT|E938.5|ICD9CM|Surface and infiltration anesthetics causing adverse effects in therapeutic use|Surface and infiltration anesthetics causing adverse effects in therapeutic use
C0261848|T037|AB|E938.6|ICD9CM|Adv eff nerve-block anes|Adv eff nerve-block anes
C0261848|T037|PT|E938.6|ICD9CM|Peripheral nerve- and plexus-blocking anesthetics causing adverse effects in therapeutic use|Peripheral nerve- and plexus-blocking anesthetics causing adverse effects in therapeutic use
C0261849|T037|AB|E938.7|ICD9CM|Adv eff spinal anesthet|Adv eff spinal anesthet
C0261849|T037|PT|E938.7|ICD9CM|Spinal anesthetics causing adverse effects in therapeutic use|Spinal anesthetics causing adverse effects in therapeutic use
C0261850|T037|AB|E938.9|ICD9CM|Adv eff loc anes NEC/NOS|Adv eff loc anes NEC/NOS
C0261850|T037|PT|E938.9|ICD9CM|Other and unspecified local anesthetics causing adverse effects in therapeutic use|Other and unspecified local anesthetics causing adverse effects in therapeutic use
C0261851|T037|HT|E939|ICD9CM|Psychotropic agents causing adverse effects in therapeutic use|Psychotropic agents causing adverse effects in therapeutic use
C0261852|T037|AB|E939.0|ICD9CM|Adv eff antidepressants|Adv eff antidepressants
C0261852|T037|PT|E939.0|ICD9CM|Antidepressants causing adverse effects in therapeutic use|Antidepressants causing adverse effects in therapeutic use
C0261853|T037|AB|E939.1|ICD9CM|Adv eff phenothiaz tranq|Adv eff phenothiaz tranq
C0261853|T037|PT|E939.1|ICD9CM|Phenothiazine-based tranquilizers causing adverse effects in therapeutic use|Phenothiazine-based tranquilizers causing adverse effects in therapeutic use
C0261854|T037|AB|E939.2|ICD9CM|Adv eff butyrophen tranq|Adv eff butyrophen tranq
C0261854|T037|PT|E939.2|ICD9CM|Butyrophenone-based tranquilizers causing adverse effects in therapeutic use|Butyrophenone-based tranquilizers causing adverse effects in therapeutic use
C0261855|T037|AB|E939.3|ICD9CM|Adv eff antipsychotc NEC|Adv eff antipsychotc NEC
C0261856|T037|AB|E939.4|ICD9CM|Adv eff benzodiaz tranq|Adv eff benzodiaz tranq
C0261856|T037|PT|E939.4|ICD9CM|Benzodiazepine-based tranquilizers causing adverse effects in therapeutic use|Benzodiazepine-based tranquilizers causing adverse effects in therapeutic use
C0261857|T037|AB|E939.5|ICD9CM|Adv eff tranquilizer NEC|Adv eff tranquilizer NEC
C0261857|T037|PT|E939.5|ICD9CM|Other tranquilizers causing adverse effects in therapeutic use|Other tranquilizers causing adverse effects in therapeutic use
C0261858|T037|AB|E939.6|ICD9CM|Adv eff hallucinogens|Adv eff hallucinogens
C0261858|T037|PT|E939.6|ICD9CM|Psychodysleptics [hallucinogens] causing adverse effects in therapeutic use|Psychodysleptics [hallucinogens] causing adverse effects in therapeutic use
C0261859|T037|AB|E939.7|ICD9CM|Adv eff psychostimulants|Adv eff psychostimulants
C0261859|T037|PT|E939.7|ICD9CM|Psychostimulants causing adverse effects in therapeutic use|Psychostimulants causing adverse effects in therapeutic use
C0261860|T037|AB|E939.8|ICD9CM|Adv eff psychotropic NEC|Adv eff psychotropic NEC
C0261860|T037|PT|E939.8|ICD9CM|Other psychotropic agents causing adverse effects in therapeutic use|Other psychotropic agents causing adverse effects in therapeutic use
C0261861|T037|AB|E939.9|ICD9CM|Adv eff psychotropic NOS|Adv eff psychotropic NOS
C0261861|T037|PT|E939.9|ICD9CM|Unspecified psychotropic agent causing adverse effects in therapeutic use|Unspecified psychotropic agent causing adverse effects in therapeutic use
C0569621|T046|HT|E940|ICD9CM|Central nervous system stimulants causing adverse effects in therapeutic use|Central nervous system stimulants causing adverse effects in therapeutic use
C0261863|T046|AB|E940.0|ICD9CM|Adv eff analeptics|Adv eff analeptics
C0261863|T046|PT|E940.0|ICD9CM|Analeptics causing adverse effects in therapeutic use|Analeptics causing adverse effects in therapeutic use
C0261864|T037|AB|E940.1|ICD9CM|Adv eff opiat antagonist|Adv eff opiat antagonist
C0261864|T037|PT|E940.1|ICD9CM|Opiate antagonists causing adverse effects in therapeutic use|Opiate antagonists causing adverse effects in therapeutic use
C0261865|T037|AB|E940.8|ICD9CM|Adv eff cns stimulnt NEC|Adv eff cns stimulnt NEC
C0261865|T037|PT|E940.8|ICD9CM|Other specified central nervous system stimulants causing adverse effects in therapeutic use|Other specified central nervous system stimulants causing adverse effects in therapeutic use
C0569621|T046|AB|E940.9|ICD9CM|Adv eff cns stimulnt NOS|Adv eff cns stimulnt NOS
C0569621|T046|PT|E940.9|ICD9CM|Unspecified central nervous system stimulant causing adverse effects in therapeutic use|Unspecified central nervous system stimulant causing adverse effects in therapeutic use
C0543418|T046|HT|E941|ICD9CM|Drugs primarily affecting the autonomic nervous system causing adverse effects in therapeutic use|Drugs primarily affecting the autonomic nervous system causing adverse effects in therapeutic use
C0261868|T037|AB|E941.0|ICD9CM|Adv eff cholinergics|Adv eff cholinergics
C0261868|T037|PT|E941.0|ICD9CM|Parasympathomimetics [cholinergics] causing adverse effects in therapeutic use|Parasympathomimetics [cholinergics] causing adverse effects in therapeutic use
C0261869|T037|AB|E941.1|ICD9CM|Adv eff parasympatholytc|Adv eff parasympatholytc
C0261870|T037|AB|E941.2|ICD9CM|Adv eff sympathomimetics|Adv eff sympathomimetics
C0261870|T037|PT|E941.2|ICD9CM|Sympathomimetics [adrenergics] causing adverse effects in therapeutic use|Sympathomimetics [adrenergics] causing adverse effects in therapeutic use
C0261871|T037|AB|E941.3|ICD9CM|Adv eff sympatholytics|Adv eff sympatholytics
C0261871|T037|PT|E941.3|ICD9CM|Sympatholytics [antiadrenergics] causing adverse effects in therapeutic use|Sympatholytics [antiadrenergics] causing adverse effects in therapeutic use
C0261872|T037|AB|E941.9|ICD9CM|Adv eff autonom agnt NOS|Adv eff autonom agnt NOS
C1533672|T046|HT|E942|ICD9CM|Agents primarily affecting the cardiovascular system causing adverse effects in therapeutic use|Agents primarily affecting the cardiovascular system causing adverse effects in therapeutic use
C0261874|T037|AB|E942.0|ICD9CM|Adv eff card rhyth regul|Adv eff card rhyth regul
C0261874|T037|PT|E942.0|ICD9CM|Cardiac rhythm regulators causing adverse effects in therapeutic use|Cardiac rhythm regulators causing adverse effects in therapeutic use
C0261875|T037|AB|E942.1|ICD9CM|Adv eff cardiotonics|Adv eff cardiotonics
C0261875|T037|PT|E942.1|ICD9CM|Cardiotonic glycosides and drugs of similar action causing adverse effects in therapeutic use|Cardiotonic glycosides and drugs of similar action causing adverse effects in therapeutic use
C0481188|T037|AB|E942.2|ICD9CM|Adv eff antilipemics|Adv eff antilipemics
C0481188|T037|PT|E942.2|ICD9CM|Antilipemic and antiarteriosclerotic drugs causing adverse effects in therapeutic use|Antilipemic and antiarteriosclerotic drugs causing adverse effects in therapeutic use
C0261877|T037|AB|E942.3|ICD9CM|Adv eff ganglion-block|Adv eff ganglion-block
C0261877|T037|PT|E942.3|ICD9CM|Ganglion-blocking agents causing adverse effects in therapeutic use|Ganglion-blocking agents causing adverse effects in therapeutic use
C0261878|T037|AB|E942.4|ICD9CM|Adv eff coronary vasodil|Adv eff coronary vasodil
C0261878|T037|PT|E942.4|ICD9CM|Coronary vasodilators causing adverse effects in therapeutic use|Coronary vasodilators causing adverse effects in therapeutic use
C0261879|T037|AB|E942.5|ICD9CM|Adv eff vasodilators NEC|Adv eff vasodilators NEC
C0261879|T037|PT|E942.5|ICD9CM|Other vasodilators causing adverse effects in therapeutic use|Other vasodilators causing adverse effects in therapeutic use
C0261880|T037|AB|E942.6|ICD9CM|Adv eff antihyperten agt|Adv eff antihyperten agt
C0261880|T037|PT|E942.6|ICD9CM|Other antihypertensive agents causing adverse effects in therapeutic use|Other antihypertensive agents causing adverse effects in therapeutic use
C0497073|T037|AB|E942.7|ICD9CM|Adv eff antivaricose|Adv eff antivaricose
C0497073|T037|PT|E942.7|ICD9CM|Antivaricose drugs, including sclerosing agents, causing adverse effects in therapeutic use|Antivaricose drugs, including sclerosing agents, causing adverse effects in therapeutic use
C0261882|T037|AB|E942.8|ICD9CM|Adv eff capillary-act|Adv eff capillary-act
C0261882|T037|PT|E942.8|ICD9CM|Capillary-active drugs causing adverse effects in therapeutic use|Capillary-active drugs causing adverse effects in therapeutic use
C0497074|T037|AB|E942.9|ICD9CM|Adv eff cardiovasc NEC|Adv eff cardiovasc NEC
C0413956|T046|HT|E943|ICD9CM|Agents primarily affecting gastrointestinal system causing adverse effects in therapeutic use|Agents primarily affecting gastrointestinal system causing adverse effects in therapeutic use
C0261885|T037|AB|E943.0|ICD9CM|Adv eff antacids|Adv eff antacids
C0261885|T037|PT|E943.0|ICD9CM|Antacids and antigastric secretion drugs causing adverse effects in therapeutic use|Antacids and antigastric secretion drugs causing adverse effects in therapeutic use
C0261886|T037|AB|E943.1|ICD9CM|Adv eff irrit cathartic|Adv eff irrit cathartic
C0261886|T037|PT|E943.1|ICD9CM|Irritant cathartics causing adverse effects in therapeutic use|Irritant cathartics causing adverse effects in therapeutic use
C0261887|T037|AB|E943.2|ICD9CM|Adv eff emoll cathartics|Adv eff emoll cathartics
C0261887|T037|PT|E943.2|ICD9CM|Emollient cathartics causing adverse effects in therapeutic use|Emollient cathartics causing adverse effects in therapeutic use
C0261888|T037|AB|E943.3|ICD9CM|Adv eff cathartics NEC|Adv eff cathartics NEC
C0261888|T037|PT|E943.3|ICD9CM|Other cathartics, including intestinal atonia drugs, causing adverse effects in therapeutic use|Other cathartics, including intestinal atonia drugs, causing adverse effects in therapeutic use
C0261889|T046|AB|E943.4|ICD9CM|Adv eff digestants|Adv eff digestants
C0261889|T046|PT|E943.4|ICD9CM|Digestants causing adverse effects in therapeutic use|Digestants causing adverse effects in therapeutic use
C0474035|T046|AB|E943.5|ICD9CM|Adv eff antidiarrhea agt|Adv eff antidiarrhea agt
C0474035|T046|PT|E943.5|ICD9CM|Antidiarrheal drugs causing adverse effects in therapeutic use|Antidiarrheal drugs causing adverse effects in therapeutic use
C0261891|T046|AB|E943.6|ICD9CM|Adv eff emetics|Adv eff emetics
C0261891|T046|PT|E943.6|ICD9CM|Emetics causing adverse effects in therapeutic use|Emetics causing adverse effects in therapeutic use
C0261892|T037|AB|E943.8|ICD9CM|Adv eff GI agent NEC|Adv eff GI agent NEC
C0413956|T046|AB|E943.9|ICD9CM|Adv eff GI agent NOS|Adv eff GI agent NOS
C0261894|T037|HT|E944|ICD9CM|Water, mineral, and uric acid metabolism drugs causing adverse effects in therapeutic use|Water, mineral, and uric acid metabolism drugs causing adverse effects in therapeutic use
C0261895|T037|AB|E944.0|ICD9CM|Adv eff mercury diuretic|Adv eff mercury diuretic
C0261895|T037|PT|E944.0|ICD9CM|Mercurial diuretics causing adverse effects in therapeutic use|Mercurial diuretics causing adverse effects in therapeutic use
C0261896|T037|AB|E944.1|ICD9CM|Adv eff purine diuretics|Adv eff purine diuretics
C0261896|T037|PT|E944.1|ICD9CM|Purine derivative diuretics causing adverse effects in therapeutic use|Purine derivative diuretics causing adverse effects in therapeutic use
C0481197|T037|AB|E944.2|ICD9CM|Adv eff acetazolamide|Adv eff acetazolamide
C0481197|T037|PT|E944.2|ICD9CM|Carbonic acid anhydrase inhibitors causing adverse effects in therapeutic use|Carbonic acid anhydrase inhibitors causing adverse effects in therapeutic use
C0261898|T037|AB|E944.3|ICD9CM|Adv eff saluretics|Adv eff saluretics
C0261898|T037|PT|E944.3|ICD9CM|Saluretics causing adverse effects in therapeutic use|Saluretics causing adverse effects in therapeutic use
C0261899|T037|AB|E944.4|ICD9CM|Adv eff diuretics NEC|Adv eff diuretics NEC
C0261899|T037|PT|E944.4|ICD9CM|Other diuretics causing adverse effects in therapeutic use|Other diuretics causing adverse effects in therapeutic use
C0497076|T046|AB|E944.5|ICD9CM|Adv eff electrolyte agnt|Adv eff electrolyte agnt
C0497076|T046|PT|E944.5|ICD9CM|Electrolytic, caloric, and water-balance agents causing adverse effects in therapeutic use|Electrolytic, caloric, and water-balance agents causing adverse effects in therapeutic use
C0261901|T037|AB|E944.6|ICD9CM|Adv eff mineral salt NEC|Adv eff mineral salt NEC
C0261901|T037|PT|E944.6|ICD9CM|Other mineral salts, not elsewhere classified, causing adverse effects in therapeutic use|Other mineral salts, not elsewhere classified, causing adverse effects in therapeutic use
C0261902|T037|AB|E944.7|ICD9CM|Adv eff uric acid metab|Adv eff uric acid metab
C0261902|T037|PT|E944.7|ICD9CM|Uric acid metabolism drugs causing adverse effects in therapeutic use|Uric acid metabolism drugs causing adverse effects in therapeutic use
C0414020|T046|AB|E945.0|ICD9CM|Adv eff oxytocic agents|Adv eff oxytocic agents
C0414020|T046|PT|E945.0|ICD9CM|Oxytocic agents causing adverse effects in therapeutic use|Oxytocic agents causing adverse effects in therapeutic use
C0261905|T037|AB|E945.1|ICD9CM|Adv eff smooth musc relx|Adv eff smooth musc relx
C0261905|T037|PT|E945.1|ICD9CM|Smooth muscle relaxants causing adverse effects in therapeutic use|Smooth muscle relaxants causing adverse effects in therapeutic use
C0481202|T037|AB|E945.2|ICD9CM|Adv eff skelet musc relx|Adv eff skelet musc relx
C0481202|T037|PT|E945.2|ICD9CM|Skeletal muscle relaxants causing adverse effects in therapeutic use|Skeletal muscle relaxants causing adverse effects in therapeutic use
C0261907|T037|AB|E945.3|ICD9CM|Adv eff musc agt NEC/NOS|Adv eff musc agt NEC/NOS
C0261907|T037|PT|E945.3|ICD9CM|Other and unspecified drugs acting on muscles causing adverse effects in therapeutic use|Other and unspecified drugs acting on muscles causing adverse effects in therapeutic use
C0261908|T046|AB|E945.4|ICD9CM|Adv eff antitussives|Adv eff antitussives
C0261908|T046|PT|E945.4|ICD9CM|Antitussives causing adverse effects in therapeutic use|Antitussives causing adverse effects in therapeutic use
C0851326|T037|AB|E945.5|ICD9CM|Adv eff expectorants|Adv eff expectorants
C0851326|T037|PT|E945.5|ICD9CM|Expectorants causing adverse effects in therapeutic use|Expectorants causing adverse effects in therapeutic use
C0414040|T046|AB|E945.6|ICD9CM|Adv eff anti-common cold|Adv eff anti-common cold
C0414040|T046|PT|E945.6|ICD9CM|Anti-common cold drugs causing adverse effects in therapeutic use|Anti-common cold drugs causing adverse effects in therapeutic use
C0261911|T037|AB|E945.7|ICD9CM|Adv eff antiasthmatics|Adv eff antiasthmatics
C0261911|T037|PT|E945.7|ICD9CM|Antiasthmatics causing adverse effects in therapeutic use|Antiasthmatics causing adverse effects in therapeutic use
C0261912|T037|AB|E945.8|ICD9CM|Adv eff resp drg NEC/NOS|Adv eff resp drg NEC/NOS
C0261912|T037|PT|E945.8|ICD9CM|Other and unspecified respiratory drugs causing adverse effects in therapeutic use|Other and unspecified respiratory drugs causing adverse effects in therapeutic use
C0261914|T037|AB|E946.0|ICD9CM|Adv eff loc anti-infectv|Adv eff loc anti-infectv
C0261914|T037|PT|E946.0|ICD9CM|Local anti-infectives and anti-inflammatory drugs causing adverse effects in therapeutic use|Local anti-infectives and anti-inflammatory drugs causing adverse effects in therapeutic use
C0261915|T046|AB|E946.1|ICD9CM|Adv eff antipruritics|Adv eff antipruritics
C0261915|T046|PT|E946.1|ICD9CM|Antipruritics causing adverse effects in therapeutic use|Antipruritics causing adverse effects in therapeutic use
C0414053|T046|AB|E946.2|ICD9CM|Adv eff local astringent|Adv eff local astringent
C0414053|T046|PT|E946.2|ICD9CM|Local astringents and local detergents causing adverse effects in therapeutic use|Local astringents and local detergents causing adverse effects in therapeutic use
C0414054|T046|AB|E946.3|ICD9CM|Adv eff emollient/demulc|Adv eff emollient/demulc
C0414054|T046|PT|E946.3|ICD9CM|Emollients, demulcents, and protectants causing adverse effects in therapeutic use|Emollients, demulcents, and protectants causing adverse effects in therapeutic use
C0414055|T046|AB|E946.4|ICD9CM|Adv eff hair/scalp prep|Adv eff hair/scalp prep
C0261919|T037|AB|E946.5|ICD9CM|Adv eff eye anti-inf/drg|Adv eff eye anti-inf/drg
C0261919|T037|PT|E946.5|ICD9CM|Eye anti-infectives and other eye drugs causing adverse effects in therapeutic use|Eye anti-infectives and other eye drugs causing adverse effects in therapeutic use
C0261920|T037|AB|E946.6|ICD9CM|Adv eff ent anti-inf/drg|Adv eff ent anti-inf/drg
C0261921|T046|AB|E946.7|ICD9CM|Adv eff topic dental drg|Adv eff topic dental drg
C0261921|T046|PT|E946.7|ICD9CM|Dental drugs topically applied causing adverse effects in therapeutic use|Dental drugs topically applied causing adverse effects in therapeutic use
C0261922|T037|AB|E946.8|ICD9CM|Adv eff skin agent NEC|Adv eff skin agent NEC
C0261922|T037|PT|E946.8|ICD9CM|Other agents primarily affecting skin and mucous membrane causing adverse effects in therapeutic use|Other agents primarily affecting skin and mucous membrane causing adverse effects in therapeutic use
C0261923|T037|AB|E946.9|ICD9CM|Adv eff skin agent NOS|Adv eff skin agent NOS
C0261930|T037|HT|E947|ICD9CM|Other and unspecified drugs and medicinal substances causing adverse effects in therapeutic use|Other and unspecified drugs and medicinal substances causing adverse effects in therapeutic use
C0261925|T037|AB|E947.0|ICD9CM|Adv eff dietetics|Adv eff dietetics
C0261925|T037|PT|E947.0|ICD9CM|Dietetics causing adverse effects in therapeutic use|Dietetics causing adverse effects in therapeutic use
C0261926|T046|AB|E947.1|ICD9CM|Adv eff lipotropic drugs|Adv eff lipotropic drugs
C0261926|T046|PT|E947.1|ICD9CM|Lipotropic drugs causing adverse effects in therapeutic use|Lipotropic drugs causing adverse effects in therapeutic use
C1963710|T037|AB|E947.2|ICD9CM|Adv eff antidotes NEC|Adv eff antidotes NEC
C1963710|T037|PT|E947.2|ICD9CM|Antidotes and chelating agents, not elsewhere classified, causing adverse effects in therapeutic use|Antidotes and chelating agents, not elsewhere classified, causing adverse effects in therapeutic use
C0261928|T046|AB|E947.3|ICD9CM|Adv eff alcohol deter|Adv eff alcohol deter
C0261928|T046|PT|E947.3|ICD9CM|Alcohol deterrents causing adverse effects in therapeutic use|Alcohol deterrents causing adverse effects in therapeutic use
C0261929|T046|AB|E947.4|ICD9CM|Adv eff pharmaceut excip|Adv eff pharmaceut excip
C0261929|T046|PT|E947.4|ICD9CM|Pharmaceutical excipients causing adverse effects in therapeutic use|Pharmaceutical excipients causing adverse effects in therapeutic use
C0261930|T037|AB|E947.8|ICD9CM|Adv eff medicinal NEC|Adv eff medicinal NEC
C0261930|T037|PT|E947.8|ICD9CM|Other drugs and medicinal substances causing adverse effects in therapeutic use|Other drugs and medicinal substances causing adverse effects in therapeutic use
C0041831|T037|AB|E947.9|ICD9CM|Adv eff medicinal NOS|Adv eff medicinal NOS
C0041831|T037|PT|E947.9|ICD9CM|Unspecified drug or medicinal substance causing adverse effects in therapeutic use|Unspecified drug or medicinal substance causing adverse effects in therapeutic use
C0851327|T037|HT|E948|ICD9CM|Bacterial vaccines causing adverse effects in therapeutic use|Bacterial vaccines causing adverse effects in therapeutic use
C0851328|T046|AB|E948.0|ICD9CM|Adv eff bcg vaccine|Adv eff bcg vaccine
C0851328|T046|PT|E948.0|ICD9CM|Bcg vaccine causing adverse effects in therapeutic use|Bcg vaccine causing adverse effects in therapeutic use
C0261933|T046|AB|E948.1|ICD9CM|Adv eff typhoid vaccine|Adv eff typhoid vaccine
C0261933|T046|PT|E948.1|ICD9CM|Typhoid and paratyphoid vaccines causing adverse effects in therapeutic use|Typhoid and paratyphoid vaccines causing adverse effects in therapeutic use
C0261934|T037|AB|E948.2|ICD9CM|Adv eff cholera vaccine|Adv eff cholera vaccine
C0261934|T037|PT|E948.2|ICD9CM|Cholera vaccine causing adverse effects in therapeutic use|Cholera vaccine causing adverse effects in therapeutic use
C0851329|T037|AB|E948.3|ICD9CM|Adv eff plague vaccine|Adv eff plague vaccine
C0851329|T037|PT|E948.3|ICD9CM|Plague vaccine causing adverse effects in therapeutic use|Plague vaccine causing adverse effects in therapeutic use
C0261936|T037|AB|E948.4|ICD9CM|Adv eff tetanus vaccine|Adv eff tetanus vaccine
C0261936|T037|PT|E948.4|ICD9CM|Tetanus vaccine causing adverse effects in therapeutic use|Tetanus vaccine causing adverse effects in therapeutic use
C0261937|T037|AB|E948.5|ICD9CM|Adv eff diphther vaccine|Adv eff diphther vaccine
C0261937|T037|PT|E948.5|ICD9CM|Diphtheria vaccine causing adverse effects in therapeutic use|Diphtheria vaccine causing adverse effects in therapeutic use
C0261938|T046|AB|E948.6|ICD9CM|Adv eff pertussis vaccin|Adv eff pertussis vaccin
C0261939|T037|AB|E948.8|ICD9CM|Adv eff bact vac NEC/NOS|Adv eff bact vac NEC/NOS
C0261939|T037|PT|E948.8|ICD9CM|Other and unspecified bacterial vaccines causing adverse effects in therapeutic use|Other and unspecified bacterial vaccines causing adverse effects in therapeutic use
C0261940|T046|AB|E948.9|ICD9CM|Adv eff mix bact vaccine|Adv eff mix bact vaccine
C0261950|T046|HT|E949|ICD9CM|Other vaccines and biological substances causing adverse effects in therapeutic use|Other vaccines and biological substances causing adverse effects in therapeutic use
C0261942|T037|AB|E949.0|ICD9CM|Adv eff smallpox vaccine|Adv eff smallpox vaccine
C0261942|T037|PT|E949.0|ICD9CM|Smallpox vaccine causing adverse effects in therapeutic use|Smallpox vaccine causing adverse effects in therapeutic use
C0261943|T037|AB|E949.1|ICD9CM|Adv eff rabies vaccine|Adv eff rabies vaccine
C0261943|T037|PT|E949.1|ICD9CM|Rabies vaccine causing adverse effects in therapeutic use|Rabies vaccine causing adverse effects in therapeutic use
C0261944|T037|AB|E949.2|ICD9CM|Adv eff typhus vaccine|Adv eff typhus vaccine
C0261944|T037|PT|E949.2|ICD9CM|Typhus vaccine causing adverse effects in therapeutic use|Typhus vaccine causing adverse effects in therapeutic use
C0261945|T037|AB|E949.3|ICD9CM|Adv eff yellow fever vac|Adv eff yellow fever vac
C0261945|T037|PT|E949.3|ICD9CM|Yellow fever vaccine causing adverse effects in therapeutic use|Yellow fever vaccine causing adverse effects in therapeutic use
C0261946|T037|AB|E949.4|ICD9CM|Adv eff measles vaccine|Adv eff measles vaccine
C0261946|T037|PT|E949.4|ICD9CM|Measles vaccine causing adverse effects in therapeutic use|Measles vaccine causing adverse effects in therapeutic use
C0261947|T037|AB|E949.5|ICD9CM|Adv eff polio vaccine|Adv eff polio vaccine
C0261947|T037|PT|E949.5|ICD9CM|Poliomyelitis vaccine causing adverse effects in therapeutic use|Poliomyelitis vaccine causing adverse effects in therapeutic use
C0261948|T037|AB|E949.6|ICD9CM|Adv eff viral vacc NEC|Adv eff viral vacc NEC
C0261948|T037|PT|E949.6|ICD9CM|Other and unspecified viral and rickettsial vaccines causing adverse effects in therapeutic use|Other and unspecified viral and rickettsial vaccines causing adverse effects in therapeutic use
C0261949|T037|AB|E949.7|ICD9CM|Adv eff mixed viral-bact|Adv eff mixed viral-bact
C0261950|T046|AB|E949.9|ICD9CM|Adv eff biologic NEC/NOS|Adv eff biologic NEC/NOS
C0261950|T046|PT|E949.9|ICD9CM|Other and unspecified vaccines and biological substances causing adverse effects in therapeutic use|Other and unspecified vaccines and biological substances causing adverse effects in therapeutic use
C0261951|T037|HT|E950|ICD9CM|Suicide and self-inflicted poisoning by solid or liquid substances|Suicide and self-inflicted poisoning by solid or liquid substances
C0178360|T037|HT|E950-E959.9|ICD9CM|SUICIDE AND SELF-INFLICTED INJURY|SUICIDE AND SELF-INFLICTED INJURY
C0261952|T037|AB|E950.0|ICD9CM|Poison-analgesics|Poison-analgesics
C0261952|T037|PT|E950.0|ICD9CM|Suicide and self-inflicted poisoning by analgesics, antipyretics, and antirheumatics|Suicide and self-inflicted poisoning by analgesics, antipyretics, and antirheumatics
C0261953|T037|AB|E950.1|ICD9CM|Poison-barbiturates|Poison-barbiturates
C0261953|T037|PT|E950.1|ICD9CM|Suicide and self-inflicted poisoning by barbiturates|Suicide and self-inflicted poisoning by barbiturates
C0261954|T037|AB|E950.2|ICD9CM|Poison-sedat/hypnotic|Poison-sedat/hypnotic
C0261954|T037|PT|E950.2|ICD9CM|Suicide and self-inflicted poisoning by other sedatives and hypnotics|Suicide and self-inflicted poisoning by other sedatives and hypnotics
C0261955|T037|AB|E950.3|ICD9CM|Poison-psychotropic agt|Poison-psychotropic agt
C0261955|T037|PT|E950.3|ICD9CM|Suicide and self-inflicted poisoning by tranquilizers and other psychotropic agents|Suicide and self-inflicted poisoning by tranquilizers and other psychotropic agents
C0261956|T037|AB|E950.4|ICD9CM|Poison-drug/medicin NEC|Poison-drug/medicin NEC
C0261956|T037|PT|E950.4|ICD9CM|Suicide and self-inflicted poisoning by other specified drugs and medicinal substances|Suicide and self-inflicted poisoning by other specified drugs and medicinal substances
C0261957|T037|AB|E950.5|ICD9CM|Poison-drug/medicin NOS|Poison-drug/medicin NOS
C0261957|T037|PT|E950.5|ICD9CM|Suicide and self-inflicted poisoning by unspecified drug or medicinal substance|Suicide and self-inflicted poisoning by unspecified drug or medicinal substance
C0261958|T037|AB|E950.6|ICD9CM|Poison-agricult agent|Poison-agricult agent
C0261959|T037|AB|E950.7|ICD9CM|Poison-corrosiv/caustic|Poison-corrosiv/caustic
C0261959|T037|PT|E950.7|ICD9CM|Suicide and self-inflicted poisoning by corrosive and caustic substances|Suicide and self-inflicted poisoning by corrosive and caustic substances
C0261960|T037|AB|E950.8|ICD9CM|Poison-arsenic|Poison-arsenic
C0261960|T037|PT|E950.8|ICD9CM|Suicide and self-inflicted poisoning by arsenic and its compounds|Suicide and self-inflicted poisoning by arsenic and its compounds
C0261961|T037|AB|E950.9|ICD9CM|Poison-solid/liquid NEC|Poison-solid/liquid NEC
C0261961|T037|PT|E950.9|ICD9CM|Suicide and self-inflicted poisoning by other and unspecified solid and liquid substances|Suicide and self-inflicted poisoning by other and unspecified solid and liquid substances
C0261962|T037|HT|E951|ICD9CM|Suicide and self-inflicted poisoning by gases in domestic use|Suicide and self-inflicted poisoning by gases in domestic use
C0261963|T037|AB|E951.0|ICD9CM|Poison-piped gas|Poison-piped gas
C0261963|T037|PT|E951.0|ICD9CM|Suicide and self-inflicted poisoning by gas distributed by pipeline|Suicide and self-inflicted poisoning by gas distributed by pipeline
C0261964|T037|AB|E951.1|ICD9CM|Poison-gas in container|Poison-gas in container
C0261964|T037|PT|E951.1|ICD9CM|Suicide and self-inflicted poisoning by liquefied petroleum gas distributed in mobile containers|Suicide and self-inflicted poisoning by liquefied petroleum gas distributed in mobile containers
C0261965|T037|AB|E951.8|ICD9CM|Poison-utility gas NEC|Poison-utility gas NEC
C0261965|T037|PT|E951.8|ICD9CM|Suicide and self-inflicted poisoning by other utility gas|Suicide and self-inflicted poisoning by other utility gas
C0261966|T037|HT|E952|ICD9CM|Suicide and self-inflicted poisoning by other gases and vapors|Suicide and self-inflicted poisoning by other gases and vapors
C0261967|T037|AB|E952.0|ICD9CM|Poison-exhaust gas|Poison-exhaust gas
C0261967|T037|PT|E952.0|ICD9CM|Suicide and self-inflicted poisoning by motor vehicle exhaust gas|Suicide and self-inflicted poisoning by motor vehicle exhaust gas
C0261968|T037|AB|E952.1|ICD9CM|Poison-co NEC|Poison-co NEC
C0261968|T037|PT|E952.1|ICD9CM|Suicide and self-inflicted poisoning by other carbon monoxide|Suicide and self-inflicted poisoning by other carbon monoxide
C0261969|T037|AB|E952.8|ICD9CM|Poison-gas/vapor NEC|Poison-gas/vapor NEC
C0261969|T037|PT|E952.8|ICD9CM|Suicide and self-inflicted poisoning by other specified gases and vapors|Suicide and self-inflicted poisoning by other specified gases and vapors
C0261970|T037|AB|E952.9|ICD9CM|Poison-gas/vapor NOS|Poison-gas/vapor NOS
C0261970|T037|PT|E952.9|ICD9CM|Suicide and self-inflicted poisoning by unspecified gases and vapors|Suicide and self-inflicted poisoning by unspecified gases and vapors
C0261971|T037|HT|E953|ICD9CM|Suicide and self-inflicted injury by hanging, strangulation, and suffocation|Suicide and self-inflicted injury by hanging, strangulation, and suffocation
C0261972|T037|AB|E953.0|ICD9CM|Injury-hanging|Injury-hanging
C0261972|T037|PT|E953.0|ICD9CM|Suicide and self-inflicted injury by hanging|Suicide and self-inflicted injury by hanging
C0261973|T037|AB|E953.1|ICD9CM|Injury-suff w plas bag|Injury-suff w plas bag
C0261973|T037|PT|E953.1|ICD9CM|Suicide and self-inflicted injury by suffocation by plastic bag|Suicide and self-inflicted injury by suffocation by plastic bag
C0261974|T037|AB|E953.8|ICD9CM|Injury-strang/suff NEC|Injury-strang/suff NEC
C0261974|T037|PT|E953.8|ICD9CM|Suicide and self-inflicted injury by other specified means|Suicide and self-inflicted injury by other specified means
C0038662|T037|AB|E953.9|ICD9CM|Injury-strang/suff NOS|Injury-strang/suff NOS
C0038662|T037|PT|E953.9|ICD9CM|Suicide and self-inflicted injury by unspecified means|Suicide and self-inflicted injury by unspecified means
C0558960|T037|AB|E954|ICD9CM|Injury-submersion|Injury-submersion
C0558960|T037|PT|E954|ICD9CM|Suicide and self-inflicted injury by submersion [drowning]|Suicide and self-inflicted injury by submersion [drowning]
C0490043|T037|HT|E955|ICD9CM|Suicide and self-inflicted injury by firearms, air guns, and explosives|Suicide and self-inflicted injury by firearms, air guns, and explosives
C0261977|T037|AB|E955.0|ICD9CM|Injury-handgun|Injury-handgun
C0261977|T037|PT|E955.0|ICD9CM|Suicide and self-inflicted injury by handgun|Suicide and self-inflicted injury by handgun
C0261978|T037|AB|E955.1|ICD9CM|Injury-shotgun|Injury-shotgun
C0261978|T037|PT|E955.1|ICD9CM|Suicide and self-inflicted injury by shotgun|Suicide and self-inflicted injury by shotgun
C0261979|T037|AB|E955.2|ICD9CM|Injury-hunting rifle|Injury-hunting rifle
C0261979|T037|PT|E955.2|ICD9CM|Suicide and self-inflicted injury by hunting rifle|Suicide and self-inflicted injury by hunting rifle
C0261980|T037|AB|E955.3|ICD9CM|Injury-military firearm|Injury-military firearm
C0261980|T037|PT|E955.3|ICD9CM|Suicide and self-inflicted injury by military firearms|Suicide and self-inflicted injury by military firearms
C0261981|T037|AB|E955.4|ICD9CM|Injury-firearm NEC|Injury-firearm NEC
C0261981|T037|PT|E955.4|ICD9CM|Suicide and self-inflicted injury by other and unspecified firearm|Suicide and self-inflicted injury by other and unspecified firearm
C0261982|T037|AB|E955.5|ICD9CM|Injury-explosives|Injury-explosives
C0261982|T037|PT|E955.5|ICD9CM|Suicide and self-inflicted injury by explosives|Suicide and self-inflicted injury by explosives
C0490036|T037|AB|E955.6|ICD9CM|Self inflict acc-air gun|Self inflict acc-air gun
C0490036|T037|PT|E955.6|ICD9CM|Suicide and self-inflicted injury by air gun|Suicide and self-inflicted injury by air gun
C1135315|T037|AB|E955.7|ICD9CM|Self inj-paintball gun|Self inj-paintball gun
C1135315|T037|PT|E955.7|ICD9CM|Suicide and self-inflicted injury by paintball gun|Suicide and self-inflicted injury by paintball gun
C0375754|T037|AB|E955.9|ICD9CM|Injury-firearm/expl NOS|Injury-firearm/expl NOS
C0375754|T037|PT|E955.9|ICD9CM|Suicide and self-inflicted injury by firearms and explosives, unspecified|Suicide and self-inflicted injury by firearms and explosives, unspecified
C0261983|T037|AB|E956|ICD9CM|Injury-cut instrument|Injury-cut instrument
C0261983|T037|PT|E956|ICD9CM|Suicide and self-inflicted injury by cutting and piercing instrument|Suicide and self-inflicted injury by cutting and piercing instrument
C0261984|T037|HT|E957|ICD9CM|Suicide and self-inflicted injuries by jumping from high place|Suicide and self-inflicted injuries by jumping from high place
C0261985|T037|AB|E957.0|ICD9CM|Injury-jump fm residence|Injury-jump fm residence
C0261985|T037|PT|E957.0|ICD9CM|Suicide and self-inflicted injuries by jumping from residential premises|Suicide and self-inflicted injuries by jumping from residential premises
C0546831|T037|AB|E957.1|ICD9CM|Injury-jump fm struc NEC|Injury-jump fm struc NEC
C0546831|T037|PT|E957.1|ICD9CM|Suicide and self-inflicted injuries by jumping from other man-made structures|Suicide and self-inflicted injuries by jumping from other man-made structures
C0261987|T037|AB|E957.2|ICD9CM|Injury-jump fm natur sit|Injury-jump fm natur sit
C0261987|T037|PT|E957.2|ICD9CM|Suicide and self-inflicted injuries by jumping from natural sites|Suicide and self-inflicted injuries by jumping from natural sites
C0261988|T037|AB|E957.9|ICD9CM|Injury-jump NEC|Injury-jump NEC
C0261988|T037|PT|E957.9|ICD9CM|Suicide and self-inflicted injuries by jumping from unspecified site|Suicide and self-inflicted injuries by jumping from unspecified site
C0261989|T037|HT|E958|ICD9CM|Suicide and self-inflicted injury by other and unspecified means|Suicide and self-inflicted injury by other and unspecified means
C0261990|T037|AB|E958.0|ICD9CM|Injury-moving object|Injury-moving object
C0261990|T037|PT|E958.0|ICD9CM|Suicide and self-inflicted injury by jumping or lying before moving object|Suicide and self-inflicted injury by jumping or lying before moving object
C0261991|T037|AB|E958.1|ICD9CM|Injury-burn, fire|Injury-burn, fire
C0261991|T037|PT|E958.1|ICD9CM|Suicide and self-inflicted injury by burns, fire|Suicide and self-inflicted injury by burns, fire
C0261992|T037|AB|E958.2|ICD9CM|Injury-scald|Injury-scald
C0261992|T037|PT|E958.2|ICD9CM|Suicide and self-inflicted injury by scald|Suicide and self-inflicted injury by scald
C0261993|T037|AB|E958.3|ICD9CM|Injury-extreme cold|Injury-extreme cold
C0261993|T037|PT|E958.3|ICD9CM|Suicide and self-inflicted injury by extremes of cold|Suicide and self-inflicted injury by extremes of cold
C0261994|T037|AB|E958.4|ICD9CM|Injury-electrocution|Injury-electrocution
C0261994|T037|PT|E958.4|ICD9CM|Suicide and self-inflicted injury by electrocution|Suicide and self-inflicted injury by electrocution
C0261995|T037|AB|E958.5|ICD9CM|Injury-motor veh crash|Injury-motor veh crash
C0261995|T037|PT|E958.5|ICD9CM|Suicide and self-inflicted injury by crashing of motor vehicle|Suicide and self-inflicted injury by crashing of motor vehicle
C0261996|T037|AB|E958.6|ICD9CM|Injury-aircraft crash|Injury-aircraft crash
C0261996|T037|PT|E958.6|ICD9CM|Suicide and self-inflicted injury by crashing of aircraft|Suicide and self-inflicted injury by crashing of aircraft
C0261997|T037|AB|E958.7|ICD9CM|Injury-caustic substance|Injury-caustic substance
C0261997|T037|PT|E958.7|ICD9CM|Suicide and self-inflicted injury by caustic substances, except poisoning|Suicide and self-inflicted injury by caustic substances, except poisoning
C0261974|T037|AB|E958.8|ICD9CM|Injury-NEC|Injury-NEC
C0261974|T037|PT|E958.8|ICD9CM|Suicide and self-inflicted injury by other specified means|Suicide and self-inflicted injury by other specified means
C0038662|T037|AB|E958.9|ICD9CM|Injury-NOS|Injury-NOS
C0038662|T037|PT|E958.9|ICD9CM|Suicide and self-inflicted injury by unspecified means|Suicide and self-inflicted injury by unspecified means
C0481358|T037|AB|E959|ICD9CM|Late eff of self-injury|Late eff of self-injury
C0481358|T037|PT|E959|ICD9CM|Late effects of self-inflicted injury|Late effects of self-inflicted injury
C0261999|T037|HT|E960|ICD9CM|Fight, brawl, rape|Fight, brawl, rape
C0178361|T033|HT|E960-E969.9|ICD9CM|HOMICIDE AND INJURY PURPOSELY INFLICTED BY OTHER PERSONS|HOMICIDE AND INJURY PURPOSELY INFLICTED BY OTHER PERSONS
C0262001|T037|PT|E961|ICD9CM|Assault by corrosive or caustic substance, except poisoning|Assault by corrosive or caustic substance, except poisoning
C0262001|T037|AB|E961|ICD9CM|Assault-corrosiv/caust|Assault-corrosiv/caust
C0262002|T037|HT|E962|ICD9CM|Assault by poisoning|Assault by poisoning
C0262003|T037|PT|E962.0|ICD9CM|Assault by drugs and medicinal substances|Assault by drugs and medicinal substances
C0262003|T037|AB|E962.0|ICD9CM|Assault-pois w medic agt|Assault-pois w medic agt
C0262004|T037|PT|E962.1|ICD9CM|Assault by other solid and liquid substances|Assault by other solid and liquid substances
C0262004|T037|AB|E962.1|ICD9CM|Assault-pois w solid/liq|Assault-pois w solid/liq
C0262005|T037|PT|E962.2|ICD9CM|Assault by other gases and vapors|Assault by other gases and vapors
C0262005|T037|AB|E962.2|ICD9CM|Assault-pois w gas/vapor|Assault-pois w gas/vapor
C0262002|T037|PT|E962.9|ICD9CM|Assault by unspecified poisoning|Assault by unspecified poisoning
C0262002|T037|AB|E962.9|ICD9CM|Assault-poisoning NOS|Assault-poisoning NOS
C0262007|T037|PT|E963|ICD9CM|Assault by hanging and strangulation|Assault by hanging and strangulation
C0262007|T037|AB|E963|ICD9CM|Assault-hanging/strangul|Assault-hanging/strangul
C0262008|T037|PT|E964|ICD9CM|Assault by submersion [drowning]|Assault by submersion [drowning]
C0262008|T037|AB|E964|ICD9CM|Assault-submersion|Assault-submersion
C0262009|T037|HT|E965|ICD9CM|Assault by firearms and explosives|Assault by firearms and explosives
C0262010|T037|PT|E965.0|ICD9CM|Assault by handgun|Assault by handgun
C0262010|T037|AB|E965.0|ICD9CM|Assault-handgun|Assault-handgun
C0262011|T037|PT|E965.1|ICD9CM|Assault by shotgun|Assault by shotgun
C0262011|T037|AB|E965.1|ICD9CM|Assault-shotgun|Assault-shotgun
C0262012|T037|PT|E965.2|ICD9CM|Assault by hunting rifle|Assault by hunting rifle
C0262012|T037|AB|E965.2|ICD9CM|Assault-hunting rifle|Assault-hunting rifle
C0262013|T037|PT|E965.3|ICD9CM|Assault by military firearms|Assault by military firearms
C0262013|T037|AB|E965.3|ICD9CM|Assault-military weapon|Assault-military weapon
C0480620|T037|PT|E965.4|ICD9CM|Assault by other and unspecified firearm|Assault by other and unspecified firearm
C0480620|T037|AB|E965.4|ICD9CM|Assault-firearm NEC|Assault-firearm NEC
C0262015|T037|PT|E965.5|ICD9CM|Assault by antipersonnel bomb|Assault by antipersonnel bomb
C0262015|T037|AB|E965.5|ICD9CM|Assault-antiperson bomb|Assault-antiperson bomb
C0418380|T037|PT|E965.6|ICD9CM|Assault by gasoline bomb|Assault by gasoline bomb
C0418380|T037|AB|E965.6|ICD9CM|Assault-gasoline bomb|Assault-gasoline bomb
C0262017|T037|PT|E965.7|ICD9CM|Assault by letter bomb|Assault by letter bomb
C0262017|T037|AB|E965.7|ICD9CM|Assault-letter bomb|Assault-letter bomb
C0262018|T037|PT|E965.8|ICD9CM|Assault by other specified explosive|Assault by other specified explosive
C0262018|T037|AB|E965.8|ICD9CM|Assault-explosive NEC|Assault-explosive NEC
C0262019|T037|PT|E965.9|ICD9CM|Assault by unspecified explosive|Assault by unspecified explosive
C0262019|T037|AB|E965.9|ICD9CM|Assault-explosive NOS|Assault-explosive NOS
C0418384|T037|PT|E966|ICD9CM|Assault by cutting and piercing instrument|Assault by cutting and piercing instrument
C0418384|T037|AB|E966|ICD9CM|Assault-cutting instr|Assault-cutting instr
C0878756|T033|HT|E967|ICD9CM|Perpetrator of child and adult abuse|Perpetrator of child and adult abuse
C0878757|T033|AB|E967.0|ICD9CM|Abuse by fther/stpfth/bf|Abuse by fther/stpfth/bf
C0878757|T033|PT|E967.0|ICD9CM|Perpetrator of child and adult abuse, by father, stepfather, or boyfriend|Perpetrator of child and adult abuse, by father, stepfather, or boyfriend
C0262023|T037|AB|E967.1|ICD9CM|Child abuse by pers NEC|Child abuse by pers NEC
C0262023|T037|PT|E967.1|ICD9CM|Perpetrator of child and adult abuse, by other specified person|Perpetrator of child and adult abuse, by other specified person
C0878758|T033|AB|E967.2|ICD9CM|Abuse by mther/stpmth/gf|Abuse by mther/stpmth/gf
C0878758|T033|PT|E967.2|ICD9CM|Perpetrator of child and adult abuse, by mother, stepmother, or girlfriend|Perpetrator of child and adult abuse, by mother, stepmother, or girlfriend
C0375757|T037|AB|E967.3|ICD9CM|Batter by spouse/partner|Batter by spouse/partner
C0375757|T037|PT|E967.3|ICD9CM|Perpetrator of child and adult abuse, by spouse or partner|Perpetrator of child and adult abuse, by spouse or partner
C0375758|T037|AB|E967.4|ICD9CM|Battering by child|Battering by child
C0375758|T037|PT|E967.4|ICD9CM|Perpetrator of child and adult abuse, by child|Perpetrator of child and adult abuse, by child
C0375759|T037|AB|E967.5|ICD9CM|Battering by sibling|Battering by sibling
C0375759|T037|PT|E967.5|ICD9CM|Perpetrator of child and adult abuse, by sibling|Perpetrator of child and adult abuse, by sibling
C0375760|T037|AB|E967.6|ICD9CM|Battering by grandparent|Battering by grandparent
C0375760|T037|PT|E967.6|ICD9CM|Perpetrator of child and adult abuse, by grandparent|Perpetrator of child and adult abuse, by grandparent
C0375761|T037|AB|E967.7|ICD9CM|Batter by other relative|Batter by other relative
C0375761|T037|PT|E967.7|ICD9CM|Perpetrator of child and adult abuse, by other relative|Perpetrator of child and adult abuse, by other relative
C0375762|T037|AB|E967.8|ICD9CM|Batter by non-relative|Batter by non-relative
C0375762|T037|PT|E967.8|ICD9CM|Perpetrator of child and adult abuse, by non-related caregiver|Perpetrator of child and adult abuse, by non-related caregiver
C0375763|T037|AB|E967.9|ICD9CM|Child abuse NOS|Child abuse NOS
C0375763|T037|PT|E967.9|ICD9CM|Perpetrator of child and adult abuse, by unspecified person|Perpetrator of child and adult abuse, by unspecified person
C0262024|T037|HT|E968|ICD9CM|Assault by other and unspecified means|Assault by other and unspecified means
C0262025|T037|PT|E968.0|ICD9CM|Assault by fire|Assault by fire
C0262025|T037|AB|E968.0|ICD9CM|Assault-fire|Assault-fire
C0480686|T037|PT|E968.1|ICD9CM|Assault by pushing from a high place|Assault by pushing from a high place
C0480686|T037|AB|E968.1|ICD9CM|Asslt-push from hi place|Asslt-push from hi place
C0262027|T037|PT|E968.2|ICD9CM|Assault by striking by blunt or thrown object|Assault by striking by blunt or thrown object
C0262027|T037|AB|E968.2|ICD9CM|Assault-striking w obj|Assault-striking w obj
C0262028|T037|PT|E968.3|ICD9CM|Assault by hot liquid|Assault by hot liquid
C0262028|T037|AB|E968.3|ICD9CM|Assault-hot liquid|Assault-hot liquid
C0418343|T033|PT|E968.4|ICD9CM|Assault by criminal neglect|Assault by criminal neglect
C0418343|T033|AB|E968.4|ICD9CM|Assault-criminal neglect|Assault-criminal neglect
C0375764|T037|PT|E968.5|ICD9CM|Assault by transport vehicle|Assault by transport vehicle
C0375764|T037|AB|E968.5|ICD9CM|Asslt-transport vehicle|Asslt-transport vehicle
C0490037|T037|AB|E968.6|ICD9CM|Assault - air gun|Assault - air gun
C0490037|T037|PT|E968.6|ICD9CM|Assault by air gun|Assault by air gun
C0418414|T037|PT|E968.7|ICD9CM|Assault by human bite|Assault by human bite
C0418414|T037|AB|E968.7|ICD9CM|Human bite - assault|Human bite - assault
C0262030|T037|PT|E968.8|ICD9CM|Assault by other specified means|Assault by other specified means
C0262030|T037|AB|E968.8|ICD9CM|Assault NEC|Assault NEC
C0004063|T037|PT|E968.9|ICD9CM|Assault by unspecified means|Assault by unspecified means
C0004063|T037|AB|E968.9|ICD9CM|Assault NOS|Assault NOS
C0418456|T037|AB|E969|ICD9CM|Late effect assault|Late effect assault
C0418456|T037|PT|E969|ICD9CM|Late effects of injury purposely inflicted by other person|Late effects of injury purposely inflicted by other person
C0262032|T037|PT|E970|ICD9CM|Injury due to legal intervention by firearms|Injury due to legal intervention by firearms
C0262032|T037|AB|E970|ICD9CM|Legal intervent-firearm|Legal intervent-firearm
C0178362|T037|HT|E970-E978.9|ICD9CM|LEGAL INTERVENTION|LEGAL INTERVENTION
C0262033|T037|PT|E971|ICD9CM|Injury due to legal intervention by explosives|Injury due to legal intervention by explosives
C0262033|T037|AB|E971|ICD9CM|Legal intervent-explosiv|Legal intervent-explosiv
C0262034|T037|PT|E972|ICD9CM|Injury due to legal intervention by gas|Injury due to legal intervention by gas
C0262034|T037|AB|E972|ICD9CM|Legal intervent-gas|Legal intervent-gas
C0262035|T037|PT|E973|ICD9CM|Injury due to legal intervention by blunt object|Injury due to legal intervention by blunt object
C0262035|T037|AB|E973|ICD9CM|Legal interven-blunt obj|Legal interven-blunt obj
C0418479|T037|PT|E974|ICD9CM|Injury due to legal intervention by cutting and piercing instrument|Injury due to legal intervention by cutting and piercing instrument
C0418479|T037|AB|E974|ICD9CM|Legal interven-cut instr|Legal interven-cut instr
C0262037|T037|PT|E975|ICD9CM|Injury due to legal intervention by other specified means|Injury due to legal intervention by other specified means
C0262037|T037|AB|E975|ICD9CM|Legal intervention NEC|Legal intervention NEC
C0262038|T037|PT|E976|ICD9CM|Injury due to legal intervention by unspecified means|Injury due to legal intervention by unspecified means
C0262038|T037|AB|E976|ICD9CM|Legal intervention NOS|Legal intervention NOS
C0481367|T037|AB|E977|ICD9CM|Late eff-legal intervent|Late eff-legal intervent
C0481367|T037|PT|E977|ICD9CM|Late effects of injuries due to legal intervention|Late effects of injuries due to legal intervention
C2077104|T037|HT|E979|ICD9CM|Terrorism|Terrorism
C2077104|T037|HT|E979-E979.9|ICD9CM|TERRORISM|TERRORISM
C1135316|T037|PT|E979.0|ICD9CM|Terrorism involving explosion of marine weapons|Terrorism involving explosion of marine weapons
C1135316|T037|AB|E979.0|ICD9CM|Terrorism,marine weapons|Terrorism,marine weapons
C1135317|T037|PT|E979.1|ICD9CM|Terrorism involving destruction of aircraft|Terrorism involving destruction of aircraft
C1135317|T037|AB|E979.1|ICD9CM|Terrorism,dest aircraft|Terrorism,dest aircraft
C1135318|T037|PT|E979.2|ICD9CM|Terrorism involving other explosions and fragments|Terrorism involving other explosions and fragments
C1135318|T037|AB|E979.2|ICD9CM|Terrorism,explosions|Terrorism,explosions
C1135319|T037|PT|E979.3|ICD9CM|Terrorism involving fires|Terrorism involving fires
C1135319|T037|AB|E979.3|ICD9CM|Terrorism, fires|Terrorism, fires
C1135320|T037|PT|E979.4|ICD9CM|Terrorism involving firearms|Terrorism involving firearms
C1135320|T037|AB|E979.4|ICD9CM|Terrorism, firearms|Terrorism, firearms
C1135321|T037|PT|E979.5|ICD9CM|Terrorism involving nuclear weapons|Terrorism involving nuclear weapons
C1135321|T037|AB|E979.5|ICD9CM|Terrorism, nuc weapons|Terrorism, nuc weapons
C1135322|T037|PT|E979.6|ICD9CM|Terrorism involving biological weapons|Terrorism involving biological weapons
C1135322|T037|AB|E979.6|ICD9CM|Terrorism, biologicals|Terrorism, biologicals
C1135323|T037|PT|E979.7|ICD9CM|Terrorism involving chemical weapons|Terrorism involving chemical weapons
C1135323|T037|AB|E979.7|ICD9CM|Terrorism, chemicals|Terrorism, chemicals
C1135324|T037|PT|E979.8|ICD9CM|Terrorism involving other means|Terrorism involving other means
C1135324|T037|AB|E979.8|ICD9CM|Terrorism, NEC/NOS|Terrorism, NEC/NOS
C1135325|T037|PT|E979.9|ICD9CM|Terrorism secondary effects|Terrorism secondary effects
C1135325|T037|AB|E979.9|ICD9CM|Terrorism, secondary|Terrorism, secondary
C0262040|T037|HT|E980|ICD9CM|Poisoning by solid or liquid substances, undetermined whether accidentally or purposely inflicted|Poisoning by solid or liquid substances, undetermined whether accidentally or purposely inflicted
C0178363|T037|HT|E980-E989.9|ICD9CM|INJURY UNDETERMINED WHETHER ACCIDENTALLY OR PURPOSELY INFLICTED|INJURY UNDETERMINED WHETHER ACCIDENTALLY OR PURPOSELY INFLICTED
C0262041|T037|AB|E980.0|ICD9CM|Undeterm pois-analgesics|Undeterm pois-analgesics
C0262042|T037|PT|E980.1|ICD9CM|Poisoning by barbiturates, undetermined whether accidentally or purposely inflicted|Poisoning by barbiturates, undetermined whether accidentally or purposely inflicted
C0262042|T037|AB|E980.1|ICD9CM|Undeterm pois-barbiturat|Undeterm pois-barbiturat
C0262043|T037|PT|E980.2|ICD9CM|Poisoning by other sedatives and hypnotics, undetermined whether accidentally or purposely inflicted|Poisoning by other sedatives and hypnotics, undetermined whether accidentally or purposely inflicted
C0262043|T037|AB|E980.2|ICD9CM|Undet pois-sed/hypn NEC|Undet pois-sed/hypn NEC
C0262044|T037|AB|E980.3|ICD9CM|Undeterm pois-psychotrop|Undeterm pois-psychotrop
C0262045|T037|AB|E980.4|ICD9CM|Undet pois-med agnt NEC|Undet pois-med agnt NEC
C0262046|T037|AB|E980.5|ICD9CM|Undet pois-med agnt NOS|Undet pois-med agnt NOS
C0262047|T037|AB|E980.6|ICD9CM|Undet pois-corros/caust|Undet pois-corros/caust
C0262048|T037|AB|E980.7|ICD9CM|Undet pois-agricult agnt|Undet pois-agricult agnt
C0262049|T037|PT|E980.8|ICD9CM|Poisoning by arsenic and its compounds, undetermined whether accidentally or purposely inflicted|Poisoning by arsenic and its compounds, undetermined whether accidentally or purposely inflicted
C0262049|T037|AB|E980.8|ICD9CM|Undeter pois-arsenic|Undeter pois-arsenic
C0262050|T037|AB|E980.9|ICD9CM|Undeter pois-sol/liq NEC|Undeter pois-sol/liq NEC
C0262051|T037|HT|E981|ICD9CM|Poisoning by gases in domestic use, undetermined whether accidentally or purposely inflicted|Poisoning by gases in domestic use, undetermined whether accidentally or purposely inflicted
C0262052|T037|PT|E981.0|ICD9CM|Poisoning by gas distributed by pipeline, undetermined whether accidentally or purposely inflicted|Poisoning by gas distributed by pipeline, undetermined whether accidentally or purposely inflicted
C0262052|T037|AB|E981.0|ICD9CM|Undeter pois-piped gas|Undeter pois-piped gas
C0262053|T037|AB|E981.1|ICD9CM|Undet pois-container gas|Undet pois-container gas
C0262054|T037|PT|E981.8|ICD9CM|Poisoning by other utility gas, undetermined whether accidentally or purposely inflicted|Poisoning by other utility gas, undetermined whether accidentally or purposely inflicted
C0262054|T037|AB|E981.8|ICD9CM|Undet pois-util gas NEC|Undet pois-util gas NEC
C0262055|T037|HT|E982|ICD9CM|Poisoning by other gases, undetermined whether accidentally or purposely inflicted|Poisoning by other gases, undetermined whether accidentally or purposely inflicted
C0262056|T037|PT|E982.0|ICD9CM|Poisoning by motor vehicle exhaust gas, undetermined whether accidentally or purposely inflicted|Poisoning by motor vehicle exhaust gas, undetermined whether accidentally or purposely inflicted
C0262056|T037|AB|E982.0|ICD9CM|Undeter pois-exhaust gas|Undeter pois-exhaust gas
C0262057|T037|PT|E982.1|ICD9CM|Poisoning by other carbon monoxide, undetermined whether accidentally or purposely inflicted|Poisoning by other carbon monoxide, undetermined whether accidentally or purposely inflicted
C0262057|T037|AB|E982.1|ICD9CM|Undetermin poison-co NEC|Undetermin poison-co NEC
C0262058|T037|AB|E982.8|ICD9CM|Undet pois-gas/vapor NEC|Undet pois-gas/vapor NEC
C0262059|T037|PT|E982.9|ICD9CM|Poisoning by unspecified gases and vapors, undetermined whether accidentally or purposely inflicted|Poisoning by unspecified gases and vapors, undetermined whether accidentally or purposely inflicted
C0262059|T037|AB|E982.9|ICD9CM|Undet pois-gas/vapor NOS|Undet pois-gas/vapor NOS
C0262060|T037|HT|E983|ICD9CM|Hanging, strangulation, or suffocation, undetermined whether accidentally or purposely inflicted|Hanging, strangulation, or suffocation, undetermined whether accidentally or purposely inflicted
C0262061|T037|PT|E983.0|ICD9CM|Hanging, undetermined whether accidentally or purposely inflicted|Hanging, undetermined whether accidentally or purposely inflicted
C0262061|T037|AB|E983.0|ICD9CM|Undetermin circ-hanging|Undetermin circ-hanging
C0262062|T037|PT|E983.1|ICD9CM|Suffocation by plastic bag, undetermined whether accidentally or purposely inflicted|Suffocation by plastic bag, undetermined whether accidentally or purposely inflicted
C0262062|T037|AB|E983.1|ICD9CM|Undet circ-suf plast bag|Undet circ-suf plast bag
C0262063|T037|AB|E983.8|ICD9CM|Undet circ-suffocate NEC|Undet circ-suffocate NEC
C0262064|T037|AB|E983.9|ICD9CM|Undet circ-suffocate NOS|Undet circ-suffocate NOS
C0262065|T037|PT|E984|ICD9CM|Submersion (drowning), undetermined whether accidentally or purposely inflicted|Submersion (drowning), undetermined whether accidentally or purposely inflicted
C0262065|T037|AB|E984|ICD9CM|Undeterm circ-submersion|Undeterm circ-submersion
C0262067|T037|PT|E985.0|ICD9CM|Injury by handgun, undetermined whether accidentally or purposely inflicted|Injury by handgun, undetermined whether accidentally or purposely inflicted
C0262067|T037|AB|E985.0|ICD9CM|Undetermin circ-handgun|Undetermin circ-handgun
C0262068|T037|PT|E985.1|ICD9CM|Injury by shotgun, undetermined whether accidentally or purposely inflicted|Injury by shotgun, undetermined whether accidentally or purposely inflicted
C0262068|T037|AB|E985.1|ICD9CM|Undetermin circ-shotgun|Undetermin circ-shotgun
C0262069|T037|PT|E985.2|ICD9CM|Injury by hunting rifle, undetermined whether accidentally or purposely inflicted|Injury by hunting rifle, undetermined whether accidentally or purposely inflicted
C0262069|T037|AB|E985.2|ICD9CM|Undet circ-hunting rifle|Undet circ-hunting rifle
C0262070|T037|PT|E985.3|ICD9CM|Injury by military firearms, undetermined whether accidentally or purposely inflicted|Injury by military firearms, undetermined whether accidentally or purposely inflicted
C0262070|T037|AB|E985.3|ICD9CM|Undet circ-military arms|Undet circ-military arms
C0262071|T037|PT|E985.4|ICD9CM|Injury by other and unspecified firearm, undetermined whether accidentally or purposely inflicted|Injury by other and unspecified firearm, undetermined whether accidentally or purposely inflicted
C0262071|T037|AB|E985.4|ICD9CM|Undeter circ-firearm NEC|Undeter circ-firearm NEC
C0262072|T037|PT|E985.5|ICD9CM|Injury by explosives, undetermined whether accidentally or purposely inflicted|Injury by explosives, undetermined whether accidentally or purposely inflicted
C0262072|T037|AB|E985.5|ICD9CM|Undeterm circ-explosive|Undeterm circ-explosive
C0490038|T037|PT|E985.6|ICD9CM|Injury by air gun, undetermined whether accidental or purposely inflicted|Injury by air gun, undetermined whether accidental or purposely inflicted
C0490038|T037|AB|E985.6|ICD9CM|Undetrmine accid-air gun|Undetrmine accid-air gun
C1135326|T037|PT|E985.7|ICD9CM|Injury by paintball gun, undetermined whether accidental or purposely inflicted|Injury by paintball gun, undetermined whether accidental or purposely inflicted
C1135326|T037|AB|E985.7|ICD9CM|Injury paintball gun NOS|Injury paintball gun NOS
C0262073|T037|PT|E986|ICD9CM|Injury by cutting and piercing instruments, undetermined whether accidentally or purposely inflicted|Injury by cutting and piercing instruments, undetermined whether accidentally or purposely inflicted
C0262073|T037|AB|E986|ICD9CM|Undet circ-cut instrumnt|Undet circ-cut instrumnt
C0262075|T037|PT|E987.0|ICD9CM|Falling from residential premises, undetermined whether accidentally or purposely inflicted|Falling from residential premises, undetermined whether accidentally or purposely inflicted
C0262075|T037|AB|E987.0|ICD9CM|Undet circ-fall residenc|Undet circ-fall residenc
C0262088|T037|HT|E988|ICD9CM|Injury by other and unspecified means, undetermined whether accidentally or purposely inflicted|Injury by other and unspecified means, undetermined whether accidentally or purposely inflicted
C0262080|T037|AB|E988.0|ICD9CM|Undeterm circ-moving obj|Undeterm circ-moving obj
C0262081|T037|PT|E988.1|ICD9CM|Injury by burns or fire, undetermined whether accidentally or purposely inflicted|Injury by burns or fire, undetermined whether accidentally or purposely inflicted
C0262081|T037|AB|E988.1|ICD9CM|Undeterm circ-burn, fire|Undeterm circ-burn, fire
C0332691|T037|PT|E988.2|ICD9CM|Injury by scald, undetermined whether accidentally or purposely inflicted|Injury by scald, undetermined whether accidentally or purposely inflicted
C0332691|T037|AB|E988.2|ICD9CM|Undeterm circ-scald|Undeterm circ-scald
C0262083|T037|PT|E988.3|ICD9CM|Injury by extremes of cold, undetermined whether accidentally or purposely inflicted|Injury by extremes of cold, undetermined whether accidentally or purposely inflicted
C0262083|T037|AB|E988.3|ICD9CM|Undeterm circ-extrm cold|Undeterm circ-extrm cold
C0262084|T037|PT|E988.4|ICD9CM|Injury by electrocution, undetermined whether accidentally or purposely inflicted|Injury by electrocution, undetermined whether accidentally or purposely inflicted
C0262084|T037|AB|E988.4|ICD9CM|Undeterm circ-electrocut|Undeterm circ-electrocut
C0262085|T037|PT|E988.5|ICD9CM|Injury by crashing of motor vehicle, undetermined whether accidentally or purposely inflicted|Injury by crashing of motor vehicle, undetermined whether accidentally or purposely inflicted
C0262085|T037|AB|E988.5|ICD9CM|Undet circ-mot veh crash|Undet circ-mot veh crash
C0262086|T037|PT|E988.6|ICD9CM|Injury by crashing of aircraft, undetermined whether accidentally or purposely inflicted|Injury by crashing of aircraft, undetermined whether accidentally or purposely inflicted
C0262086|T037|AB|E988.6|ICD9CM|Undet circ-aircrft crash|Undet circ-aircrft crash
C0262087|T037|AB|E988.7|ICD9CM|Undet circ-caustic subst|Undet circ-caustic subst
C0262088|T037|PT|E988.8|ICD9CM|Injury by other specified means, undetermined whether accidentally or purposely inflicted|Injury by other specified means, undetermined whether accidentally or purposely inflicted
C0262088|T037|AB|E988.8|ICD9CM|Undetermin circumst NEC|Undetermin circumst NEC
C0262089|T037|PT|E988.9|ICD9CM|Injury by unspecified means, undetermined whether accidentally or purposely inflicted|Injury by unspecified means, undetermined whether accidentally or purposely inflicted
C0262089|T037|AB|E988.9|ICD9CM|Undetermin circumst NOS|Undetermin circumst NOS
C0481360|T037|AB|E989|ICD9CM|Late eff inj-undet circ|Late eff inj-undet circ
C0481360|T037|PT|E989|ICD9CM|Late effects of injury, undetermined whether accidentally or purposely inflicted|Late effects of injury, undetermined whether accidentally or purposely inflicted
C0262091|T037|HT|E990|ICD9CM|Injury due to war operations by fires and conflagrations|Injury due to war operations by fires and conflagrations
C0178364|T037|HT|E990-E999.9|ICD9CM|INJURY RESULTING FROM OPERATIONS OF WAR|INJURY RESULTING FROM OPERATIONS OF WAR
C0262092|T037|PT|E990.0|ICD9CM|Injury due to war operations from gasoline bomb|Injury due to war operations from gasoline bomb
C0262092|T037|AB|E990.0|ICD9CM|War inj:gasoline bomb|War inj:gasoline bomb
C2712482|T037|PT|E990.1|ICD9CM|Injury due to war operations from flamethrower|Injury due to war operations from flamethrower
C2712482|T037|AB|E990.1|ICD9CM|War inj:flamethrower|War inj:flamethrower
C2712483|T037|PT|E990.2|ICD9CM|Injury due to war operations from incendiary bullet|Injury due to war operations from incendiary bullet
C2712483|T037|AB|E990.2|ICD9CM|War inj:incndiary bullet|War inj:incndiary bullet
C2712484|T037|PT|E990.3|ICD9CM|Injury due to war operations from fire caused indirectly from conventional weapon|Injury due to war operations from fire caused indirectly from conventional weapon
C2712484|T037|AB|E990.3|ICD9CM|War inj:ind convn weapn|War inj:ind convn weapn
C0262093|T037|PT|E990.9|ICD9CM|Injury due to war operations from other and unspecified source|Injury due to war operations from other and unspecified source
C0262093|T037|AB|E990.9|ICD9CM|War injury:fire NEC|War injury:fire NEC
C0262094|T037|HT|E991|ICD9CM|Injury due to war operations by bullets and fragments|Injury due to war operations by bullets and fragments
C0262095|T037|PT|E991.0|ICD9CM|Injury due to war operations from rubber bullets (rifle)|Injury due to war operations from rubber bullets (rifle)
C0262095|T037|AB|E991.0|ICD9CM|War inj:rubber bullet|War inj:rubber bullet
C0262096|T037|PT|E991.1|ICD9CM|Injury due to war operations from pellets (rifle)|Injury due to war operations from pellets (rifle)
C0262096|T037|AB|E991.1|ICD9CM|War injury:pellets|War injury:pellets
C0262097|T037|PT|E991.2|ICD9CM|Injury due to war operations from other bullets|Injury due to war operations from other bullets
C0262097|T037|AB|E991.2|ICD9CM|War injury:bullet NEC|War injury:bullet NEC
C0262098|T037|PT|E991.3|ICD9CM|Injury due to war operations from antipersonnel bomb (fragments)|Injury due to war operations from antipersonnel bomb (fragments)
C0262098|T037|AB|E991.3|ICD9CM|War inj:antiperson bomb|War inj:antiperson bomb
C2712485|T037|PT|E991.4|ICD9CM|Injury due to war operations by fragments from munitions|Injury due to war operations by fragments from munitions
C2712485|T037|AB|E991.4|ICD9CM|War inj:munition fragmnt|War inj:munition fragmnt
C2712486|T037|PT|E991.5|ICD9CM|Injury due to war operations by fragments from person-borne improvised explosive device [IED]|Injury due to war operations by fragments from person-borne improvised explosive device [IED]
C2712486|T037|AB|E991.5|ICD9CM|War inj:prsn-brn fragmnt|War inj:prsn-brn fragmnt
C2712487|T037|PT|E991.6|ICD9CM|Injury due to war operations by fragments from vehicle-borne improvised explosive device [IED]|Injury due to war operations by fragments from vehicle-borne improvised explosive device [IED]
C2712487|T037|AB|E991.6|ICD9CM|War inj:vehic-borne IED|War inj:vehic-borne IED
C2712488|T037|PT|E991.7|ICD9CM|Injury due to war operations by fragments from other improvised explosive device [IED]|Injury due to war operations by fragments from other improvised explosive device [IED]
C2712488|T037|AB|E991.7|ICD9CM|War inj:fragment IED NEC|War inj:fragment IED NEC
C2712489|T037|PT|E991.8|ICD9CM|Injury due to war operations by fragments from weapons|Injury due to war operations by fragments from weapons
C2712489|T037|AB|E991.8|ICD9CM|War inj:weapon fragments|War inj:weapon fragments
C0262099|T037|PT|E991.9|ICD9CM|Injury due to war operations from other and unspecified fragments|Injury due to war operations from other and unspecified fragments
C0262099|T037|AB|E991.9|ICD9CM|War inj:fragments NEC|War inj:fragments NEC
C0262100|T037|HT|E992|ICD9CM|Injury due to war operations by explosion of marine weapons|Injury due to war operations by explosion of marine weapons
C2712490|T037|PT|E992.0|ICD9CM|Injury due to torpedo|Injury due to torpedo
C2712490|T037|AB|E992.0|ICD9CM|War inj:torpedo|War inj:torpedo
C2712491|T037|PT|E992.1|ICD9CM|Injury due to depth charge|Injury due to depth charge
C2712491|T037|AB|E992.1|ICD9CM|War inj:depth charge|War inj:depth charge
C2712492|T037|PT|E992.2|ICD9CM|Injury due to marine mines|Injury due to marine mines
C2712492|T037|AB|E992.2|ICD9CM|War inj:marine mines|War inj:marine mines
C2712493|T037|PT|E992.3|ICD9CM|Injury due to sea-based artillery shell|Injury due to sea-based artillery shell
C2712493|T037|AB|E992.3|ICD9CM|War inj:seabase art shel|War inj:seabase art shel
C2712494|T037|PT|E992.8|ICD9CM|Injury due to war operations by other marine weapons|Injury due to war operations by other marine weapons
C2712494|T037|AB|E992.8|ICD9CM|War inj:marine weapn NEC|War inj:marine weapn NEC
C2712495|T037|PT|E992.9|ICD9CM|Injury due to war operations by unspecified marine weapon|Injury due to war operations by unspecified marine weapon
C2712495|T037|AB|E992.9|ICD9CM|War inj:marine weapn NOS|War inj:marine weapn NOS
C0262101|T037|HT|E993|ICD9CM|Injury due to war operations by other explosion|Injury due to war operations by other explosion
C2712496|T037|PT|E993.0|ICD9CM|Injury due to war operations by aerial bomb|Injury due to war operations by aerial bomb
C2712496|T037|AB|E993.0|ICD9CM|War inj:aerial bomb|War inj:aerial bomb
C2712497|T037|PT|E993.1|ICD9CM|Injury due to war operations by guided missile|Injury due to war operations by guided missile
C2712497|T037|AB|E993.1|ICD9CM|War inj:guided missile|War inj:guided missile
C2712498|T037|PT|E993.2|ICD9CM|Injury due to war operations by mortar|Injury due to war operations by mortar
C2712498|T037|AB|E993.2|ICD9CM|War inj:mortar|War inj:mortar
C2712499|T037|PT|E993.3|ICD9CM|Injury due to war operations by person-borne improvised explosive device [IED]|Injury due to war operations by person-borne improvised explosive device [IED]
C2712499|T037|AB|E993.3|ICD9CM|War inj:person IED|War inj:person IED
C2712500|T037|PT|E993.4|ICD9CM|Injury due to war operations by vehicle-borne improvised explosive device [IED]|Injury due to war operations by vehicle-borne improvised explosive device [IED]
C2712500|T037|AB|E993.4|ICD9CM|War inj:vehicle IED|War inj:vehicle IED
C2712501|T037|PT|E993.5|ICD9CM|Injury due to war operations by other improvised explosive device [IED]|Injury due to war operations by other improvised explosive device [IED]
C2712501|T037|AB|E993.5|ICD9CM|War inj:IED NEC|War inj:IED NEC
C2712502|T037|PT|E993.6|ICD9CM|Injury due to war operations by unintentional detonation of own munitions|Injury due to war operations by unintentional detonation of own munitions
C2712502|T037|AB|E993.6|ICD9CM|War inj:acc own munition|War inj:acc own munition
C2712503|T037|PT|E993.7|ICD9CM|Injury due to war operations by unintentional discharge of own munitions launch device|Injury due to war operations by unintentional discharge of own munitions launch device
C2712503|T037|AB|E993.7|ICD9CM|War inj:acc disch launch|War inj:acc disch launch
C2712504|T037|PT|E993.8|ICD9CM|Injury due to war operations by other specified explosion|Injury due to war operations by other specified explosion
C2712504|T037|AB|E993.8|ICD9CM|War inj:explosion NEC|War inj:explosion NEC
C0418717|T037|PT|E993.9|ICD9CM|Injury due to war operations by unspecified explosion|Injury due to war operations by unspecified explosion
C0418717|T037|AB|E993.9|ICD9CM|War inj:explosion NOS|War inj:explosion NOS
C0262102|T037|HT|E994|ICD9CM|Injury due to war operations by destruction of aircraft|Injury due to war operations by destruction of aircraft
C2712505|T037|PT|E994.0|ICD9CM|Injury due to war operations by destruction of aircraft due to enemy fire or explosives|Injury due to war operations by destruction of aircraft due to enemy fire or explosives
C2712505|T037|AB|E994.0|ICD9CM|War inj:aircrft des-enmy|War inj:aircrft des-enmy
C2712506|T037|PT|E994.1|ICD9CM|Injury due to war operations by unintentional destruction of aircraft due to own onboard explosives|Injury due to war operations by unintentional destruction of aircraft due to own onboard explosives
C2712506|T037|AB|E994.1|ICD9CM|War inj:aircrft-own expl|War inj:aircrft-own expl
C2712507|T037|PT|E994.2|ICD9CM|Injury due to war operations by destruction of aircraft due to collision with other aircraft|Injury due to war operations by destruction of aircraft due to collision with other aircraft
C2712507|T037|AB|E994.2|ICD9CM|War inj:aircrft collisn|War inj:aircrft collisn
C2712508|T037|PT|E994.3|ICD9CM|Injury due to war operations by destruction of aircraft due to onboard fire|Injury due to war operations by destruction of aircraft due to onboard fire
C2712508|T037|AB|E994.3|ICD9CM|War inj:aircraft fire|War inj:aircraft fire
C2712509|T037|PT|E994.8|ICD9CM|Injury due to war operations by other destruction of aircraft|Injury due to war operations by other destruction of aircraft
C2712509|T037|AB|E994.8|ICD9CM|War inj:aircrft dest NEC|War inj:aircrft dest NEC
C2712510|T037|PT|E994.9|ICD9CM|Injury due to war operations by unspecified destruction of aircraft|Injury due to war operations by unspecified destruction of aircraft
C2712510|T037|AB|E994.9|ICD9CM|War inj:aircrft dest NOS|War inj:aircrft dest NOS
C0262103|T037|HT|E995|ICD9CM|Injury due to war operations by other and unspecified forms of conventional warfare|Injury due to war operations by other and unspecified forms of conventional warfare
C2712511|T037|PT|E995.0|ICD9CM|Injury due to war operations by unarmed hand-to-hand combat|Injury due to war operations by unarmed hand-to-hand combat
C2712511|T037|AB|E995.0|ICD9CM|War inj:hnd-hnd combat|War inj:hnd-hnd combat
C2712512|T037|PT|E995.1|ICD9CM|Injury due to war operations, struck by blunt object|Injury due to war operations, struck by blunt object
C2712512|T037|AB|E995.1|ICD9CM|War inj:blunt object|War inj:blunt object
C2712513|T037|PT|E995.2|ICD9CM|Injury due to war operations by piercing object|Injury due to war operations by piercing object
C2712513|T037|AB|E995.2|ICD9CM|War inj:piercing object|War inj:piercing object
C2712514|T037|PT|E995.3|ICD9CM|Injury due to war operations by intentional restriction of air and airway|Injury due to war operations by intentional restriction of air and airway
C2712514|T037|AB|E995.3|ICD9CM|War inj:intn restrct air|War inj:intn restrct air
C2712515|T037|PT|E995.4|ICD9CM|Injury due to war operations by unintentional drowning due to inability to surface or obtain air|Injury due to war operations by unintentional drowning due to inability to surface or obtain air
C2712515|T037|AB|E995.4|ICD9CM|War inj:unintentl drown|War inj:unintentl drown
C2712516|T037|PT|E995.8|ICD9CM|Injury due to war operations by other forms of conventional warfare|Injury due to war operations by other forms of conventional warfare
C2712516|T037|AB|E995.8|ICD9CM|War inj:con warfare NEC|War inj:con warfare NEC
C2712517|T037|PT|E995.9|ICD9CM|Injury due to war operations by unspecified form of conventional warfare|Injury due to war operations by unspecified form of conventional warfare
C2712517|T037|AB|E995.9|ICD9CM|War inj:con warfare NOS|War inj:con warfare NOS
C0418710|T037|HT|E996|ICD9CM|Injury due to war operations by nuclear weapons|Injury due to war operations by nuclear weapons
C2712518|T037|PT|E996.0|ICD9CM|Injury due to war operations by direct blast effect of nuclear weapon|Injury due to war operations by direct blast effect of nuclear weapon
C2712518|T037|AB|E996.0|ICD9CM|War inj:dir nucl weapon|War inj:dir nucl weapon
C2712519|T037|PT|E996.1|ICD9CM|Injury due to war operations by indirect blast effect of nuclear weapon|Injury due to war operations by indirect blast effect of nuclear weapon
C2712519|T037|AB|E996.1|ICD9CM|War inj:indir nucl weapn|War inj:indir nucl weapn
C2712520|T037|PT|E996.2|ICD9CM|Injury due to war operations by thermal radiation effect of nuclear weapon|Injury due to war operations by thermal radiation effect of nuclear weapon
C2712520|T037|AB|E996.2|ICD9CM|War inj:therml radiation|War inj:therml radiation
C2712521|T037|PT|E996.3|ICD9CM|Injury due to war operations by nuclear radiation effects|Injury due to war operations by nuclear radiation effects
C2712521|T037|AB|E996.3|ICD9CM|War inj:nuclear rad eff|War inj:nuclear rad eff
C2712522|T037|PT|E996.8|ICD9CM|Injury due to war operations by other effects of nuclear weapons|Injury due to war operations by other effects of nuclear weapons
C2712522|T037|AB|E996.8|ICD9CM|War inj:nucl weapon NEC|War inj:nucl weapon NEC
C2712523|T037|PT|E996.9|ICD9CM|Injury due to war operations by unspecified effect of nuclear weapon|Injury due to war operations by unspecified effect of nuclear weapon
C2712523|T037|AB|E996.9|ICD9CM|War inj:nucl weapon NOS|War inj:nucl weapon NOS
C0262105|T037|HT|E997|ICD9CM|Injury due to war operations by other forms of unconventional warfare|Injury due to war operations by other forms of unconventional warfare
C0262106|T037|PT|E997.0|ICD9CM|Injury due to war operations by lasers|Injury due to war operations by lasers
C0262106|T037|AB|E997.0|ICD9CM|War injury:lasers|War injury:lasers
C0262107|T037|PT|E997.1|ICD9CM|Injury due to war operations by biological warfare|Injury due to war operations by biological warfare
C0262107|T037|AB|E997.1|ICD9CM|War injury:biol warfare|War injury:biol warfare
C0262108|T037|PT|E997.2|ICD9CM|Injury due to war operations by gases, fumes, and chemicals|Injury due to war operations by gases, fumes, and chemicals
C0262108|T037|AB|E997.2|ICD9CM|War injury:gas/fum/chem|War injury:gas/fum/chem
C2712524|T037|PT|E997.3|ICD9CM|Injury due to war operations by weapon of mass destruction [WMD], unspecified|Injury due to war operations by weapon of mass destruction [WMD], unspecified
C2712524|T037|AB|E997.3|ICD9CM|War inj:WMD NOS|War inj:WMD NOS
C0262109|T037|PT|E997.8|ICD9CM|Injury due to other specified forms of unconventional warfare|Injury due to other specified forms of unconventional warfare
C0262109|T037|AB|E997.8|ICD9CM|War inj-unconven war NEC|War inj-unconven war NEC
C0262110|T037|PT|E997.9|ICD9CM|Injury due to unspecified form of unconventional warfare|Injury due to unspecified form of unconventional warfare
C0262110|T037|AB|E997.9|ICD9CM|War inj-unconven war NOS|War inj-unconven war NOS
C0262111|T037|HT|E998|ICD9CM|Injury due to war operations but occurring after cessation of hostilities|Injury due to war operations but occurring after cessation of hostilities
C2712525|T037|PT|E998.0|ICD9CM|Injury due to war operations but occurring after cessation of hostilities by explosion of mines|Injury due to war operations but occurring after cessation of hostilities by explosion of mines
C2712525|T037|AB|E998.0|ICD9CM|War inj:expl mine-cease|War inj:expl mine-cease
C2712526|T037|PT|E998.1|ICD9CM|Injury due to war operations but occurring after cessation of hostilities by explosion of bombs|Injury due to war operations but occurring after cessation of hostilities by explosion of bombs
C2712526|T037|AB|E998.1|ICD9CM|War inj:expl bomb-cease|War inj:expl bomb-cease
C2712527|T037|PT|E998.8|ICD9CM|Injury due to other war operations but occurring after cessation of hostilities|Injury due to other war operations but occurring after cessation of hostilities
C2712527|T037|AB|E998.8|ICD9CM|War inj:after cease NEC|War inj:after cease NEC
C2712528|T037|PT|E998.9|ICD9CM|Injury due to unspecified war operations but occurring after cessation of hostilities|Injury due to unspecified war operations but occurring after cessation of hostilities
C2712528|T037|AB|E998.9|ICD9CM|War inj:after cease NOS|War inj:after cease NOS
C1135340|T037|HT|E999|ICD9CM|Late effect of injury due to war operations and terrorism|Late effect of injury due to war operations and terrorism
C0481368|T046|PT|E999.0|ICD9CM|Late effect of injury due to war operations|Late effect of injury due to war operations
C0481368|T046|AB|E999.0|ICD9CM|Late effect, war injury|Late effect, war injury
C1135327|T046|PT|E999.1|ICD9CM|Late effect of injury due to terrorism|Late effect of injury due to terrorism
C1135327|T046|AB|E999.1|ICD9CM|Late effect, terrorism|Late effect, terrorism
C0260339|T033|HT|V01|ICD9CM|Contact with or exposure to communicable diseases|Contact with or exposure to communicable diseases
C0178337|T033|HT|V01-V06.99|ICD9CM|PERSONS WITH POTENTIAL HEALTH HAZARDS RELATED TO COMMUNICABLE DISEASES|PERSONS WITH POTENTIAL HEALTH HAZARDS RELATED TO COMMUNICABLE DISEASES
C0260340|T033|AB|V01.0|ICD9CM|Cholera contact|Cholera contact
C0260340|T033|PT|V01.0|ICD9CM|Contact with or exposure to cholera|Contact with or exposure to cholera
C0260341|T033|PT|V01.1|ICD9CM|Contact with or exposure to tuberculosis|Contact with or exposure to tuberculosis
C0260341|T033|AB|V01.1|ICD9CM|Tuberculosis contact|Tuberculosis contact
C0260342|T033|PT|V01.2|ICD9CM|Contact with or exposure to poliomyelitis|Contact with or exposure to poliomyelitis
C0260342|T033|AB|V01.2|ICD9CM|Poliomyelitis contact|Poliomyelitis contact
C0260343|T033|PT|V01.3|ICD9CM|Contact with or exposure to smallpox|Contact with or exposure to smallpox
C0260343|T033|AB|V01.3|ICD9CM|Smallpox contact|Smallpox contact
C0260344|T033|PT|V01.4|ICD9CM|Contact with or exposure to rubella|Contact with or exposure to rubella
C0260344|T033|AB|V01.4|ICD9CM|Rubella contact|Rubella contact
C0260345|T033|PT|V01.5|ICD9CM|Contact with or exposure to rabies|Contact with or exposure to rabies
C0260345|T033|AB|V01.5|ICD9CM|Rabies contact|Rabies contact
C0260346|T033|PT|V01.6|ICD9CM|Contact with or exposure to venereal diseases|Contact with or exposure to venereal diseases
C0260346|T033|AB|V01.6|ICD9CM|Venereal dis contact|Venereal dis contact
C0260347|T033|HT|V01.7|ICD9CM|Contact with or exposure to other viral diseases|Contact with or exposure to other viral diseases
C1455968|T033|PT|V01.71|ICD9CM|Contact with or exposure to varicella|Contact with or exposure to varicella
C1455968|T033|AB|V01.71|ICD9CM|Varicella contact/exp|Varicella contact/exp
C0260347|T033|PT|V01.79|ICD9CM|Contact with or exposure to other viral diseases|Contact with or exposure to other viral diseases
C0260347|T033|AB|V01.79|ICD9CM|Viral dis contact NEC|Viral dis contact NEC
C0260348|T033|HT|V01.8|ICD9CM|Contact with or exposure to other communicable diseases|Contact with or exposure to other communicable diseases
C1135271|T033|PT|V01.81|ICD9CM|Contact with or exposure to anthrax|Contact with or exposure to anthrax
C1135271|T033|AB|V01.81|ICD9CM|Contact/exposure-anthrax|Contact/exposure-anthrax
C1260451|T033|AB|V01.82|ICD9CM|Exposure to SARS|Exposure to SARS
C1260451|T033|PT|V01.82|ICD9CM|Exposure to SARS-associated coronavirus|Exposure to SARS-associated coronavirus
C1455969|T033|PT|V01.83|ICD9CM|Contact with or exposure to escherichia coli (E. coli)|Contact with or exposure to escherichia coli (E. coli)
C1455969|T033|AB|V01.83|ICD9CM|E. coli contact/exp|E. coli contact/exp
C1455970|T033|PT|V01.84|ICD9CM|Contact with or exposure to meningococcus|Contact with or exposure to meningococcus
C1455970|T033|AB|V01.84|ICD9CM|Meningococcus contact|Meningococcus contact
C0260348|T033|AB|V01.89|ICD9CM|Communic dis contact NEC|Communic dis contact NEC
C0260348|T033|PT|V01.89|ICD9CM|Contact with or exposure to other communicable diseases|Contact with or exposure to other communicable diseases
C0260339|T033|AB|V01.9|ICD9CM|Communic dis contact NOS|Communic dis contact NOS
C0260339|T033|PT|V01.9|ICD9CM|Contact with or exposure to unspecified communicable disease|Contact with or exposure to unspecified communicable disease
C0481551|T033|HT|V02|ICD9CM|Carrier or suspected carrier of infectious diseases|Carrier or suspected carrier of infectious diseases
C0260351|T033|PT|V02.0|ICD9CM|Carrier or suspected carrier of cholera|Carrier or suspected carrier of cholera
C0260351|T033|AB|V02.0|ICD9CM|Cholera carrier|Cholera carrier
C0260352|T033|PT|V02.1|ICD9CM|Carrier or suspected carrier of typhoid|Carrier or suspected carrier of typhoid
C0260352|T033|AB|V02.1|ICD9CM|Typhoid carrier|Typhoid carrier
C0481434|T033|AB|V02.2|ICD9CM|Amebiasis carrier|Amebiasis carrier
C0481434|T033|PT|V02.2|ICD9CM|Carrier or suspected carrier of amebiasis|Carrier or suspected carrier of amebiasis
C0260354|T033|PT|V02.3|ICD9CM|Carrier or suspected carrier of other gastrointestinal pathogens|Carrier or suspected carrier of other gastrointestinal pathogens
C0260354|T033|AB|V02.3|ICD9CM|GI pathogen carrier NEC|GI pathogen carrier NEC
C0260355|T033|PT|V02.4|ICD9CM|Carrier or suspected carrier of diphtheria|Carrier or suspected carrier of diphtheria
C0260355|T033|AB|V02.4|ICD9CM|Diphtheria carrier|Diphtheria carrier
C0260356|T033|HT|V02.5|ICD9CM|Carrier or suspected carrier of other specified bacterial diseases|Carrier or suspected carrier of other specified bacterial diseases
C0700297|T033|PT|V02.51|ICD9CM|Carrier or suspected carrier of group B streptococcus|Carrier or suspected carrier of group B streptococcus
C0700297|T033|AB|V02.51|ICD9CM|Group b streptoc carrier|Group b streptoc carrier
C0695257|T033|PT|V02.52|ICD9CM|Carrier or suspected carrier of other streptococcus|Carrier or suspected carrier of other streptococcus
C0695257|T033|AB|V02.52|ICD9CM|Streptococus carrier NEC|Streptococus carrier NEC
C2355591|T033|PT|V02.53|ICD9CM|Carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus|Carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus
C2355591|T033|AB|V02.53|ICD9CM|Meth susc Staph carrier|Meth susc Staph carrier
C2350012|T033|PT|V02.54|ICD9CM|Carrier or suspected carrier of Methicillin resistant Staphylococcus aureus|Carrier or suspected carrier of Methicillin resistant Staphylococcus aureus
C2350012|T033|AB|V02.54|ICD9CM|Meth resis Staph carrier|Meth resis Staph carrier
C0260356|T033|AB|V02.59|ICD9CM|Bacteria dis carrier NEC|Bacteria dis carrier NEC
C0260356|T033|PT|V02.59|ICD9CM|Carrier or suspected carrier of other specified bacterial diseases|Carrier or suspected carrier of other specified bacterial diseases
C0543428|T033|HT|V02.6|ICD9CM|Carrier or suspected carrier of viral hepatitis|Carrier or suspected carrier of viral hepatitis
C0549126|T033|AB|V02.60|ICD9CM|Viral hep carrier NOS|Viral hep carrier NOS
C0549126|T033|PT|V02.60|ICD9CM|Viral hepatitis carrier, unspecified|Viral hepatitis carrier, unspecified
C2911652|T033|AB|V02.61|ICD9CM|Hepatitis B carrier|Hepatitis B carrier
C2911652|T033|PT|V02.61|ICD9CM|Hepatitis B carrier|Hepatitis B carrier
C0840990|T033|AB|V02.62|ICD9CM|Hepatitis C carrier|Hepatitis C carrier
C0840990|T033|PT|V02.62|ICD9CM|Hepatitis C carrier|Hepatitis C carrier
C0490013|T033|PT|V02.69|ICD9CM|Other viral hepatitis carrier|Other viral hepatitis carrier
C0490013|T033|AB|V02.69|ICD9CM|Viral hep carrier NEC|Viral hep carrier NEC
C0481436|T033|PT|V02.7|ICD9CM|Carrier or suspected carrier of gonorrhea|Carrier or suspected carrier of gonorrhea
C0481436|T033|AB|V02.7|ICD9CM|Gonorrhea carrier|Gonorrhea carrier
C0260359|T033|PT|V02.8|ICD9CM|Carrier or suspected carrier of other venereal diseases|Carrier or suspected carrier of other venereal diseases
C0260359|T033|AB|V02.8|ICD9CM|Venereal dis carrier NEC|Venereal dis carrier NEC
C0260360|T033|AB|V02.9|ICD9CM|Carrier NEC|Carrier NEC
C0260360|T033|PT|V02.9|ICD9CM|Carrier or suspected carrier of other specified infectious organism|Carrier or suspected carrier of other specified infectious organism
C0260361|T033|HT|V03|ICD9CM|Need for prophylactic vaccination and inoculation against bacterial diseases|Need for prophylactic vaccination and inoculation against bacterial diseases
C0260362|T033|PT|V03.0|ICD9CM|Need for prophylactic vaccination and inoculation against cholera alone|Need for prophylactic vaccination and inoculation against cholera alone
C0260362|T033|AB|V03.0|ICD9CM|Vaccin for cholera|Vaccin for cholera
C0260363|T033|PT|V03.1|ICD9CM|Need for prophylactic vaccination and inoculation against typhoid-paratyphoid alone [TAB]|Need for prophylactic vaccination and inoculation against typhoid-paratyphoid alone [TAB]
C0260363|T033|AB|V03.1|ICD9CM|Vacc-typhoid-paratyphoid|Vacc-typhoid-paratyphoid
C0260364|T033|PT|V03.2|ICD9CM|Need for prophylactic vaccination and inoculation against tuberculosis [BCG]|Need for prophylactic vaccination and inoculation against tuberculosis [BCG]
C0260364|T033|AB|V03.2|ICD9CM|Vaccin for tuberculosis|Vaccin for tuberculosis
C0496613|T033|PT|V03.3|ICD9CM|Need for prophylactic vaccination and inoculation against plague|Need for prophylactic vaccination and inoculation against plague
C0496613|T033|AB|V03.3|ICD9CM|Vaccin for plague|Vaccin for plague
C0496614|T033|PT|V03.4|ICD9CM|Need for prophylactic vaccination and inoculation against tularemia|Need for prophylactic vaccination and inoculation against tularemia
C0496614|T033|AB|V03.4|ICD9CM|Vaccin for tularemia|Vaccin for tularemia
C0260367|T033|PT|V03.5|ICD9CM|Need for prophylactic vaccination and inoculation against diphtheria alone|Need for prophylactic vaccination and inoculation against diphtheria alone
C0260367|T033|AB|V03.5|ICD9CM|Vaccin for diphtheria|Vaccin for diphtheria
C0260368|T033|PT|V03.6|ICD9CM|Need for prophylactic vaccination and inoculation against pertussis alone|Need for prophylactic vaccination and inoculation against pertussis alone
C0260368|T033|AB|V03.6|ICD9CM|Vaccin for pertussis|Vaccin for pertussis
C0496615|T033|PT|V03.7|ICD9CM|Need for prophylactic vaccination and inoculation against tetanus toxoid alone|Need for prophylactic vaccination and inoculation against tetanus toxoid alone
C0496615|T033|AB|V03.7|ICD9CM|Tetanus toxoid inoculat|Tetanus toxoid inoculat
C0740080|T033|HT|V03.8|ICD9CM|Need for other specified vaccinations against single bacterial diseases|Need for other specified vaccinations against single bacterial diseases
C0375765|T033|AB|V03.81|ICD9CM|Nd vac hmophlus inflnz b|Nd vac hmophlus inflnz b
C0375765|T033|PT|V03.81|ICD9CM|Other specified vaccinations against hemophilus influenza, type B [Hib]|Other specified vaccinations against hemophilus influenza, type B [Hib]
C0375766|T033|AB|V03.82|ICD9CM|Nd vac strptcs pneumni b|Nd vac strptcs pneumni b
C0375766|T033|PT|V03.82|ICD9CM|Other specified vaccinations against streptococcus pneumoniae [pneumococcus]|Other specified vaccinations against streptococcus pneumoniae [pneumococcus]
C0478550|T033|AB|V03.89|ICD9CM|Nd other specf vacnation|Nd other specf vacnation
C0478550|T033|PT|V03.89|ICD9CM|Other specified vaccination|Other specified vaccination
C0260371|T033|PT|V03.9|ICD9CM|Need for prophylactic vaccination and inoculation against unspecified single bacterial disease|Need for prophylactic vaccination and inoculation against unspecified single bacterial disease
C0260371|T033|AB|V03.9|ICD9CM|Vaccin for bact dis NOS|Vaccin for bact dis NOS
C0375767|T033|HT|V04|ICD9CM|Need for prophylactic vaccination and inoculation against certain diseases|Need for prophylactic vaccination and inoculation against certain diseases
C1962940|T033|PT|V04.0|ICD9CM|Need for prophylactic vaccination and inoculation against poliomyelitis|Need for prophylactic vaccination and inoculation against poliomyelitis
C1962940|T033|AB|V04.0|ICD9CM|Vaccin for poliomyelitis|Vaccin for poliomyelitis
C0260374|T033|PT|V04.1|ICD9CM|Need for prophylactic vaccination and inoculation against smallpox|Need for prophylactic vaccination and inoculation against smallpox
C0260374|T033|AB|V04.1|ICD9CM|Vaccin for smallpox|Vaccin for smallpox
C0700173|T033|PT|V04.2|ICD9CM|Need for prophylactic vaccination and inoculation against measles alone|Need for prophylactic vaccination and inoculation against measles alone
C0700173|T033|AB|V04.2|ICD9CM|Vaccin for measles|Vaccin for measles
C0700174|T033|PT|V04.3|ICD9CM|Need for prophylactic vaccination and inoculation against rubella alone|Need for prophylactic vaccination and inoculation against rubella alone
C0700174|T033|AB|V04.3|ICD9CM|Vaccin for rubella|Vaccin for rubella
C0496621|T033|PT|V04.4|ICD9CM|Need for prophylactic vaccination and inoculation against yellow fever|Need for prophylactic vaccination and inoculation against yellow fever
C0496621|T033|AB|V04.4|ICD9CM|Vaccin for yellow fever|Vaccin for yellow fever
C0728859|T033|PT|V04.5|ICD9CM|Need for prophylactic vaccination and inoculation against rabies|Need for prophylactic vaccination and inoculation against rabies
C0728859|T033|AB|V04.5|ICD9CM|Vaccin for rabies|Vaccin for rabies
C0700172|T033|PT|V04.6|ICD9CM|Need for prophylactic vaccination and inoculation against mumps alone|Need for prophylactic vaccination and inoculation against mumps alone
C0700172|T033|AB|V04.6|ICD9CM|Vaccin for mumps|Vaccin for mumps
C0260380|T033|PT|V04.7|ICD9CM|Need for prophylactic vaccination and inoculation against common cold|Need for prophylactic vaccination and inoculation against common cold
C0260380|T033|AB|V04.7|ICD9CM|Vaccin for common cold|Vaccin for common cold
C1260454|T033|HT|V04.8|ICD9CM|Need for prophylactic vaccination and inoculation against other viral diseases|Need for prophylactic vaccination and inoculation against other viral diseases
C1260452|T033|PT|V04.81|ICD9CM|Need for prophylactic vaccination and inoculation against influenza|Need for prophylactic vaccination and inoculation against influenza
C1260452|T033|AB|V04.81|ICD9CM|Vaccin for influenza|Vaccin for influenza
C1260453|T033|PT|V04.82|ICD9CM|Need for prophylactic vaccination and inoculation against respiratory syncytial virus (RSV)|Need for prophylactic vaccination and inoculation against respiratory syncytial virus (RSV)
C1260453|T033|AB|V04.82|ICD9CM|Vaccination for RSV|Vaccination for RSV
C1260454|T033|PT|V04.89|ICD9CM|Need for prophylactic vaccination and inoculation against other viral diseases|Need for prophylactic vaccination and inoculation against other viral diseases
C1260454|T033|AB|V04.89|ICD9CM|Vaccn/inoc viral dis NEC|Vaccn/inoc viral dis NEC
C0375768|T033|HT|V05|ICD9CM|Need for prophylactic vaccination and inoculation against single diseases|Need for prophylactic vaccination and inoculation against single diseases
C1962938|T033|AB|V05.0|ICD9CM|Arbovirus enceph vaccin|Arbovirus enceph vaccin
C1962938|T033|PT|V05.0|ICD9CM|Need for prophylactic vaccination and inoculation against arthropod-borne viral encephalitis|Need for prophylactic vaccination and inoculation against arthropod-borne viral encephalitis
C0260384|T033|PT|V05.1|ICD9CM|Need for prophylactic vaccination and inoculation against other arthropod-borne viral diseases|Need for prophylactic vaccination and inoculation against other arthropod-borne viral diseases
C0260384|T033|AB|V05.1|ICD9CM|Vacc arboviral dis NEC|Vacc arboviral dis NEC
C0476556|T033|PT|V05.2|ICD9CM|Need for prophylactic vaccination and inoculation against leishmaniasis|Need for prophylactic vaccination and inoculation against leishmaniasis
C0476556|T033|AB|V05.2|ICD9CM|Vaccin for leishmaniasis|Vaccin for leishmaniasis
C0476555|T033|PT|V05.3|ICD9CM|Need for prophylactic vaccination and inoculation against viral hepatitis|Need for prophylactic vaccination and inoculation against viral hepatitis
C0476555|T033|AB|V05.3|ICD9CM|Need prphyl vc vrl hepat|Need prphyl vc vrl hepat
C0375770|T033|PT|V05.4|ICD9CM|Need for prophylactic vaccination and inoculation against varicella|Need for prophylactic vaccination and inoculation against varicella
C0375770|T033|AB|V05.4|ICD9CM|Need prphyl vc varicella|Need prphyl vc varicella
C0260386|T033|PT|V05.8|ICD9CM|Need for prophylactic vaccination and inoculation against other specified disease|Need for prophylactic vaccination and inoculation against other specified disease
C0260386|T033|AB|V05.8|ICD9CM|Vaccin for disease NEC|Vaccin for disease NEC
C0260387|T033|PT|V05.9|ICD9CM|Need for prophylactic vaccination and inoculation against unspecified single disease|Need for prophylactic vaccination and inoculation against unspecified single disease
C0260387|T033|AB|V05.9|ICD9CM|Vaccin for singl dis NOS|Vaccin for singl dis NOS
C0260388|T033|HT|V06|ICD9CM|Need for prophylactic vaccination and inoculation against combinations of diseases|Need for prophylactic vaccination and inoculation against combinations of diseases
C0260389|T033|AB|V06.0|ICD9CM|Vaccin for cholera + tab|Vaccin for cholera + tab
C0260390|T033|AB|V06.1|ICD9CM|Vaccination for DTP-DTaP|Vaccination for DTP-DTaP
C0260391|T033|AB|V06.2|ICD9CM|Vaccin for dtp + tab|Vaccin for dtp + tab
C0260392|T033|AB|V06.3|ICD9CM|Vaccin for dtp + polio|Vaccin for dtp + polio
C0496634|T033|PT|V06.4|ICD9CM|Need for prophylactic vaccination and inoculation against measles-mumps-rubella (MMR)|Need for prophylactic vaccination and inoculation against measles-mumps-rubella (MMR)
C0496634|T033|AB|V06.4|ICD9CM|Vac-measle-mumps-rubella|Vac-measle-mumps-rubella
C0375771|T033|PT|V06.5|ICD9CM|Need for prophylactic vaccination and inoculation against tetanus-diphtheria [Td] (DT)|Need for prophylactic vaccination and inoculation against tetanus-diphtheria [Td] (DT)
C0375771|T033|AB|V06.5|ICD9CM|Vaccination for Td-DT|Vaccination for Td-DT
C0375772|T033|AB|V06.6|ICD9CM|Nd vac strp pnumn/inflnz|Nd vac strp pnumn/inflnz
C0260394|T033|PT|V06.8|ICD9CM|Need for prophylactic vaccination and inoculation against other combinations of diseases|Need for prophylactic vaccination and inoculation against other combinations of diseases
C0260394|T033|AB|V06.8|ICD9CM|Vac-dis combinations NEC|Vac-dis combinations NEC
C0260395|T033|PT|V06.9|ICD9CM|Unspecified combined vaccine|Unspecified combined vaccine
C0260395|T033|AB|V06.9|ICD9CM|Vac-dis combinations NOS|Vac-dis combinations NOS
C2921269|T033|HT|V07|ICD9CM|Need for isolation and other prophylactic or treatment measures|Need for isolation and other prophylactic or treatment measures
C0260397|T033|PT|V07.0|ICD9CM|Need for isolation|Need for isolation
C0260397|T033|AB|V07.0|ICD9CM|Prophylactic isolation|Prophylactic isolation
C0260398|T033|AB|V07.1|ICD9CM|Desensitiza to allergens|Desensitiza to allergens
C0260398|T033|PT|V07.1|ICD9CM|Need for desensitization to allergens|Need for desensitization to allergens
C0260399|T033|PT|V07.2|ICD9CM|Need for prophylactic immunotherapy|Need for prophylactic immunotherapy
C0260399|T033|AB|V07.2|ICD9CM|Prophylact immunotherapy|Prophylact immunotherapy
C0260400|T033|HT|V07.3|ICD9CM|Need for other prophylactic chemotherapy|Need for other prophylactic chemotherapy
C0260400|T033|PT|V07.39|ICD9CM|Need for other prophylactic chemotherapy|Need for other prophylactic chemotherapy
C0260400|T033|AB|V07.39|ICD9CM|Other prophylac chemothr|Other prophylac chemothr
C2911677|T033|AB|V07.4|ICD9CM|Hormone replace postmeno|Hormone replace postmeno
C2911677|T033|PT|V07.4|ICD9CM|Hormone replacement therapy (postmenopausal)|Hormone replacement therapy (postmenopausal)
C2921270|T033|HT|V07.5|ICD9CM|Use of agents affecting estrogen receptors and estrogen levels|Use of agents affecting estrogen receptors and estrogen levels
C2921271|T033|PT|V07.51|ICD9CM|Use of selective estrogen receptor modulators (SERMs)|Use of selective estrogen receptor modulators (SERMs)
C2921271|T033|AB|V07.51|ICD9CM|Use of SERMs|Use of SERMs
C2349826|T033|AB|V07.52|ICD9CM|Use aromatase inhibitors|Use aromatase inhibitors
C2349826|T033|PT|V07.52|ICD9CM|Use of aromatase inhibitors|Use of aromatase inhibitors
C2349833|T033|PT|V07.59|ICD9CM|Use of other agents affecting estrogen receptors and estrogen levels|Use of other agents affecting estrogen receptors and estrogen levels
C2349833|T033|AB|V07.59|ICD9CM|Use oth agnt af estrogen|Use oth agnt af estrogen
C2921272|T033|PT|V07.8|ICD9CM|Other specified prophylactic or treatment measure|Other specified prophylactic or treatment measure
C2921272|T033|AB|V07.8|ICD9CM|Prophyl or tx meas NEC|Prophyl or tx meas NEC
C0260402|T033|AB|V07.9|ICD9CM|Prophyl or tx meas NOS|Prophyl or tx meas NOS
C0260402|T033|PT|V07.9|ICD9CM|Unspecified prophylactic or treatment measure|Unspecified prophylactic or treatment measure
C0476550|T033|AB|V08|ICD9CM|Asymp hiv infectn status|Asymp hiv infectn status
C0476550|T033|PT|V08|ICD9CM|Asymptomatic human immunodeficiency virus [HIV] infection status|Asymptomatic human immunodeficiency virus [HIV] infection status
C0375792|T033|HT|V09|ICD9CM|Infection with drug-resistant microorganisms|Infection with drug-resistant microorganisms
C0375777|T033|AB|V09.0|ICD9CM|Inf mcrg rstn pncllins|Inf mcrg rstn pncllins
C0375777|T033|PT|V09.0|ICD9CM|Infection with microorganisms resistant to penicillins|Infection with microorganisms resistant to penicillins
C0375778|T033|AB|V09.1|ICD9CM|Inf mcrg rstn b-lactam|Inf mcrg rstn b-lactam
C0375778|T033|PT|V09.1|ICD9CM|Infection with microorganisms resistant to cephalosporins and other B-lactam antibiotics|Infection with microorganisms resistant to cephalosporins and other B-lactam antibiotics
C0375779|T033|AB|V09.2|ICD9CM|Inf mcrg rstn macrolides|Inf mcrg rstn macrolides
C0375779|T033|PT|V09.2|ICD9CM|Infection with microorganisms resistant to macrolides|Infection with microorganisms resistant to macrolides
C0375780|T033|AB|V09.3|ICD9CM|Inf mcrg rstn ttrcycln|Inf mcrg rstn ttrcycln
C0375780|T033|PT|V09.3|ICD9CM|Infection with microorganisms resistant to tetracyclines|Infection with microorganisms resistant to tetracyclines
C0375781|T033|AB|V09.4|ICD9CM|Inf mcrg rstn amnglcsds|Inf mcrg rstn amnglcsds
C0375781|T033|PT|V09.4|ICD9CM|Infection with microorganisms resistant to aminoglycosides|Infection with microorganisms resistant to aminoglycosides
C0375782|T033|HT|V09.5|ICD9CM|Infection with microorganisms resistant to quinolones and fluoroquinolones|Infection with microorganisms resistant to quinolones and fluoroquinolones
C0375783|T033|AB|V09.50|ICD9CM|Inf mcr rst qn flr nt ml|Inf mcr rst qn flr nt ml
C0375784|T033|AB|V09.51|ICD9CM|Inf mcrg rstn qn flrq ml|Inf mcrg rstn qn flrq ml
C0375784|T033|PT|V09.51|ICD9CM|Infection with microorganisms with resistance to multiple quinolones and fluroquinolones|Infection with microorganisms with resistance to multiple quinolones and fluroquinolones
C0375785|T033|AB|V09.6|ICD9CM|Inf mcrg rstn sulfnmides|Inf mcrg rstn sulfnmides
C0375785|T033|PT|V09.6|ICD9CM|Infection with microorganisms resistant to sulfonamides|Infection with microorganisms resistant to sulfonamides
C0375786|T033|HT|V09.7|ICD9CM|Infection with microorganisms resistant to other specified antimycobacterial agents|Infection with microorganisms resistant to other specified antimycobacterial agents
C0375787|T033|AB|V09.70|ICD9CM|Inf mcr rst oth ag nt ml|Inf mcr rst oth ag nt ml
C0375787|T033|PT|V09.70|ICD9CM|Infection with microorganisms without mention of resistance to multiple antimycobacterial agents|Infection with microorganisms without mention of resistance to multiple antimycobacterial agents
C0375788|T033|AB|V09.71|ICD9CM|Inf mcrg rstn oth ag mlt|Inf mcrg rstn oth ag mlt
C0375788|T033|PT|V09.71|ICD9CM|Infection with microorganisms with resistance to multiple antimycobacterial agents|Infection with microorganisms with resistance to multiple antimycobacterial agents
C0375789|T033|HT|V09.8|ICD9CM|Infection with microorganisms resistant to other specified drugs|Infection with microorganisms resistant to other specified drugs
C0375790|T033|AB|V09.80|ICD9CM|Inf mcr rst ot drg nt ml|Inf mcr rst ot drg nt ml
C0375790|T033|PT|V09.80|ICD9CM|Infection with microorganisms without mention of resistance to multiple drugs|Infection with microorganisms without mention of resistance to multiple drugs
C0375791|T033|AB|V09.81|ICD9CM|Inf mcrg rstn oth drg ml|Inf mcrg rstn oth drg ml
C0375791|T033|PT|V09.81|ICD9CM|Infection with microorganisms with resistance to multiple drugs|Infection with microorganisms with resistance to multiple drugs
C0375792|T033|HT|V09.9|ICD9CM|Infection with drug-resistant microorganisms, unspecified|Infection with drug-resistant microorganisms, unspecified
C0375793|T033|AB|V09.90|ICD9CM|Infc mcrg drgrst nt mult|Infc mcrg drgrst nt mult
C0375794|T033|AB|V09.91|ICD9CM|Infc mcrg drgrst mult|Infc mcrg drgrst mult
C0375794|T033|PT|V09.91|ICD9CM|Infection with drug-resistant microorganisms, unspecified, with multiple drug resistance|Infection with drug-resistant microorganisms, unspecified, with multiple drug resistance
C0260455|T033|HT|V10|ICD9CM|Personal history of malignant neoplasm|Personal history of malignant neoplasm
C0260405|T033|HT|V10.0|ICD9CM|Personal history of malignant neoplasm of gastrointestinal tract|Personal history of malignant neoplasm of gastrointestinal tract
C0260405|T033|AB|V10.00|ICD9CM|Hx of GI malignancy NOS|Hx of GI malignancy NOS
C0260405|T033|PT|V10.00|ICD9CM|Personal history of malignant neoplasm of gastrointestinal tract, unspecified|Personal history of malignant neoplasm of gastrointestinal tract, unspecified
C0260406|T033|AB|V10.01|ICD9CM|Hx of tongue malignancy|Hx of tongue malignancy
C0260406|T033|PT|V10.01|ICD9CM|Personal history of malignant neoplasm of tongue|Personal history of malignant neoplasm of tongue
C0260407|T033|AB|V10.02|ICD9CM|Hx-oral/pharynx malg NEC|Hx-oral/pharynx malg NEC
C0260407|T033|PT|V10.02|ICD9CM|Personal history of malignant neoplasm of other and unspecified oral cavity and pharynx|Personal history of malignant neoplasm of other and unspecified oral cavity and pharynx
C0260408|T033|AB|V10.03|ICD9CM|Hx-esophageal malignancy|Hx-esophageal malignancy
C0260408|T033|PT|V10.03|ICD9CM|Personal history of malignant neoplasm of esophagus|Personal history of malignant neoplasm of esophagus
C0260409|T033|AB|V10.04|ICD9CM|Hx of gastric malignancy|Hx of gastric malignancy
C0260409|T033|PT|V10.04|ICD9CM|Personal history of malignant neoplasm of stomach|Personal history of malignant neoplasm of stomach
C0260410|T033|AB|V10.05|ICD9CM|Hx of colonic malignancy|Hx of colonic malignancy
C0260410|T033|PT|V10.05|ICD9CM|Personal history of malignant neoplasm of large intestine|Personal history of malignant neoplasm of large intestine
C0260411|T033|AB|V10.06|ICD9CM|Hx-rectal & anal malign|Hx-rectal & anal malign
C0260411|T033|PT|V10.06|ICD9CM|Personal history of malignant neoplasm of rectum, rectosigmoid junction, and anus|Personal history of malignant neoplasm of rectum, rectosigmoid junction, and anus
C0260412|T033|AB|V10.07|ICD9CM|Hx of liver malignancy|Hx of liver malignancy
C0260412|T033|PT|V10.07|ICD9CM|Personal history of malignant neoplasm of liver|Personal history of malignant neoplasm of liver
C0260413|T033|AB|V10.09|ICD9CM|Hx of GI malignancy NEC|Hx of GI malignancy NEC
C0260413|T033|PT|V10.09|ICD9CM|Personal history of malignant neoplasm of other gastrointestinal tract|Personal history of malignant neoplasm of other gastrointestinal tract
C0260414|T033|HT|V10.1|ICD9CM|Personal history of malignant neoplasm of trachea, bronchus, and lung|Personal history of malignant neoplasm of trachea, bronchus, and lung
C0260415|T033|AB|V10.11|ICD9CM|Hx-bronchogenic malignan|Hx-bronchogenic malignan
C0260415|T033|PT|V10.11|ICD9CM|Personal history of malignant neoplasm of bronchus and lung|Personal history of malignant neoplasm of bronchus and lung
C0260416|T033|AB|V10.12|ICD9CM|Hx-tracheal malignancy|Hx-tracheal malignancy
C0260416|T033|PT|V10.12|ICD9CM|Personal history of malignant neoplasm of trachea|Personal history of malignant neoplasm of trachea
C0260417|T033|HT|V10.2|ICD9CM|Personal history of malignant neoplasm of other respiratory and intrathoracic organs|Personal history of malignant neoplasm of other respiratory and intrathoracic organs
C0260418|T033|AB|V10.20|ICD9CM|Hx-resp org malignan NOS|Hx-resp org malignan NOS
C0260418|T033|PT|V10.20|ICD9CM|Personal history of malignant neoplasm of respiratory organ, unspecified|Personal history of malignant neoplasm of respiratory organ, unspecified
C0260419|T033|AB|V10.21|ICD9CM|Hx-laryngeal malignancy|Hx-laryngeal malignancy
C0260419|T033|PT|V10.21|ICD9CM|Personal history of malignant neoplasm of larynx|Personal history of malignant neoplasm of larynx
C0260420|T033|AB|V10.22|ICD9CM|Hx-nose/ear/sinus malig|Hx-nose/ear/sinus malig
C0260420|T033|PT|V10.22|ICD9CM|Personal history of malignant neoplasm of nasal cavities, middle ear, and accessory sinuses|Personal history of malignant neoplasm of nasal cavities, middle ear, and accessory sinuses
C0260417|T033|AB|V10.29|ICD9CM|Hx-intrathoracic mal NEC|Hx-intrathoracic mal NEC
C0260417|T033|PT|V10.29|ICD9CM|Personal history of malignant neoplasm of other respiratory and intrathoracic organs|Personal history of malignant neoplasm of other respiratory and intrathoracic organs
C0260421|T033|AB|V10.3|ICD9CM|Hx of breast malignancy|Hx of breast malignancy
C0260421|T033|PT|V10.3|ICD9CM|Personal history of malignant neoplasm of breast|Personal history of malignant neoplasm of breast
C0260422|T033|HT|V10.4|ICD9CM|Personal history of malignant neoplasm of genital organs|Personal history of malignant neoplasm of genital organs
C0260423|T033|AB|V10.40|ICD9CM|Hx-female genit malg NOS|Hx-female genit malg NOS
C0260423|T033|PT|V10.40|ICD9CM|Personal history of malignant neoplasm of female genital organ, unspecified|Personal history of malignant neoplasm of female genital organ, unspecified
C0260424|T033|AB|V10.41|ICD9CM|Hx-cervical malignancy|Hx-cervical malignancy
C0260424|T033|PT|V10.41|ICD9CM|Personal history of malignant neoplasm of cervix uteri|Personal history of malignant neoplasm of cervix uteri
C0260425|T033|AB|V10.42|ICD9CM|Hx-uterus malignancy NEC|Hx-uterus malignancy NEC
C0260425|T033|PT|V10.42|ICD9CM|Personal history of malignant neoplasm of other parts of uterus|Personal history of malignant neoplasm of other parts of uterus
C0260426|T033|AB|V10.43|ICD9CM|Hx of ovarian malignancy|Hx of ovarian malignancy
C0260426|T033|PT|V10.43|ICD9CM|Personal history of malignant neoplasm of ovary|Personal history of malignant neoplasm of ovary
C0260427|T033|AB|V10.44|ICD9CM|Hx-female genit malg NEC|Hx-female genit malg NEC
C0260427|T033|PT|V10.44|ICD9CM|Personal history of malignant neoplasm of other female genital organs|Personal history of malignant neoplasm of other female genital organs
C0260428|T033|AB|V10.45|ICD9CM|Hx-male genit malig NOS|Hx-male genit malig NOS
C0260428|T033|PT|V10.45|ICD9CM|Personal history of malignant neoplasm of male genital organ, unspecified|Personal history of malignant neoplasm of male genital organ, unspecified
C0260429|T033|AB|V10.46|ICD9CM|Hx-prostatic malignancy|Hx-prostatic malignancy
C0260429|T033|PT|V10.46|ICD9CM|Personal history of malignant neoplasm of prostate|Personal history of malignant neoplasm of prostate
C0260430|T033|AB|V10.47|ICD9CM|Hx-testicular malignancy|Hx-testicular malignancy
C0260430|T033|PT|V10.47|ICD9CM|Personal history of malignant neoplasm of testis|Personal history of malignant neoplasm of testis
C0700112|T033|AB|V10.48|ICD9CM|Hx-epididymis malignancy|Hx-epididymis malignancy
C0700112|T033|PT|V10.48|ICD9CM|Personal history of malignant neoplasm of epididymis|Personal history of malignant neoplasm of epididymis
C0260431|T033|AB|V10.49|ICD9CM|Hx-male genit malig NEC|Hx-male genit malig NEC
C0260431|T033|PT|V10.49|ICD9CM|Personal history of malignant neoplasm of other male genital organs|Personal history of malignant neoplasm of other male genital organs
C0260432|T033|HT|V10.5|ICD9CM|Personal history of malignant neoplasm of urinary organs|Personal history of malignant neoplasm of urinary organs
C0260433|T033|AB|V10.50|ICD9CM|Hx-urinary malignan NOS|Hx-urinary malignan NOS
C0260433|T033|PT|V10.50|ICD9CM|Personal history of malignant neoplasm of urinary organ, unspecified|Personal history of malignant neoplasm of urinary organ, unspecified
C0260434|T033|AB|V10.51|ICD9CM|Hx of bladder malignancy|Hx of bladder malignancy
C0260434|T033|PT|V10.51|ICD9CM|Personal history of malignant neoplasm of bladder|Personal history of malignant neoplasm of bladder
C0260435|T033|AB|V10.52|ICD9CM|Hx of kidney malignancy|Hx of kidney malignancy
C0260435|T033|PT|V10.52|ICD9CM|Personal history of malignant neoplasm of kidney|Personal history of malignant neoplasm of kidney
C0949153|T033|AB|V10.53|ICD9CM|Hx malig renal pelvis|Hx malig renal pelvis
C0949153|T033|PT|V10.53|ICD9CM|Personal history of malignant neoplasm of renal pelvis|Personal history of malignant neoplasm of renal pelvis
C2911290|T033|AB|V10.59|ICD9CM|Hx-urinary malignan NEC|Hx-urinary malignan NEC
C2911290|T033|PT|V10.59|ICD9CM|Personal history of malignant neoplasm of other urinary organs|Personal history of malignant neoplasm of other urinary organs
C0260437|T033|HT|V10.6|ICD9CM|Personal history of leukemia|Personal history of leukemia
C0475686|T033|AB|V10.60|ICD9CM|Hx of leukemia NOS|Hx of leukemia NOS
C0475686|T033|PT|V10.60|ICD9CM|Personal history of leukemia, unspecified|Personal history of leukemia, unspecified
C0260439|T033|AB|V10.61|ICD9CM|Hx of lymphoid leukemia|Hx of lymphoid leukemia
C0260439|T033|PT|V10.61|ICD9CM|Personal history of lymphoid leukemia|Personal history of lymphoid leukemia
C0260440|T033|AB|V10.62|ICD9CM|Hx of myeloid leukemia|Hx of myeloid leukemia
C0260440|T033|PT|V10.62|ICD9CM|Personal history of myeloid leukemia|Personal history of myeloid leukemia
C0260441|T033|AB|V10.63|ICD9CM|Hx of monocytic leukemia|Hx of monocytic leukemia
C0260441|T033|PT|V10.63|ICD9CM|Personal history of monocytic leukemia|Personal history of monocytic leukemia
C0260442|T033|AB|V10.69|ICD9CM|Hx of leukemia NEC|Hx of leukemia NEC
C0260442|T033|PT|V10.69|ICD9CM|Personal history of other leukemia|Personal history of other leukemia
C0349403|T033|HT|V10.7|ICD9CM|Personal history of other lymphatic and hematopoietic neoplasms|Personal history of other lymphatic and hematopoietic neoplasms
C0260444|T033|AB|V10.71|ICD9CM|Hx-lymphosarcoma|Hx-lymphosarcoma
C0260444|T033|PT|V10.71|ICD9CM|Personal history of lymphosarcoma and reticulosarcoma|Personal history of lymphosarcoma and reticulosarcoma
C0260445|T033|AB|V10.72|ICD9CM|Hx-hodgkin's disease|Hx-hodgkin's disease
C0260445|T033|PT|V10.72|ICD9CM|Personal history of hodgkin's disease|Personal history of hodgkin's disease
C0349403|T033|AB|V10.79|ICD9CM|Hx-lymphatic malign NEC|Hx-lymphatic malign NEC
C0349403|T033|PT|V10.79|ICD9CM|Personal history of other lymphatic and hematopoietic neoplasms|Personal history of other lymphatic and hematopoietic neoplasms
C0260446|T033|HT|V10.8|ICD9CM|Personal history of malignant neoplasm of other sites|Personal history of malignant neoplasm of other sites
C0260447|T033|AB|V10.81|ICD9CM|Hx of bone malignancy|Hx of bone malignancy
C0260447|T033|PT|V10.81|ICD9CM|Personal history of malignant neoplasm of bone|Personal history of malignant neoplasm of bone
C0260448|T033|AB|V10.82|ICD9CM|Hx-malig skin melanoma|Hx-malig skin melanoma
C0260448|T033|PT|V10.82|ICD9CM|Personal history of malignant melanoma of skin|Personal history of malignant melanoma of skin
C0260449|T033|AB|V10.83|ICD9CM|Hx-skin malignancy NEC|Hx-skin malignancy NEC
C0260449|T033|PT|V10.83|ICD9CM|Personal history of other malignant neoplasm of skin|Personal history of other malignant neoplasm of skin
C0260450|T033|AB|V10.84|ICD9CM|Hx of eye malignancy|Hx of eye malignancy
C0260450|T033|PT|V10.84|ICD9CM|Personal history of malignant neoplasm of eye|Personal history of malignant neoplasm of eye
C0260451|T033|AB|V10.85|ICD9CM|Hx of brain malignancy|Hx of brain malignancy
C0260451|T033|PT|V10.85|ICD9CM|Personal history of malignant neoplasm of brain|Personal history of malignant neoplasm of brain
C0260452|T033|AB|V10.86|ICD9CM|Hx-malign nerve syst NEC|Hx-malign nerve syst NEC
C0260452|T033|PT|V10.86|ICD9CM|Personal history of malignant neoplasm of other parts of nervous system|Personal history of malignant neoplasm of other parts of nervous system
C0260453|T033|AB|V10.87|ICD9CM|Hx of thyroid malignancy|Hx of thyroid malignancy
C0260453|T033|PT|V10.87|ICD9CM|Personal history of malignant neoplasm of thyroid|Personal history of malignant neoplasm of thyroid
C0260454|T033|AB|V10.88|ICD9CM|Hx-endocrine malign NEC|Hx-endocrine malign NEC
C0260454|T033|PT|V10.88|ICD9CM|Personal history of malignant neoplasm of other endocrine glands and related structures|Personal history of malignant neoplasm of other endocrine glands and related structures
C0260446|T033|AB|V10.89|ICD9CM|Hx of malignancy NEC|Hx of malignancy NEC
C0260446|T033|PT|V10.89|ICD9CM|Personal history of malignant neoplasm of other sites|Personal history of malignant neoplasm of other sites
C2712731|T033|HT|V10.9|ICD9CM|Other and unspecified personal history of malignant neoplasm|Other and unspecified personal history of malignant neoplasm
C0260455|T033|AB|V10.90|ICD9CM|Hx malig neoplasm NOS|Hx malig neoplasm NOS
C0260455|T033|PT|V10.90|ICD9CM|Personal history of unspecified malignant neoplasm|Personal history of unspecified malignant neoplasm
C2712771|T033|AB|V10.91|ICD9CM|Hx malig neuroendo tumor|Hx malig neuroendo tumor
C2712771|T033|PT|V10.91|ICD9CM|Personal history of malignant neuroendocrine tumor|Personal history of malignant neuroendocrine tumor
C0260462|T033|HT|V11|ICD9CM|Personal history of mental disorder|Personal history of mental disorder
C0260457|T033|AB|V11.0|ICD9CM|Hx of schizophrenia|Hx of schizophrenia
C0260457|T033|PT|V11.0|ICD9CM|Personal history of schizophrenia|Personal history of schizophrenia
C0260458|T033|AB|V11.1|ICD9CM|Hx of affective disorder|Hx of affective disorder
C0260458|T033|PT|V11.1|ICD9CM|Personal history of affective disorders|Personal history of affective disorders
C0260459|T033|AB|V11.2|ICD9CM|Hx of neurosis|Hx of neurosis
C0260459|T033|PT|V11.2|ICD9CM|Personal history of neurosis|Personal history of neurosis
C0260460|T033|AB|V11.3|ICD9CM|Hx of alcoholism|Hx of alcoholism
C0260460|T033|PT|V11.3|ICD9CM|Personal history of alcoholism|Personal history of alcoholism
C2921273|T033|AB|V11.4|ICD9CM|Hx combat/stress reactn|Hx combat/stress reactn
C2921273|T033|PT|V11.4|ICD9CM|Personal history of combat and operational stress reaction|Personal history of combat and operational stress reaction
C0260461|T033|AB|V11.8|ICD9CM|Hx-mental disorder NEC|Hx-mental disorder NEC
C0260461|T033|PT|V11.8|ICD9CM|Personal history of other mental disorders|Personal history of other mental disorders
C0260462|T033|AB|V11.9|ICD9CM|Hx-mental disorder NOS|Hx-mental disorder NOS
C0260462|T033|PT|V11.9|ICD9CM|Personal history of unspecified mental disorder|Personal history of unspecified mental disorder
C0260463|T033|HT|V12|ICD9CM|Personal history of certain other diseases|Personal history of certain other diseases
C0260464|T033|HT|V12.0|ICD9CM|Personal history of infectious and parasitic diseases|Personal history of infectious and parasitic diseases
C0375795|T033|PT|V12.00|ICD9CM|Personal history of unspecified infectious and parasitic disease|Personal history of unspecified infectious and parasitic disease
C0375795|T033|AB|V12.00|ICD9CM|Prsnl hst unsp nfct prst|Prsnl hst unsp nfct prst
C0375796|T033|PT|V12.01|ICD9CM|Personal history of tuberculosis|Personal history of tuberculosis
C0375796|T033|AB|V12.01|ICD9CM|Prsnl hst tuberculosis|Prsnl hst tuberculosis
C0375797|T033|PT|V12.02|ICD9CM|Personal history of poliomyelitis|Personal history of poliomyelitis
C0375797|T033|AB|V12.02|ICD9CM|Prsnl hst poliomyelitis|Prsnl hst poliomyelitis
C0375798|T033|PT|V12.03|ICD9CM|Personal history of malaria|Personal history of malaria
C0375798|T033|AB|V12.03|ICD9CM|Personal histry malaria|Personal histry malaria
C2350012|T033|AB|V12.04|ICD9CM|Hx Methicln resist Staph|Hx Methicln resist Staph
C2350012|T033|PT|V12.04|ICD9CM|Personal history of Methicillin resistant Staphylococcus aureus|Personal history of Methicillin resistant Staphylococcus aureus
C0375799|T033|PT|V12.09|ICD9CM|Personal history of other infectious and parasitic diseases|Personal history of other infectious and parasitic diseases
C0375799|T033|AB|V12.09|ICD9CM|Prsnl hst oth nfct parst|Prsnl hst oth nfct parst
C0260465|T033|AB|V12.1|ICD9CM|Hx-nutrition deficiency|Hx-nutrition deficiency
C0260465|T033|PT|V12.1|ICD9CM|Personal history of nutritional deficiency|Personal history of nutritional deficiency
C0260466|T033|HT|V12.2|ICD9CM|Personal history of endocrine, metabolic, and immunity disorders|Personal history of endocrine, metabolic, and immunity disorders
C3161145|T033|AB|V12.21|ICD9CM|Hx gestational diabetes|Hx gestational diabetes
C3161145|T033|PT|V12.21|ICD9CM|Personal history of gestational diabetes|Personal history of gestational diabetes
C3161146|T033|AB|V12.29|ICD9CM|Hx-endocr/meta/immun dis|Hx-endocr/meta/immun dis
C3161146|T033|PT|V12.29|ICD9CM|Personal history of other endocrine, metabolic, and immunity disorders|Personal history of other endocrine, metabolic, and immunity disorders
C0260467|T033|AB|V12.3|ICD9CM|Hx-blood diseases|Hx-blood diseases
C0260467|T033|PT|V12.3|ICD9CM|Personal history of diseases of blood and blood-forming organs|Personal history of diseases of blood and blood-forming organs
C0496723|T033|HT|V12.4|ICD9CM|Personal history of disorders of nervous system and sense organs|Personal history of disorders of nervous system and sense organs
C0496723|T033|AB|V12.40|ICD9CM|Hx nerv sys/snse org NOS|Hx nerv sys/snse org NOS
C0496723|T033|PT|V12.40|ICD9CM|Personal history of unspecified disorder of nervous system and sense organs|Personal history of unspecified disorder of nervous system and sense organs
C0490014|T033|AB|V12.41|ICD9CM|Hx benign neoplasm brain|Hx benign neoplasm brain
C0490014|T033|PT|V12.41|ICD9CM|Personal history of benign neoplasm of the brain|Personal history of benign neoplasm of the brain
C2921394|T033|PT|V12.42|ICD9CM|Personal history of infections of the central nervous system|Personal history of infections of the central nervous system
C2921394|T033|AB|V12.42|ICD9CM|Personl hx infection CNS|Personl hx infection CNS
C0490015|T033|AB|V12.49|ICD9CM|Hx nerv sys/snse org NEC|Hx nerv sys/snse org NEC
C0490015|T033|PT|V12.49|ICD9CM|Personal history of other disorders of nervous system and sense organs|Personal history of other disorders of nervous system and sense organs
C0260469|T033|HT|V12.5|ICD9CM|Personal history of diseases of circulatory system|Personal history of diseases of circulatory system
C0740088|T033|AB|V12.50|ICD9CM|Hx-circulatory dis NOS|Hx-circulatory dis NOS
C0740088|T033|PT|V12.50|ICD9CM|Personal history of unspecified circulatory disease|Personal history of unspecified circulatory disease
C0375800|T033|AB|V12.51|ICD9CM|Hx-ven thrombosis/embols|Hx-ven thrombosis/embols
C0375800|T033|PT|V12.51|ICD9CM|Personal history of venous thrombosis and embolism|Personal history of venous thrombosis and embolism
C0375801|T033|AB|V12.52|ICD9CM|Hx-thrombophlebitis|Hx-thrombophlebitis
C0375801|T033|PT|V12.52|ICD9CM|Personal history of thrombophlebitis|Personal history of thrombophlebitis
C1961116|T033|AB|V12.53|ICD9CM|Hx sudden cardiac arrest|Hx sudden cardiac arrest
C1961116|T033|PT|V12.53|ICD9CM|Personal history of sudden cardiac arrest|Personal history of sudden cardiac arrest
C1955570|T033|AB|V12.54|ICD9CM|Hx TIA/stroke w/o resid|Hx TIA/stroke w/o resid
C0585968|T033|AB|V12.55|ICD9CM|Hx pulmonary embolism|Hx pulmonary embolism
C0585968|T033|PT|V12.55|ICD9CM|Personal history of pulmonary embolism|Personal history of pulmonary embolism
C0375802|T033|AB|V12.59|ICD9CM|Hx-circulatory dis NEC|Hx-circulatory dis NEC
C0375802|T033|PT|V12.59|ICD9CM|Personal history of other diseases of circulatory system|Personal history of other diseases of circulatory system
C0260470|T033|HT|V12.6|ICD9CM|Personal history of diseases of respiratory system|Personal history of diseases of respiratory system
C0035204|T047|AB|V12.60|ICD9CM|Hx resp system dis NOS|Hx resp system dis NOS
C0035204|T047|PT|V12.60|ICD9CM|Personal history of unspecified disease of respiratory system|Personal history of unspecified disease of respiratory system
C2911331|T033|PT|V12.61|ICD9CM|Personal history of pneumonia (recurrent)|Personal history of pneumonia (recurrent)
C2911331|T033|AB|V12.61|ICD9CM|Prsnl hx recur pneumonia|Prsnl hx recur pneumonia
C2921392|T033|AB|V12.69|ICD9CM|Hx resp system dis NEC|Hx resp system dis NEC
C2921392|T033|PT|V12.69|ICD9CM|Personal history of other diseases of respiratory system|Personal history of other diseases of respiratory system
C0260471|T033|HT|V12.7|ICD9CM|Personal history of diseases of digestive system|Personal history of diseases of digestive system
C0740089|T033|PT|V12.70|ICD9CM|Personal history of unspecified digestive disease|Personal history of unspecified digestive disease
C0740089|T033|AB|V12.70|ICD9CM|Prsnl hst unspc dgstv ds|Prsnl hst unspc dgstv ds
C0375803|T033|PT|V12.71|ICD9CM|Personal history of peptic ulcer disease|Personal history of peptic ulcer disease
C0375803|T033|AB|V12.71|ICD9CM|Prsnl hst peptic ulcr ds|Prsnl hst peptic ulcr ds
C0375804|T033|PT|V12.72|ICD9CM|Personal history of colonic polyps|Personal history of colonic polyps
C0375804|T033|AB|V12.72|ICD9CM|Prsnl hst colonic polyps|Prsnl hst colonic polyps
C0375805|T033|PT|V12.79|ICD9CM|Personal history of other diseases of digestive system|Personal history of other diseases of digestive system
C0375805|T033|AB|V12.79|ICD9CM|Prsnl hst ot spf dgst ds|Prsnl hst ot spf dgst ds
C0260472|T033|HT|V13|ICD9CM|Personal history of other diseases|Personal history of other diseases
C0700516|T033|HT|V13.0|ICD9CM|Personal history of disorders of urinary system|Personal history of disorders of urinary system
C0260473|T033|PT|V13.00|ICD9CM|Personal history of unspecified urinary disorder|Personal history of unspecified urinary disorder
C0260473|T033|AB|V13.00|ICD9CM|Prsnl hst urnr dsrd unsp|Prsnl hst urnr dsrd unsp
C0375806|T033|PT|V13.01|ICD9CM|Personal history of urinary calculi|Personal history of urinary calculi
C0375806|T033|AB|V13.01|ICD9CM|Prsnl hst urnr dsrd calc|Prsnl hst urnr dsrd calc
C2921372|T033|AB|V13.02|ICD9CM|Personal history UTI|Personal history UTI
C2921372|T033|PT|V13.02|ICD9CM|Personal history, urinary (tract) infection|Personal history, urinary (tract) infection
C2921393|T033|PT|V13.03|ICD9CM|Personal history, nephrotic syndrome|Personal history, nephrotic syndrome
C2921393|T033|AB|V13.03|ICD9CM|Personl hx nephrotic syn|Personl hx nephrotic syn
C0375807|T033|PT|V13.09|ICD9CM|Personal history of other specified urinary system disorders|Personal history of other specified urinary system disorders
C0375807|T033|AB|V13.09|ICD9CM|Prsn hst ot spf urn dsrd|Prsn hst ot spf urn dsrd
C0260474|T033|AB|V13.1|ICD9CM|Hx-trophoblastic disease|Hx-trophoblastic disease
C0260474|T033|PT|V13.1|ICD9CM|Personal history of trophoblastic disease|Personal history of trophoblastic disease
C0260475|T033|HT|V13.2|ICD9CM|Personal history of other genital system and obstetric disorders|Personal history of other genital system and obstetric disorders
C1135273|T033|AB|V13.21|ICD9CM|History-pre-term labor|History-pre-term labor
C1135273|T033|PT|V13.21|ICD9CM|Personal history of pre-term labor|Personal history of pre-term labor
C1955573|T033|AB|V13.22|ICD9CM|Hx of cervical dysplasia|Hx of cervical dysplasia
C1955573|T033|PT|V13.22|ICD9CM|Personal history of cervical dysplasia|Personal history of cervical dysplasia
C2921279|T033|AB|V13.23|ICD9CM|Hx vaginal dysplasia|Hx vaginal dysplasia
C2921279|T033|PT|V13.23|ICD9CM|Personal history of vaginal dysplasia|Personal history of vaginal dysplasia
C2921281|T033|AB|V13.24|ICD9CM|Hx vulvar dysplasia|Hx vulvar dysplasia
C2921281|T033|PT|V13.24|ICD9CM|Personal history of vulvar dysplasia|Personal history of vulvar dysplasia
C0260475|T033|AB|V13.29|ICD9CM|Hx-genital/obs dis NEC|Hx-genital/obs dis NEC
C0260475|T033|PT|V13.29|ICD9CM|Personal history of other genital system and obstetric disorders|Personal history of other genital system and obstetric disorders
C0260476|T033|AB|V13.3|ICD9CM|Hx-skin/subcutan tis dis|Hx-skin/subcutan tis dis
C0260476|T033|PT|V13.3|ICD9CM|Personal history of diseases of skin and subcutaneous tissue|Personal history of diseases of skin and subcutaneous tissue
C0260477|T033|AB|V13.4|ICD9CM|Hx of arthritis|Hx of arthritis
C0260477|T033|PT|V13.4|ICD9CM|Personal history of arthritis|Personal history of arthritis
C0260478|T033|HT|V13.5|ICD9CM|Personal history of other musculoskeletal disorders|Personal history of other musculoskeletal disorders
C0016663|T046|AB|V13.51|ICD9CM|Hx pathological fracture|Hx pathological fracture
C0016663|T046|PT|V13.51|ICD9CM|Personal history of pathologic fracture|Personal history of pathologic fracture
C2921408|T033|AB|V13.52|ICD9CM|Hx stress fracture|Hx stress fracture
C2921408|T033|PT|V13.52|ICD9CM|Personal history of stress fracture|Personal history of stress fracture
C0260478|T033|AB|V13.59|ICD9CM|Hx musculoskletl dis NEC|Hx musculoskletl dis NEC
C0260478|T033|PT|V13.59|ICD9CM|Personal history of other musculoskeletal disorders|Personal history of other musculoskeletal disorders
C2921283|T033|HT|V13.6|ICD9CM|Personal history of congenital (corrected) malformations|Personal history of congenital (corrected) malformations
C2921284|T033|AB|V13.61|ICD9CM|Hx-hypospadias|Hx-hypospadias
C2921284|T033|PT|V13.61|ICD9CM|Personal history of (corrected) hypospadias|Personal history of (corrected) hypospadias
C2921285|T033|AB|V13.62|ICD9CM|Hx-cong malform-gu|Hx-cong malform-gu
C2921285|T033|PT|V13.62|ICD9CM|Personal history of other (corrected) congenital malformations of genitourinary system|Personal history of other (corrected) congenital malformations of genitourinary system
C2921286|T033|AB|V13.63|ICD9CM|Hx-cong malform-nervous|Hx-cong malform-nervous
C2921286|T033|PT|V13.63|ICD9CM|Personal history of (corrected) congenital malformations of nervous system|Personal history of (corrected) congenital malformations of nervous system
C2921288|T033|AB|V13.64|ICD9CM|Hx-cong malform-eye,face|Hx-cong malform-eye,face
C2921288|T033|PT|V13.64|ICD9CM|Personal history of (corrected) congenital malformations of eye, ear, face and neck|Personal history of (corrected) congenital malformations of eye, ear, face and neck
C2921289|T033|AB|V13.65|ICD9CM|Hx-cong malform-heart|Hx-cong malform-heart
C2921289|T033|PT|V13.65|ICD9CM|Personal history of (corrected) congenital malformations of heart and circulatory system|Personal history of (corrected) congenital malformations of heart and circulatory system
C2921290|T033|AB|V13.66|ICD9CM|Hx-cong malform-resp sys|Hx-cong malform-resp sys
C2921290|T033|PT|V13.66|ICD9CM|Personal history of (corrected) congenital malformations of respiratory system|Personal history of (corrected) congenital malformations of respiratory system
C2921291|T033|AB|V13.67|ICD9CM|Hx-cong malform-digest|Hx-cong malform-digest
C2921291|T033|PT|V13.67|ICD9CM|Personal history of (corrected) congenital malformations of digestive system|Personal history of (corrected) congenital malformations of digestive system
C2921292|T033|AB|V13.68|ICD9CM|Hx-cong malform-skin,ms|Hx-cong malform-skin,ms
C0700232|T033|AB|V13.69|ICD9CM|Hx-congenital malfor NEC|Hx-congenital malfor NEC
C0700232|T033|PT|V13.69|ICD9CM|Personal history of other (corrected) congenital malformations|Personal history of other (corrected) congenital malformations
C0260480|T033|AB|V13.7|ICD9CM|Hx-perinatal problems|Hx-perinatal problems
C0260480|T033|PT|V13.7|ICD9CM|Personal history of perinatal problems|Personal history of perinatal problems
C0260481|T033|HT|V13.8|ICD9CM|Personal history of other specified diseases|Personal history of other specified diseases
C3161147|T033|AB|V13.81|ICD9CM|Hx of anaphylaxis|Hx of anaphylaxis
C3161147|T033|PT|V13.81|ICD9CM|Personal history of anaphylaxis|Personal history of anaphylaxis
C0260481|T033|AB|V13.89|ICD9CM|Hx diseases NEC|Hx diseases NEC
C0260481|T033|PT|V13.89|ICD9CM|Personal history of other specified diseases|Personal history of other specified diseases
C0260482|T033|AB|V13.9|ICD9CM|Hx of disease NOS|Hx of disease NOS
C0260482|T033|PT|V13.9|ICD9CM|Personal history of unspecified disease|Personal history of unspecified disease
C0260483|T033|HT|V14|ICD9CM|Personal history of allergy to medicinal agents|Personal history of allergy to medicinal agents
C0260484|T033|AB|V14.0|ICD9CM|Hx-penicillin allergy|Hx-penicillin allergy
C0260484|T033|PT|V14.0|ICD9CM|Personal history of allergy to penicillin|Personal history of allergy to penicillin
C0260485|T033|AB|V14.1|ICD9CM|Hx-antibiot allergy NEC|Hx-antibiot allergy NEC
C0260485|T033|PT|V14.1|ICD9CM|Personal history of allergy to other antibiotic agent|Personal history of allergy to other antibiotic agent
C0260486|T033|AB|V14.2|ICD9CM|Hx-sulfonamides allergy|Hx-sulfonamides allergy
C0260486|T033|PT|V14.2|ICD9CM|Personal history of allergy to sulfonamides|Personal history of allergy to sulfonamides
C0260487|T033|AB|V14.3|ICD9CM|Hx-anti-infect allergy|Hx-anti-infect allergy
C0260487|T033|PT|V14.3|ICD9CM|Personal history of allergy to other anti-infective agent|Personal history of allergy to other anti-infective agent
C0260488|T033|AB|V14.4|ICD9CM|Hx-anesthetic allergy|Hx-anesthetic allergy
C0260488|T033|PT|V14.4|ICD9CM|Personal history of allergy to anesthetic agent|Personal history of allergy to anesthetic agent
C0260489|T033|AB|V14.5|ICD9CM|Hx-narcotic allergy|Hx-narcotic allergy
C0260489|T033|PT|V14.5|ICD9CM|Personal history of allergy to narcotic agent|Personal history of allergy to narcotic agent
C0260490|T033|AB|V14.6|ICD9CM|Hx-analgesic allergy|Hx-analgesic allergy
C0260490|T033|PT|V14.6|ICD9CM|Personal history of allergy to analgesic agent|Personal history of allergy to analgesic agent
C0260491|T033|AB|V14.7|ICD9CM|Hx-vaccine allergy|Hx-vaccine allergy
C0260491|T033|PT|V14.7|ICD9CM|Personal history of allergy to serum or vaccine|Personal history of allergy to serum or vaccine
C0260492|T033|AB|V14.8|ICD9CM|Hx-drug allergy NEC|Hx-drug allergy NEC
C0260492|T033|PT|V14.8|ICD9CM|Personal history of allergy to other specified medicinal agents|Personal history of allergy to other specified medicinal agents
C0260493|T033|AB|V14.9|ICD9CM|Hx-drug allergy NOS|Hx-drug allergy NOS
C0260493|T033|PT|V14.9|ICD9CM|Personal history of allergy to unspecified medicinal agent|Personal history of allergy to unspecified medicinal agent
C0260494|T033|HT|V15|ICD9CM|Other personal history presenting hazards to health|Other personal history presenting hazards to health
C0877841|T033|HT|V15.0|ICD9CM|Personal history of allergy, other than to medicinal agents, presenting hazards to health|Personal history of allergy, other than to medicinal agents, presenting hazards to health
C0917918|T033|PT|V15.01|ICD9CM|Allergy to peanuts|Allergy to peanuts
C0917918|T033|AB|V15.01|ICD9CM|Hx-peanut allergy|Hx-peanut allergy
C0878710|T033|PT|V15.02|ICD9CM|Allergy to milk products|Allergy to milk products
C0878710|T033|AB|V15.02|ICD9CM|Hx-milk prod allergy|Hx-milk prod allergy
C0917919|T033|PT|V15.03|ICD9CM|Allergy to eggs|Allergy to eggs
C0917919|T033|AB|V15.03|ICD9CM|Hx-eggs allergy|Hx-eggs allergy
C0917920|T033|PT|V15.04|ICD9CM|Allergy to seafood|Allergy to seafood
C0917920|T033|AB|V15.04|ICD9CM|Hx-seafood allergy|Hx-seafood allergy
C0878711|T033|PT|V15.05|ICD9CM|Allergy to other foods|Allergy to other foods
C0878711|T033|AB|V15.05|ICD9CM|Hx-other food allergy|Hx-other food allergy
C2712538|T033|PT|V15.06|ICD9CM|Allergy to insects and arachnids|Allergy to insects and arachnids
C2712538|T033|AB|V15.06|ICD9CM|Hx-allergy insct/arachnd|Hx-allergy insct/arachnd
C0917921|T033|PT|V15.07|ICD9CM|Allergy to latex|Allergy to latex
C0917921|T033|AB|V15.07|ICD9CM|Hx-latex allergy|Hx-latex allergy
C0878713|T033|PT|V15.08|ICD9CM|Allergy to radiographic dye|Allergy to radiographic dye
C0878713|T033|AB|V15.08|ICD9CM|Hx-radiogrphc dye allrgy|Hx-radiogrphc dye allrgy
C0878714|T033|AB|V15.09|ICD9CM|Hx-allergy NEC|Hx-allergy NEC
C0878714|T033|PT|V15.09|ICD9CM|Other allergy, other than to medicinal agents|Other allergy, other than to medicinal agents
C0260495|T033|AB|V15.1|ICD9CM|Hx-major cardiovasc surg|Hx-major cardiovasc surg
C0260495|T033|PT|V15.1|ICD9CM|Personal history of surgery to heart and great vessels, presenting hazards to health|Personal history of surgery to heart and great vessels, presenting hazards to health
C0260496|T033|HT|V15.2|ICD9CM|Personal history of surgery to other organs, presenting hazards to health|Personal history of surgery to other organs, presenting hazards to health
C2911571|T033|AB|V15.21|ICD9CM|Hx in utero proc in preg|Hx in utero proc in preg
C2911571|T033|PT|V15.21|ICD9CM|Personal history of undergoing in utero procedure during pregnancy|Personal history of undergoing in utero procedure during pregnancy
C2911572|T033|AB|V15.22|ICD9CM|Hx in utero proc fetus|Hx in utero proc fetus
C2911572|T033|PT|V15.22|ICD9CM|Personal history of undergoing in utero procedure while a fetus|Personal history of undergoing in utero procedure while a fetus
C0260496|T033|AB|V15.29|ICD9CM|Hx surgery to organs NEC|Hx surgery to organs NEC
C0260496|T033|PT|V15.29|ICD9CM|Personal history of surgery to other organs|Personal history of surgery to other organs
C0260497|T033|AB|V15.3|ICD9CM|Hx of irradiation|Hx of irradiation
C0260497|T033|PT|V15.3|ICD9CM|Personal history of irradiation, presenting hazards to health|Personal history of irradiation, presenting hazards to health
C0260498|T033|HT|V15.4|ICD9CM|Personal history of psychological trauma, presenting hazards to health|Personal history of psychological trauma, presenting hazards to health
C0730554|T033|PT|V15.41|ICD9CM|History of physical abuse|History of physical abuse
C0730554|T033|AB|V15.41|ICD9CM|Hx of physical abuse|Hx of physical abuse
C0730556|T033|PT|V15.42|ICD9CM|History of emotional abuse|History of emotional abuse
C0730556|T033|AB|V15.42|ICD9CM|Hx of emotional abuse|Hx of emotional abuse
C0375810|T033|PT|V15.49|ICD9CM|Other psychological trauma|Other psychological trauma
C0375810|T033|AB|V15.49|ICD9CM|Psychological trauma NEC|Psychological trauma NEC
C0260499|T033|HT|V15.5|ICD9CM|Personal history of injury, presenting hazards to health|Personal history of injury, presenting hazards to health
C2349852|T033|AB|V15.51|ICD9CM|Hx traumatic fracture|Hx traumatic fracture
C2349852|T033|PT|V15.51|ICD9CM|Personal history of traumatic fracture|Personal history of traumatic fracture
C2712539|T033|AB|V15.52|ICD9CM|Hx traumatc brain injury|Hx traumatc brain injury
C2712539|T033|PT|V15.52|ICD9CM|Personal history of traumatic brain injury|Personal history of traumatic brain injury
C2921301|T033|AB|V15.53|ICD9CM|Hx retained FB, rem|Hx retained FB, rem
C2921301|T033|PT|V15.53|ICD9CM|Personal history of retained foreign body fully removed|Personal history of retained foreign body fully removed
C2349854|T033|AB|V15.59|ICD9CM|Hx injury NEC|Hx injury NEC
C2349854|T033|PT|V15.59|ICD9CM|Personal history of other injury|Personal history of other injury
C0260500|T033|AB|V15.6|ICD9CM|Hx of poisoning|Hx of poisoning
C0260500|T033|PT|V15.6|ICD9CM|Personal history of poisoning, presenting hazards to health|Personal history of poisoning, presenting hazards to health
C0260501|T033|AB|V15.7|ICD9CM|Hx of contraception|Hx of contraception
C0260501|T033|PT|V15.7|ICD9CM|Personal history of contraception, presenting hazards to health|Personal history of contraception, presenting hazards to health
C0260502|T033|HT|V15.8|ICD9CM|Other specified personal history presenting hazards to health|Other specified personal history presenting hazards to health
C2712540|T033|AB|V15.80|ICD9CM|Hx failed mod sedation|Hx failed mod sedation
C2712540|T033|PT|V15.80|ICD9CM|Personal history of failed moderate sedation|Personal history of failed moderate sedation
C0260503|T033|AB|V15.81|ICD9CM|Hx of past noncompliance|Hx of past noncompliance
C0260503|T033|PT|V15.81|ICD9CM|Personal history of noncompliance with medical treatment, presenting hazards to health|Personal history of noncompliance with medical treatment, presenting hazards to health
C0040335|T033|AB|V15.82|ICD9CM|History of tobacco use|History of tobacco use
C0040335|T033|PT|V15.82|ICD9CM|Personal history of tobacco use|Personal history of tobacco use
C2712541|T033|AB|V15.83|ICD9CM|Hx underimmunizn status|Hx underimmunizn status
C2712541|T033|PT|V15.83|ICD9CM|Personal history of underimmunization status|Personal history of underimmunization status
C2712542|T033|AB|V15.84|ICD9CM|Hx-contct/expos asbestos|Hx-contct/expos asbestos
C2712542|T033|PT|V15.84|ICD9CM|Personal history of contact with and (suspected) exposure to asbestos|Personal history of contact with and (suspected) exposure to asbestos
C2712543|T033|AB|V15.85|ICD9CM|Hx-cont/exps haz bdy fld|Hx-cont/exps haz bdy fld
C2712543|T033|PT|V15.85|ICD9CM|Personal history of contact with and (suspected) exposure to potentially hazardous body fluids|Personal history of contact with and (suspected) exposure to potentially hazardous body fluids
C2911144|T033|AB|V15.86|ICD9CM|Hx-contact/exposure lead|Hx-contact/exposure lead
C2911144|T033|PT|V15.86|ICD9CM|Personal history of contact with and (suspected) exposure to lead|Personal history of contact with and (suspected) exposure to lead
C1260455|T033|PT|V15.87|ICD9CM|History of extracorporeal membrane oxygenation (ECMO)|History of extracorporeal membrane oxygenation (ECMO)
C1260455|T033|AB|V15.87|ICD9CM|Hx of ECMO|Hx of ECMO
C2919132|T033|PT|V15.88|ICD9CM|History of fall|History of fall
C2919132|T033|AB|V15.88|ICD9CM|Personal history of fall|Personal history of fall
C0260502|T033|AB|V15.89|ICD9CM|Hx-health hazards NEC|Hx-health hazards NEC
C0260502|T033|PT|V15.89|ICD9CM|Other specified personal history presenting hazards to health|Other specified personal history presenting hazards to health
C0260504|T033|AB|V15.9|ICD9CM|Hx-health hazard NOS|Hx-health hazard NOS
C0260504|T033|PT|V15.9|ICD9CM|Unspecified personal history presenting hazards to health|Unspecified personal history presenting hazards to health
C1261378|T033|HT|V16|ICD9CM|Family history of malignant neoplasm|Family history of malignant neoplasm
C0260506|T033|PT|V16.0|ICD9CM|Family history of malignant neoplasm of gastrointestinal tract|Family history of malignant neoplasm of gastrointestinal tract
C0260506|T033|AB|V16.0|ICD9CM|Family hx-gi malignancy|Family hx-gi malignancy
C0260507|T033|PT|V16.1|ICD9CM|Family history of malignant neoplasm of trachea, bronchus, and lung|Family history of malignant neoplasm of trachea, bronchus, and lung
C0260507|T033|AB|V16.1|ICD9CM|Fm hx-trach/bronchog mal|Fm hx-trach/bronchog mal
C0260508|T033|AB|V16.2|ICD9CM|Fam hx-intrathoracic mal|Fam hx-intrathoracic mal
C0260508|T033|PT|V16.2|ICD9CM|Family history of malignant neoplasm of other respiratory and intrathoracic organs|Family history of malignant neoplasm of other respiratory and intrathoracic organs
C1261325|T033|PT|V16.3|ICD9CM|Family history of malignant neoplasm of breast|Family history of malignant neoplasm of breast
C1261325|T033|AB|V16.3|ICD9CM|Family hx-breast malig|Family hx-breast malig
C0260510|T033|HT|V16.4|ICD9CM|Family history of malignant neoplasm of genital organs|Family history of malignant neoplasm of genital organs
C0260510|T033|PT|V16.40|ICD9CM|Family history of malignant neoplasm of genital organ, unspecified|Family history of malignant neoplasm of genital organ, unspecified
C0260510|T033|AB|V16.40|ICD9CM|Fm hx genital malig NOS|Fm hx genital malig NOS
C0490017|T033|PT|V16.41|ICD9CM|Family history of malignant neoplasm of ovary|Family history of malignant neoplasm of ovary
C0490017|T033|AB|V16.41|ICD9CM|Fm hx ovary malignancy|Fm hx ovary malignancy
C1532320|T033|PT|V16.42|ICD9CM|Family history of malignant neoplasm of prostate|Family history of malignant neoplasm of prostate
C1532320|T033|AB|V16.42|ICD9CM|Fm hx prostate malig|Fm hx prostate malig
C0490019|T033|PT|V16.43|ICD9CM|Family history of malignant neoplasm of testis|Family history of malignant neoplasm of testis
C0490019|T033|AB|V16.43|ICD9CM|Fm hx testis malig|Fm hx testis malig
C0490020|T033|PT|V16.49|ICD9CM|Family history of malignant neoplasm of other genital organs|Family history of malignant neoplasm of other genital organs
C0490020|T033|AB|V16.49|ICD9CM|Fm hx genital malig NEC|Fm hx genital malig NEC
C0260511|T033|HT|V16.5|ICD9CM|Family history of malignant neoplasm of urinary organs|Family history of malignant neoplasm of urinary organs
C0700102|T033|PT|V16.51|ICD9CM|Family history of malignant neoplasm of kidney|Family history of malignant neoplasm of kidney
C0700102|T033|AB|V16.51|ICD9CM|Family hx-kidney malig|Family hx-kidney malig
C1955574|T033|AB|V16.52|ICD9CM|Fam hx-bladder malig|Fam hx-bladder malig
C1955574|T033|PT|V16.52|ICD9CM|Family history of malignant neoplasm, bladder|Family history of malignant neoplasm, bladder
C2911212|T033|AB|V16.59|ICD9CM|Fam hx-urinry malig NEC|Fam hx-urinry malig NEC
C2911212|T033|PT|V16.59|ICD9CM|Family history of malignant neoplasm of other urinary organs|Family history of malignant neoplasm of other urinary organs
C0260512|T033|PT|V16.6|ICD9CM|Family history of leukemia|Family history of leukemia
C0260512|T033|AB|V16.6|ICD9CM|Family hx-leukemia|Family hx-leukemia
C2586326|T033|AB|V16.7|ICD9CM|Fam hx-lymph neoplas NEC|Fam hx-lymph neoplas NEC
C2586326|T033|PT|V16.7|ICD9CM|Family history of other lymphatic and hematopoietic neoplasms|Family history of other lymphatic and hematopoietic neoplasms
C0260514|T033|PT|V16.8|ICD9CM|Family history of other specified malignant neoplasm|Family history of other specified malignant neoplasm
C0260514|T033|AB|V16.8|ICD9CM|Family hx-malignancy NEC|Family hx-malignancy NEC
C1261378|T033|PT|V16.9|ICD9CM|Family history of unspecified malignant neoplasm|Family history of unspecified malignant neoplasm
C1261378|T033|AB|V16.9|ICD9CM|Family hx-malignancy NOS|Family hx-malignancy NOS
C0260516|T033|HT|V17|ICD9CM|Family history of certain chronic disabling diseases|Family history of certain chronic disabling diseases
C0260517|T033|AB|V17.0|ICD9CM|Fam hx-psychiatric cond|Fam hx-psychiatric cond
C0260517|T033|PT|V17.0|ICD9CM|Family history of psychiatric condition|Family history of psychiatric condition
C0260518|T033|PT|V17.1|ICD9CM|Family history of stroke (cerebrovascular)|Family history of stroke (cerebrovascular)
C0260518|T033|AB|V17.1|ICD9CM|Family hx-stroke|Family hx-stroke
C0260519|T033|AB|V17.2|ICD9CM|Fam hx-neurolog dis NEC|Fam hx-neurolog dis NEC
C0260519|T033|PT|V17.2|ICD9CM|Family history of other neurological diseases|Family history of other neurological diseases
C0260520|T033|AB|V17.3|ICD9CM|Fam hx-ischem heart dis|Fam hx-ischem heart dis
C0260520|T033|PT|V17.3|ICD9CM|Family history of ischemic heart disease|Family history of ischemic heart disease
C1963706|T033|HT|V17.4|ICD9CM|Family history of other cardiovascular diseases|Family history of other cardiovascular diseases
C2825161|T033|AB|V17.41|ICD9CM|Fam hx sudden card death|Fam hx sudden card death
C2825161|T033|PT|V17.41|ICD9CM|Family history of sudden cardiac death (SCD)|Family history of sudden cardiac death (SCD)
C1963707|T033|AB|V17.49|ICD9CM|Fam hx-cardiovas dis NEC|Fam hx-cardiovas dis NEC
C1963707|T033|PT|V17.49|ICD9CM|Family history of other cardiovascular diseases|Family history of other cardiovascular diseases
C0260522|T033|PT|V17.5|ICD9CM|Family history of asthma|Family history of asthma
C0260522|T033|AB|V17.5|ICD9CM|Family hx-asthma|Family hx-asthma
C0260523|T033|AB|V17.6|ICD9CM|Fam hx-chr resp cond NEC|Fam hx-chr resp cond NEC
C0260523|T033|PT|V17.6|ICD9CM|Family history of other chronic respiratory conditions|Family history of other chronic respiratory conditions
C0221565|T033|PT|V17.7|ICD9CM|Family history of arthritis|Family history of arthritis
C0221565|T033|AB|V17.7|ICD9CM|Family hx-arthritis|Family hx-arthritis
C0260524|T033|HT|V17.8|ICD9CM|Family history of other musculoskeletal diseases|Family history of other musculoskeletal diseases
C2911643|T033|PT|V17.81|ICD9CM|Family history of osteoporosis|Family history of osteoporosis
C2911643|T033|AB|V17.81|ICD9CM|Family hx osteoporosis|Family hx osteoporosis
C0260524|T033|AB|V17.89|ICD9CM|Fam hx musculosk dis NEC|Fam hx musculosk dis NEC
C0260524|T033|PT|V17.89|ICD9CM|Family history of other musculoskeletal diseases|Family history of other musculoskeletal diseases
C0260525|T033|HT|V18|ICD9CM|Family history of certain other specific conditions|Family history of certain other specific conditions
C0260526|T033|AB|V18.0|ICD9CM|Fam hx-diabetes mellitus|Fam hx-diabetes mellitus
C0260526|T033|PT|V18.0|ICD9CM|Family history of diabetes mellitus|Family history of diabetes mellitus
C1955577|T033|HT|V18.1|ICD9CM|Family history of other endocrine and metabolic diseases|Family history of other endocrine and metabolic diseases
C1955576|T033|AB|V18.11|ICD9CM|Fam hx MEN syndrome|Fam hx MEN syndrome
C1955576|T033|PT|V18.11|ICD9CM|Family history of multiple endocrine neoplasia [MEN] syndrome|Family history of multiple endocrine neoplasia [MEN] syndrome
C1955577|T033|PT|V18.19|ICD9CM|Family history of other endocrine and metabolic diseases|Family history of other endocrine and metabolic diseases
C1955577|T033|AB|V18.19|ICD9CM|Fm hx endo/metab dis NEC|Fm hx endo/metab dis NEC
C0260528|T033|PT|V18.2|ICD9CM|Family history of anemia|Family history of anemia
C0260528|T033|AB|V18.2|ICD9CM|Family hx-anemia|Family hx-anemia
C0260529|T033|AB|V18.3|ICD9CM|Fam hx-blood disord NEC|Fam hx-blood disord NEC
C0260529|T033|PT|V18.3|ICD9CM|Family history of other blood disorders|Family history of other blood disorders
C0260530|T033|PT|V18.4|ICD9CM|Family history of intellectual disabilities|Family history of intellectual disabilities
C0260530|T033|AB|V18.4|ICD9CM|Fm hx-intellect disablty|Fm hx-intellect disablty
C0496716|T033|HT|V18.5|ICD9CM|Family history of digestive disorders|Family history of digestive disorders
C2911243|T033|PT|V18.51|ICD9CM|Family history of colonic polyps|Family history of colonic polyps
C2911243|T033|AB|V18.51|ICD9CM|Family hx colonic polyps|Family hx colonic polyps
C2911244|T033|AB|V18.59|ICD9CM|Fam hx digest disord NEC|Fam hx digest disord NEC
C2911244|T033|PT|V18.59|ICD9CM|Family history of other digestive disorders|Family history of other digestive disorders
C1261328|T033|HT|V18.6|ICD9CM|Family history of kidney diseases|Family history of kidney diseases
C0455422|T033|AB|V18.61|ICD9CM|Fam hx-polycystic kidney|Fam hx-polycystic kidney
C0455422|T033|PT|V18.61|ICD9CM|Family history of polycystic kidney|Family history of polycystic kidney
C0695259|T033|AB|V18.69|ICD9CM|Fam hx-kidney dis NEC|Fam hx-kidney dis NEC
C0695259|T033|PT|V18.69|ICD9CM|Family history of other kidney diseases|Family history of other kidney diseases
C0260533|T033|PT|V18.7|ICD9CM|Family history of other genitourinary diseases|Family history of other genitourinary diseases
C0260533|T033|AB|V18.7|ICD9CM|Family hx-gu disease NEC|Family hx-gu disease NEC
C0260534|T033|PT|V18.8|ICD9CM|Family history of infectious and parasitic diseases|Family history of infectious and parasitic diseases
C0260534|T033|AB|V18.8|ICD9CM|Fm hx-infect/parasit dis|Fm hx-infect/parasit dis
C0007294|T033|AB|V18.9|ICD9CM|Fam hx genet dis carrier|Fam hx genet dis carrier
C0007294|T033|PT|V18.9|ICD9CM|Family history of genetic disease carrier|Family history of genetic disease carrier
C0260535|T033|HT|V19|ICD9CM|Family history of other conditions|Family history of other conditions
C0496709|T033|PT|V19.0|ICD9CM|Family history of blindness or visual loss|Family history of blindness or visual loss
C0496709|T033|AB|V19.0|ICD9CM|Family hx-blindness|Family hx-blindness
C0260537|T033|HT|V19.1|ICD9CM|Family history of other eye disorders|Family history of other eye disorders
C0455397|T033|AB|V19.11|ICD9CM|Family history glaucoma|Family history glaucoma
C0455397|T033|PT|V19.11|ICD9CM|Family history of glaucoma|Family history of glaucoma
C3161148|T033|PT|V19.19|ICD9CM|Family history of other specified eye disorder|Family history of other specified eye disorder
C3161148|T033|AB|V19.19|ICD9CM|Family hx-eye disord NEC|Family hx-eye disord NEC
C0260538|T033|PT|V19.2|ICD9CM|Family history of deafness or hearing loss|Family history of deafness or hearing loss
C0260538|T033|AB|V19.2|ICD9CM|Family hx-deafness|Family hx-deafness
C0260539|T033|PT|V19.3|ICD9CM|Family history of other ear disorders|Family history of other ear disorders
C0260539|T033|AB|V19.3|ICD9CM|Family hx-ear disord NEC|Family hx-ear disord NEC
C0260540|T033|PT|V19.4|ICD9CM|Family history of skin conditions|Family history of skin conditions
C0260540|T033|AB|V19.4|ICD9CM|Family hx-skin condition|Family hx-skin condition
C0260541|T033|AB|V19.5|ICD9CM|Fam hx-congen anomalies|Fam hx-congen anomalies
C0260541|T033|PT|V19.5|ICD9CM|Family history of congenital anomalies|Family history of congenital anomalies
C0260542|T033|PT|V19.6|ICD9CM|Family history of allergic disorders|Family history of allergic disorders
C0260542|T033|AB|V19.6|ICD9CM|Family hx-allergic dis|Family hx-allergic dis
C0015584|T033|AB|V19.7|ICD9CM|Consanguinity|Consanguinity
C0015584|T033|PT|V19.7|ICD9CM|Family history of consanguinity|Family history of consanguinity
C0260535|T033|PT|V19.8|ICD9CM|Family history of other condition|Family history of other condition
C0260535|T033|AB|V19.8|ICD9CM|Family hx-condition NEC|Family hx-condition NEC
C0260543|T033|HT|V20|ICD9CM|Health supervision of infant or child|Health supervision of infant or child
C0476707|T033|AB|V20.0|ICD9CM|Foundling health care|Foundling health care
C0476707|T033|PT|V20.0|ICD9CM|Health supervision of foundling|Health supervision of foundling
C0029629|T033|AB|V20.1|ICD9CM|Care of healthy chld NEC|Care of healthy chld NEC
C0029629|T033|PT|V20.1|ICD9CM|Other healthy infant or child receiving care|Other healthy infant or child receiving care
C0260545|T033|AB|V20.2|ICD9CM|Routin child health exam|Routin child health exam
C0260545|T033|PT|V20.2|ICD9CM|Routine infant or child health check|Routine infant or child health check
C2712857|T033|HT|V20.3|ICD9CM|Newborn health supervision|Newborn health supervision
C2712545|T033|PT|V20.31|ICD9CM|Health supervision for newborn under 8 days old|Health supervision for newborn under 8 days old
C2712545|T033|AB|V20.31|ICD9CM|Health supvsn nb <8 days|Health supvsn nb <8 days
C2712546|T033|PT|V20.32|ICD9CM|Health supervision for newborn 8 to 28 days old|Health supervision for newborn 8 to 28 days old
C2712546|T033|AB|V20.32|ICD9CM|Health supv nb 8-28 days|Health supv nb 8-28 days
C0260546|T033|HT|V21|ICD9CM|Constitutional states in development|Constitutional states in development
C1399001|T033|PT|V21.0|ICD9CM|Period of rapid growth in childhood|Period of rapid growth in childhood
C1399001|T033|AB|V21.0|ICD9CM|Rapid childhood growth|Rapid childhood growth
C0677548|T033|AB|V21.1|ICD9CM|Puberty|Puberty
C0677548|T033|PT|V21.1|ICD9CM|Puberty|Puberty
C0029575|T033|AB|V21.2|ICD9CM|Adolescence growth NEC|Adolescence growth NEC
C0029575|T033|PT|V21.2|ICD9CM|Other development of adolescence|Other development of adolescence
C0878715|T033|HT|V21.3|ICD9CM|Low birth weight status|Low birth weight status
C0878716|T033|PT|V21.30|ICD9CM|Low birth weight status, unspecified|Low birth weight status, unspecified
C0878716|T033|AB|V21.30|ICD9CM|Low birthwt status NOS|Low birthwt status NOS
C0878717|T033|PT|V21.31|ICD9CM|Low birth weight status, less than 500 grams|Low birth weight status, less than 500 grams
C0878717|T033|AB|V21.31|ICD9CM|Low birthwt status <500g|Low birthwt status <500g
C0878718|T033|PT|V21.32|ICD9CM|Low birth weight status, 500-999 grams|Low birth weight status, 500-999 grams
C0878718|T033|AB|V21.32|ICD9CM|Low birthwt 500-999g|Low birthwt 500-999g
C0878719|T033|PT|V21.33|ICD9CM|Low birth weight status, 1000-1499 grams|Low birth weight status, 1000-1499 grams
C0878719|T033|AB|V21.33|ICD9CM|Low birthwt 1000-1499g|Low birthwt 1000-1499g
C0878720|T033|PT|V21.34|ICD9CM|Low birth weight status, 1500-1999 grams|Low birth weight status, 1500-1999 grams
C0878720|T033|AB|V21.34|ICD9CM|Low birthwt 1500-1999g|Low birthwt 1500-1999g
C0878721|T033|PT|V21.35|ICD9CM|Low birth weight status, 2000-2500 grams|Low birth weight status, 2000-2500 grams
C0878721|T033|AB|V21.35|ICD9CM|Low birthwt 2000-2500g|Low birthwt 2000-2500g
C0260548|T033|AB|V21.8|ICD9CM|Constit state in dev NEC|Constit state in dev NEC
C0260548|T033|PT|V21.8|ICD9CM|Other specified constitutional states in development|Other specified constitutional states in development
C0260549|T033|AB|V21.9|ICD9CM|Constit state in dev NOS|Constit state in dev NOS
C0260549|T033|PT|V21.9|ICD9CM|Unspecified constitutional state in development|Unspecified constitutional state in development
C0700573|T033|HT|V22|ICD9CM|Normal pregnancy|Normal pregnancy
C0260550|T033|AB|V22.0|ICD9CM|Supervis normal 1st preg|Supervis normal 1st preg
C0260550|T033|PT|V22.0|ICD9CM|Supervision of normal first pregnancy|Supervision of normal first pregnancy
C0038843|T033|AB|V22.1|ICD9CM|Supervis oth normal preg|Supervis oth normal preg
C0038843|T033|PT|V22.1|ICD9CM|Supervision of other normal pregnancy|Supervision of other normal pregnancy
C0451636|T033|AB|V22.2|ICD9CM|Preg state, incidental|Preg state, incidental
C0451636|T033|PT|V22.2|ICD9CM|Pregnant state, incidental|Pregnant state, incidental
C0260551|T033|HT|V23|ICD9CM|Supervision of high-risk pregnancy|Supervision of high-risk pregnancy
C0260552|T033|AB|V23.0|ICD9CM|Preg w hx of infertility|Preg w hx of infertility
C0260552|T033|PT|V23.0|ICD9CM|Supervision of high-risk pregnancy with history of infertility|Supervision of high-risk pregnancy with history of infertility
C0260553|T033|AB|V23.1|ICD9CM|Preg w hx-trophoblas dis|Preg w hx-trophoblas dis
C0260553|T033|PT|V23.1|ICD9CM|Supervision of high-risk pregnancy with history of trophoblastic disease|Supervision of high-risk pregnancy with history of trophoblastic disease
C0260554|T033|AB|V23.2|ICD9CM|Preg w hx of abortion|Preg w hx of abortion
C0260554|T033|PT|V23.2|ICD9CM|Supervision of high-risk pregnancy with history of abortion|Supervision of high-risk pregnancy with history of abortion
C0260555|T033|AB|V23.3|ICD9CM|Grand multiparity|Grand multiparity
C0260555|T033|PT|V23.3|ICD9CM|Supervision of high-risk pregnancy with grand multiparity|Supervision of high-risk pregnancy with grand multiparity
C0260556|T033|HT|V23.4|ICD9CM|Supervision of high-risk pregnancy with other poor obstetric history|Supervision of high-risk pregnancy with other poor obstetric history
C1135275|T033|AB|V23.41|ICD9CM|Preg w hx pre-term labor|Preg w hx pre-term labor
C1135275|T033|PT|V23.41|ICD9CM|Pregnancy with history of pre-term labor|Pregnancy with history of pre-term labor
C3161149|T033|AB|V23.42|ICD9CM|Preg w hx ectopic preg|Preg w hx ectopic preg
C3161149|T033|PT|V23.42|ICD9CM|Pregnancy with history of ectopic pregnancy|Pregnancy with history of ectopic pregnancy
C0481651|T033|AB|V23.49|ICD9CM|Preg w poor obs hx NEC|Preg w poor obs hx NEC
C0481651|T033|PT|V23.49|ICD9CM|Pregnancy with other poor obstetric history|Pregnancy with other poor obstetric history
C0260557|T033|AB|V23.5|ICD9CM|Preg w poor reproduct hx|Preg w poor reproduct hx
C0260557|T033|PT|V23.5|ICD9CM|Supervision of high-risk pregnancy with other poor reproductive history|Supervision of high-risk pregnancy with other poor reproductive history
C0695231|T033|AB|V23.7|ICD9CM|Insufficnt prenatal care|Insufficnt prenatal care
C0695231|T033|PT|V23.7|ICD9CM|Supervision of high-risk pregnancy with insufficient prenatal care|Supervision of high-risk pregnancy with insufficient prenatal care
C0260559|T033|HT|V23.8|ICD9CM|Supervision of other high-risk pregnancy|Supervision of other high-risk pregnancy
C0740177|T033|PT|V23.81|ICD9CM|Supervision of high-risk pregnancy with elderly primigravida|Supervision of high-risk pregnancy with elderly primigravida
C0740177|T033|AB|V23.81|ICD9CM|Suprv elderly primigrav|Suprv elderly primigrav
C0695244|T033|PT|V23.82|ICD9CM|Supervision of high-risk pregnancy with elderly multigravida|Supervision of high-risk pregnancy with elderly multigravida
C0695244|T033|AB|V23.82|ICD9CM|Suprv elderly multigrav|Suprv elderly multigrav
C0695260|T033|PT|V23.83|ICD9CM|Supervision of high-risk pregnancy with young primigravida|Supervision of high-risk pregnancy with young primigravida
C0695260|T033|AB|V23.83|ICD9CM|Suprv young primigravida|Suprv young primigravida
C0695261|T033|PT|V23.84|ICD9CM|Supervision of high-risk pregnancy with young multigravida|Supervision of high-risk pregnancy with young multigravida
C0695261|T033|AB|V23.84|ICD9CM|Suprv young multigravida|Suprv young multigravida
C2349859|T033|PT|V23.85|ICD9CM|Pregnancy resulting from assisted reproductive technology|Pregnancy resulting from assisted reproductive technology
C2349859|T033|AB|V23.85|ICD9CM|Pregnt-assist repro tech|Pregnt-assist repro tech
C2349861|T047|AB|V23.86|ICD9CM|Preg-hx in utro prev prg|Preg-hx in utro prev prg
C2349861|T047|PT|V23.86|ICD9CM|Pregnancy with history of in utero procedure during previous pregnancy|Pregnancy with history of in utero procedure during previous pregnancy
C3161150|T033|AB|V23.87|ICD9CM|Preg w incon fetl viabil|Preg w incon fetl viabil
C3161150|T033|PT|V23.87|ICD9CM|Pregnancy with inconclusive fetal viability|Pregnancy with inconclusive fetal viability
C0260559|T033|PT|V23.89|ICD9CM|Supervision of other high-risk pregnancy|Supervision of other high-risk pregnancy
C0260559|T033|AB|V23.89|ICD9CM|Suprv high-risk preg NEC|Suprv high-risk preg NEC
C3714588|T033|PT|V23.9|ICD9CM|Supervision of unspecified high-risk pregnancy|Supervision of unspecified high-risk pregnancy
C3714588|T033|AB|V23.9|ICD9CM|Suprv high-risk preg NOS|Suprv high-risk preg NOS
C0260561|T033|HT|V24|ICD9CM|Postpartum care and examination|Postpartum care and examination
C0496662|T033|AB|V24.0|ICD9CM|Postpart care after del|Postpart care after del
C0496662|T033|PT|V24.0|ICD9CM|Postpartum care and examination immediately after delivery|Postpartum care and examination immediately after delivery
C0260563|T033|AB|V24.1|ICD9CM|Postpart care-lactation|Postpart care-lactation
C0260563|T033|PT|V24.1|ICD9CM|Postpartum care and examination of lactating mother|Postpartum care and examination of lactating mother
C0260564|T033|AB|V24.2|ICD9CM|Rout postpart follow-up|Rout postpart follow-up
C0260564|T033|PT|V24.2|ICD9CM|Routine postpartum follow-up|Routine postpartum follow-up
C0375815|T033|HT|V25|ICD9CM|Encounter for contraceptive management|Encounter for contraceptive management
C0375816|T033|HT|V25.0|ICD9CM|Encounter for general counseling and advice on contraceptive management|Encounter for general counseling and advice on contraceptive management
C0375817|T033|PT|V25.01|ICD9CM|General counseling on prescription of oral contraceptives|General counseling on prescription of oral contraceptives
C0375817|T033|AB|V25.01|ICD9CM|Prescrip-oral contracept|Prescrip-oral contracept
C0375818|T033|PT|V25.02|ICD9CM|General counseling on initiation of other contraceptive measures|General counseling on initiation of other contraceptive measures
C0375818|T033|AB|V25.02|ICD9CM|Initiate contracept NEC|Initiate contracept NEC
C1955578|T033|PT|V25.04|ICD9CM|Counseling and instruction in natural family planning to avoid pregnancy|Counseling and instruction in natural family planning to avoid pregnancy
C1955578|T033|AB|V25.04|ICD9CM|Natrl fam pln-avoid preg|Natrl fam pln-avoid preg
C0029624|T033|AB|V25.09|ICD9CM|Contraceptive mangmt NEC|Contraceptive mangmt NEC
C0029624|T033|PT|V25.09|ICD9CM|Other general counseling and advice on contraceptive management|Other general counseling and advice on contraceptive management
C2921302|T033|HT|V25.1|ICD9CM|Encounter for insertion or removal of intrauterine contraceptive device|Encounter for insertion or removal of intrauterine contraceptive device
C0375820|T033|PT|V25.11|ICD9CM|Encounter for insertion of intrauterine contraceptive device|Encounter for insertion of intrauterine contraceptive device
C0375820|T033|AB|V25.11|ICD9CM|Insertion of iud|Insertion of iud
C2921303|T033|PT|V25.12|ICD9CM|Encounter for removal of intrauterine contraceptive device|Encounter for removal of intrauterine contraceptive device
C2921303|T033|AB|V25.12|ICD9CM|Removal of iud|Removal of iud
C2921304|T033|PT|V25.13|ICD9CM|Encounter for removal and reinsertion of intrauterine contraceptive device|Encounter for removal and reinsertion of intrauterine contraceptive device
C2921304|T033|AB|V25.13|ICD9CM|Remove/insert iud|Remove/insert iud
C0362065|T033|AB|V25.2|ICD9CM|Sterilization|Sterilization
C0362065|T033|PT|V25.2|ICD9CM|Sterilization|Sterilization
C0362068|T033|AB|V25.3|ICD9CM|Menstrual extraction|Menstrual extraction
C0362068|T033|PT|V25.3|ICD9CM|Menstrual extraction|Menstrual extraction
C0375823|T033|HT|V25.4|ICD9CM|Encounter for surveillance of previously prescribed contraceptive methods|Encounter for surveillance of previously prescribed contraceptive methods
C0375824|T033|AB|V25.40|ICD9CM|Contracept surveill NOS|Contracept surveill NOS
C0375824|T033|PT|V25.40|ICD9CM|Contraceptive surveillance, unspecified|Contraceptive surveillance, unspecified
C0375825|T033|AB|V25.41|ICD9CM|Contracept pill surveill|Contracept pill surveill
C0375825|T033|PT|V25.41|ICD9CM|Surveillance of contraceptive pill|Surveillance of contraceptive pill
C0260572|T033|AB|V25.42|ICD9CM|Iud surveillance|Iud surveillance
C0260572|T033|PT|V25.42|ICD9CM|Surveillance of intrauterine contraceptive device|Surveillance of intrauterine contraceptive device
C0375827|T033|AB|V25.43|ICD9CM|Srvl mplnt sbdrm cntrcep|Srvl mplnt sbdrm cntrcep
C0375827|T033|PT|V25.43|ICD9CM|Surveillance of implantable subdermal contraceptive|Surveillance of implantable subdermal contraceptive
C0375828|T033|AB|V25.49|ICD9CM|Contracept surveill NEC|Contracept surveill NEC
C0375828|T033|PT|V25.49|ICD9CM|Surveillance of other contraceptive method|Surveillance of other contraceptive method
C0375829|T033|PT|V25.5|ICD9CM|Insertion of implantable subdermal contraceptive|Insertion of implantable subdermal contraceptive
C0375829|T033|AB|V25.5|ICD9CM|Nsrt mplnt sbdrm cntrcep|Nsrt mplnt sbdrm cntrcep
C0260574|T033|AB|V25.8|ICD9CM|Contraceptive mangmt NEC|Contraceptive mangmt NEC
C0260574|T033|PT|V25.8|ICD9CM|Other specified contraceptive management|Other specified contraceptive management
C0375815|T033|AB|V25.9|ICD9CM|Contraceptive mangmt NOS|Contraceptive mangmt NOS
C0375815|T033|PT|V25.9|ICD9CM|Unspecified contraceptive management|Unspecified contraceptive management
C0260576|T033|HT|V26|ICD9CM|Procreative management|Procreative management
C1961128|T033|AB|V26.0|ICD9CM|Tuboplasty or vasoplasty|Tuboplasty or vasoplasty
C1961128|T033|PT|V26.0|ICD9CM|Tuboplasty or vasoplasty after previous sterilization|Tuboplasty or vasoplasty after previous sterilization
C0699895|T033|AB|V26.1|ICD9CM|Artificial insemination|Artificial insemination
C0699895|T033|PT|V26.1|ICD9CM|Artificial insemination|Artificial insemination
C0877842|T033|HT|V26.2|ICD9CM|Procreation management investigation and testing|Procreation management investigation and testing
C0886496|T033|AB|V26.21|ICD9CM|Fertility testing|Fertility testing
C0886496|T033|PT|V26.21|ICD9CM|Fertility testing|Fertility testing
C0878722|T033|PT|V26.22|ICD9CM|Aftercare following sterilization reversal|Aftercare following sterilization reversal
C0878722|T033|AB|V26.22|ICD9CM|Sterilzation rev aftcare|Sterilzation rev aftcare
C0878723|T033|AB|V26.29|ICD9CM|Investigate & test NEC|Investigate & test NEC
C0878723|T033|PT|V26.29|ICD9CM|Other investigation and testing|Other investigation and testing
C0878754|T033|HT|V26.3|ICD9CM|Genetic counseling and testing on procreative management|Genetic counseling and testing on procreative management
C0599986|T033|AB|V26.33|ICD9CM|Genetic counseling|Genetic counseling
C0599986|T033|PT|V26.33|ICD9CM|Genetic counseling|Genetic counseling
C2921306|T033|PT|V26.35|ICD9CM|Encounter for testing of male partner of female with recurrent pregnancy loss|Encounter for testing of male partner of female with recurrent pregnancy loss
C2921306|T033|AB|V26.35|ICD9CM|Test male/fem preg loss|Test male/fem preg loss
C0496640|T033|HT|V26.4|ICD9CM|General counseling and advice on procreative management|General counseling and advice on procreative management
C1955579|T033|AB|V26.41|ICD9CM|Natrl family plan counsl|Natrl family plan counsl
C1955579|T033|PT|V26.41|ICD9CM|Procreative counseling and advice using natural family planning|Procreative counseling and advice using natural family planning
C2712547|T033|PT|V26.42|ICD9CM|Encounter for fertility preservation counseling|Encounter for fertility preservation counseling
C2712547|T033|AB|V26.42|ICD9CM|Fertlity preserv counsel|Fertlity preserv counsel
C1955580|T033|PT|V26.49|ICD9CM|Other procreative management counseling and advice|Other procreative management counseling and advice
C1955580|T033|AB|V26.49|ICD9CM|Procr mgmt cnsl/adv NEC|Procr mgmt cnsl/adv NEC
C0695263|T033|HT|V26.5|ICD9CM|Sterilization status|Sterilization status
C0695264|T033|AB|V26.51|ICD9CM|Tubal ligation status|Tubal ligation status
C0695264|T033|PT|V26.51|ICD9CM|Tubal ligation status|Tubal ligation status
C0695265|T033|AB|V26.52|ICD9CM|Vasectomy status|Vasectomy status
C0695265|T033|PT|V26.52|ICD9CM|Vasectomy status|Vasectomy status
C0478559|T033|HT|V26.8|ICD9CM|Other specified procreative management|Other specified procreative management
C1955581|T033|AB|V26.81|ICD9CM|Assist repro fertility|Assist repro fertility
C1955581|T033|PT|V26.81|ICD9CM|Encounter for assisted reproductive fertility procedure cycle|Encounter for assisted reproductive fertility procedure cycle
C2712548|T033|PT|V26.82|ICD9CM|Encounter for fertility preservation procedure|Encounter for fertility preservation procedure
C2712548|T033|AB|V26.82|ICD9CM|Fertility preserv proc|Fertility preserv proc
C1955583|T033|PT|V26.89|ICD9CM|Other specified procreative management|Other specified procreative management
C1955583|T033|AB|V26.89|ICD9CM|Procreative managemt NEC|Procreative managemt NEC
C0260576|T033|AB|V26.9|ICD9CM|Procreative mangmt NOS|Procreative mangmt NOS
C0260576|T033|PT|V26.9|ICD9CM|Unspecified procreative management|Unspecified procreative management
C1313895|T033|AB|V27.0|ICD9CM|Deliver-single liveborn|Deliver-single liveborn
C1313895|T033|PT|V27.0|ICD9CM|Outcome of delivery, single liveborn|Outcome of delivery, single liveborn
C1313896|T033|AB|V27.1|ICD9CM|Deliver-single stillborn|Deliver-single stillborn
C1313896|T033|PT|V27.1|ICD9CM|Outcome of delivery, single stillborn|Outcome of delivery, single stillborn
C0481459|T033|AB|V27.2|ICD9CM|Deliver-twins, both live|Deliver-twins, both live
C0481459|T033|PT|V27.2|ICD9CM|Outcome of delivery, twins, both liveborn|Outcome of delivery, twins, both liveborn
C0481466|T033|AB|V27.3|ICD9CM|Del-twins, 1 nb, 1 sb|Del-twins, 1 nb, 1 sb
C0481466|T033|PT|V27.3|ICD9CM|Outcome of delivery, twins, one liveborn and one stillborn|Outcome of delivery, twins, one liveborn and one stillborn
C0419377|T033|AB|V27.4|ICD9CM|Deliver-twins, both sb|Deliver-twins, both sb
C0419377|T033|PT|V27.4|ICD9CM|Outcome of delivery, twins, both stillborn|Outcome of delivery, twins, both stillborn
C0260587|T033|AB|V27.5|ICD9CM|Del-mult birth, all live|Del-mult birth, all live
C0260587|T033|PT|V27.5|ICD9CM|Outcome of delivery, other multiple birth, all liveborn|Outcome of delivery, other multiple birth, all liveborn
C0260588|T033|AB|V27.6|ICD9CM|Del-mult brth, some live|Del-mult brth, some live
C0260588|T033|PT|V27.6|ICD9CM|Outcome of delivery, other multiple birth, some liveborn|Outcome of delivery, other multiple birth, some liveborn
C0481671|T033|AB|V27.7|ICD9CM|Del-mult birth, all sb|Del-mult birth, all sb
C0481671|T033|PT|V27.7|ICD9CM|Outcome of delivery, other multiple birth, all stillborn|Outcome of delivery, other multiple birth, all stillborn
C0260590|T033|AB|V27.9|ICD9CM|Outcome of delivery NOS|Outcome of delivery NOS
C0260590|T033|PT|V27.9|ICD9CM|Outcome of delivery, unspecified outcome of delivery|Outcome of delivery, unspecified outcome of delivery
C1719685|T033|HT|V28|ICD9CM|Encounter for antenatal screening of mother|Encounter for antenatal screening of mother
C1962919|T033|PT|V28.0|ICD9CM|Antenatal screening for chromosomal anomalies by amniocentesis|Antenatal screening for chromosomal anomalies by amniocentesis
C1962919|T033|AB|V28.0|ICD9CM|Screening-chromosom anom|Screening-chromosom anom
C0496648|T033|PT|V28.1|ICD9CM|Antenatal screening for raised alpha-fetoprotein levels in amniotic fluid|Antenatal screening for raised alpha-fetoprotein levels in amniotic fluid
C0496648|T033|AB|V28.1|ICD9CM|Screen-alphafetoprotein|Screen-alphafetoprotein
C0260594|T033|PT|V28.2|ICD9CM|Other antenatal screening based on amniocentesis|Other antenatal screening based on amniocentesis
C0260594|T033|AB|V28.2|ICD9CM|Screen by amniocent NEC|Screen by amniocent NEC
C2349862|T033|PT|V28.3|ICD9CM|Encounter for routine screening for malformation using ultrasonics|Encounter for routine screening for malformation using ultrasonics
C2349862|T033|AB|V28.3|ICD9CM|Scr fetl malfrm-ultrasnd|Scr fetl malfrm-ultrasnd
C0260596|T033|PT|V28.4|ICD9CM|Antenatal screening for fetal growth retardation using ultrasonics|Antenatal screening for fetal growth retardation using ultrasonics
C0260596|T033|AB|V28.4|ICD9CM|Screen-fetal retardation|Screen-fetal retardation
C0490021|T033|AB|V28.6|ICD9CM|Antenatal screen strep b|Antenatal screen strep b
C0490021|T033|PT|V28.6|ICD9CM|Antenatal screening for Streptococcus B|Antenatal screening for Streptococcus B
C0260598|T033|HT|V28.8|ICD9CM|Other specified antenatal screening|Other specified antenatal screening
C2349864|T033|PT|V28.81|ICD9CM|Encounter for fetal anatomic survey|Encounter for fetal anatomic survey
C2349864|T033|AB|V28.81|ICD9CM|Scrn fetal anatmc survey|Scrn fetal anatmc survey
C2349865|T033|PT|V28.82|ICD9CM|Encounter for screening for risk of pre-term labor|Encounter for screening for risk of pre-term labor
C2349865|T033|AB|V28.82|ICD9CM|Scrn risk preterm labor|Scrn risk preterm labor
C0260598|T033|AB|V28.89|ICD9CM|Antenatal screening NEC|Antenatal screening NEC
C0260598|T033|PT|V28.89|ICD9CM|Other specified antenatal screening|Other specified antenatal screening
C0260591|T033|AB|V28.9|ICD9CM|Antenatal screening NOS|Antenatal screening NOS
C0260591|T033|PT|V28.9|ICD9CM|Unspecified antenatal screening|Unspecified antenatal screening
C0375832|T033|HT|V29|ICD9CM|Observation and evaluation of newborns for suspected condition not found|Observation and evaluation of newborns for suspected condition not found
C0375833|T033|AB|V29.0|ICD9CM|NB obsrv suspct infect|NB obsrv suspct infect
C0375833|T033|PT|V29.0|ICD9CM|Observation for suspected infectious condition|Observation for suspected infectious condition
C0375834|T033|AB|V29.1|ICD9CM|NB obsrv suspct neurlgcl|NB obsrv suspct neurlgcl
C0375834|T033|PT|V29.1|ICD9CM|Observation for suspected neurological conditions|Observation for suspected neurological conditions
C0375835|T033|PT|V29.2|ICD9CM|Observation and evaluation of newborn for suspected respiratory condition|Observation and evaluation of newborn for suspected respiratory condition
C0375835|T033|AB|V29.2|ICD9CM|Obsrv NB suspc resp cond|Obsrv NB suspc resp cond
C0695266|T033|AB|V29.3|ICD9CM|NB obs genetc/metabl cnd|NB obs genetc/metabl cnd
C0695266|T033|PT|V29.3|ICD9CM|Observation for suspected genetic or metabolic condition|Observation for suspected genetic or metabolic condition
C0481850|T033|AB|V29.8|ICD9CM|NB obsrv oth suspct cond|NB obsrv oth suspct cond
C0481850|T033|PT|V29.8|ICD9CM|Observation for other specified suspected conditions|Observation for other specified suspected conditions
C0490064|T033|AB|V29.9|ICD9CM|NB obsrv unsp suspct cnd|NB obsrv unsp suspct cnd
C0490064|T033|PT|V29.9|ICD9CM|Observation for unspecified suspected conditions|Observation for unspecified suspected conditions
C1313895|T033|HT|V30|ICD9CM|Single liveborn|Single liveborn
C0260601|T033|HT|V30.0|ICD9CM|Single liveborn, born in hospital|Single liveborn, born in hospital
C0260602|T033|AB|V30.00|ICD9CM|Single lb in-hosp w/o cs|Single lb in-hosp w/o cs
C0260602|T033|PT|V30.00|ICD9CM|Single liveborn, born in hospital, delivered without mention of cesarean section|Single liveborn, born in hospital, delivered without mention of cesarean section
C0260603|T033|AB|V30.01|ICD9CM|Single lb in-hosp w cs|Single lb in-hosp w cs
C0260603|T033|PT|V30.01|ICD9CM|Single liveborn, born in hospital, delivered by cesarean section|Single liveborn, born in hospital, delivered by cesarean section
C0260604|T033|AB|V30.1|ICD9CM|Singl livebrn-before adm|Singl livebrn-before adm
C0260604|T033|PT|V30.1|ICD9CM|Single liveborn, born before admission to hospital|Single liveborn, born before admission to hospital
C0481686|T033|AB|V30.2|ICD9CM|Single liveborn-nonhosp|Single liveborn-nonhosp
C0481686|T033|PT|V30.2|ICD9CM|Single liveborn, born outside hospital and not hospitalized|Single liveborn, born outside hospital and not hospitalized
C0481689|T033|HT|V31|ICD9CM|Twin birth, mate liveborn|Twin birth, mate liveborn
C0260607|T033|HT|V31.0|ICD9CM|Twin, mate liveborn, born in hospital|Twin, mate liveborn, born in hospital
C0260608|T033|PT|V31.00|ICD9CM|Twin birth, mate liveborn, born in hospital, delivered without mention of cesarean section|Twin birth, mate liveborn, born in hospital, delivered without mention of cesarean section
C0260608|T033|AB|V31.00|ICD9CM|Twin-mate lb-hosp w/o cs|Twin-mate lb-hosp w/o cs
C0260609|T033|PT|V31.01|ICD9CM|Twin birth, mate liveborn, born in hospital, delivered by cesarean section|Twin birth, mate liveborn, born in hospital, delivered by cesarean section
C0260609|T033|AB|V31.01|ICD9CM|Twin-mate lb-in hos w cs|Twin-mate lb-in hos w cs
C0260610|T033|PT|V31.1|ICD9CM|Twin birth, mate liveborn, born before admission to hospital|Twin birth, mate liveborn, born before admission to hospital
C0260610|T033|AB|V31.1|ICD9CM|Twin, mate lb-before adm|Twin, mate lb-before adm
C0260611|T033|PT|V31.2|ICD9CM|Twin birth, mate liveborn, born outside hospital and not hospitalized|Twin birth, mate liveborn, born outside hospital and not hospitalized
C0260611|T033|AB|V31.2|ICD9CM|Twin, mate lb-nonhosp|Twin, mate lb-nonhosp
C0260612|T033|HT|V32|ICD9CM|Twin birth, mate stillborn|Twin birth, mate stillborn
C0260613|T033|HT|V32.0|ICD9CM|Twin, mate stillborn, born in hospital|Twin, mate stillborn, born in hospital
C0260614|T033|PT|V32.00|ICD9CM|Twin birth, mate stillborn, born in hospital, delivered without mention of cesarean section|Twin birth, mate stillborn, born in hospital, delivered without mention of cesarean section
C0260614|T033|AB|V32.00|ICD9CM|Twin-mate sb-hosp w/o cs|Twin-mate sb-hosp w/o cs
C0260615|T033|PT|V32.01|ICD9CM|Twin birth, mate stillborn, born in hospital, delivered by cesarean section|Twin birth, mate stillborn, born in hospital, delivered by cesarean section
C0260615|T033|AB|V32.01|ICD9CM|Twin-mate sb-hosp w cs|Twin-mate sb-hosp w cs
C0260616|T033|PT|V32.1|ICD9CM|Twin birth, mate stillborn, born before admission to hospital|Twin birth, mate stillborn, born before admission to hospital
C0260616|T033|AB|V32.1|ICD9CM|Twin, mate sb-before adm|Twin, mate sb-before adm
C0260617|T033|PT|V32.2|ICD9CM|Twin birth, mate stillborn, born outside hospital and not hospitalized|Twin birth, mate stillborn, born outside hospital and not hospitalized
C0260617|T033|AB|V32.2|ICD9CM|Twin, mate sb-nonhosp|Twin, mate sb-nonhosp
C0041423|T033|HT|V33|ICD9CM|Twin birth, unspecified whether mate liveborn or stillborn|Twin birth, unspecified whether mate liveborn or stillborn
C0496656|T033|HT|V33.0|ICD9CM|Twin, unspecified, born in hospital|Twin, unspecified, born in hospital
C0260619|T033|AB|V33.00|ICD9CM|Twin-NOS-in hosp w/o cs|Twin-NOS-in hosp w/o cs
C0260620|T033|AB|V33.01|ICD9CM|Twin-NOS-in hosp w cs|Twin-NOS-in hosp w cs
C0260621|T033|PT|V33.1|ICD9CM|Twin birth, unspecified whether mate liveborn or stillborn, born before admission to hospital|Twin birth, unspecified whether mate liveborn or stillborn, born before admission to hospital
C0260621|T033|AB|V33.1|ICD9CM|Twin NOS-before admissn|Twin NOS-before admissn
C0260622|T033|AB|V33.2|ICD9CM|Twin NOS-nonhosp|Twin NOS-nonhosp
C0260623|T033|HT|V34|ICD9CM|Other multiple birth (three or more), mates all liveborn|Other multiple birth (three or more), mates all liveborn
C0260624|T033|HT|V34.0|ICD9CM|Other multiple, mates all liveborn, born in hospital|Other multiple, mates all liveborn, born in hospital
C0260625|T033|AB|V34.00|ICD9CM|Oth mult lb-hosp w/o cs|Oth mult lb-hosp w/o cs
C0260626|T033|AB|V34.01|ICD9CM|Oth mult lb-in hosp w cs|Oth mult lb-in hosp w cs
C0260627|T033|AB|V34.1|ICD9CM|Oth mult nb-before adm|Oth mult nb-before adm
C0260627|T033|PT|V34.1|ICD9CM|Other multiple birth (three or more), mates all liveborn, born before admission to hospital|Other multiple birth (three or more), mates all liveborn, born before admission to hospital
C0260628|T033|AB|V34.2|ICD9CM|Oth multiple nb-nonhosp|Oth multiple nb-nonhosp
C0260628|T033|PT|V34.2|ICD9CM|Other multiple birth (three or more), mates all liveborn, born outside hospital and not hospitalized|Other multiple birth (three or more), mates all liveborn, born outside hospital and not hospitalized
C0260629|T033|HT|V35|ICD9CM|Other multiple birth (three or more), mates all stillborn|Other multiple birth (three or more), mates all stillborn
C0260630|T033|HT|V35.0|ICD9CM|Other multiple, mates all stillborn, born in hospital|Other multiple, mates all stillborn, born in hospital
C0260631|T033|AB|V35.00|ICD9CM|Oth mult sb-hosp w/o cs|Oth mult sb-hosp w/o cs
C0260632|T033|AB|V35.01|ICD9CM|Oth mult sb-in hosp w cs|Oth mult sb-in hosp w cs
C0260633|T033|AB|V35.1|ICD9CM|Oth mult sb-before adm|Oth mult sb-before adm
C0260633|T033|PT|V35.1|ICD9CM|Other multiple birth (three or more), mates all stillborn, born before admission to hospital|Other multiple birth (three or more), mates all stillborn, born before admission to hospital
C0260634|T033|AB|V35.2|ICD9CM|Oth multiple sb-nonhosp|Oth multiple sb-nonhosp
C0260635|T033|HT|V36|ICD9CM|Other multiple birth (three or more), mates liveborn and stillborn|Other multiple birth (three or more), mates liveborn and stillborn
C0260636|T033|HT|V36.0|ICD9CM|Other multiple, mates liveborn and stillborn, born in hospital|Other multiple, mates liveborn and stillborn, born in hospital
C0260637|T033|AB|V36.00|ICD9CM|Mult lb/sb-in hos w/o cs|Mult lb/sb-in hos w/o cs
C0260638|T033|AB|V36.01|ICD9CM|Mult lb/sb-in hosp w cs|Mult lb/sb-in hosp w cs
C0260639|T033|AB|V36.1|ICD9CM|Mult nb/sb-before adm|Mult nb/sb-before adm
C0260640|T033|AB|V36.2|ICD9CM|Multiple nb/sb-nonhosp|Multiple nb/sb-nonhosp
C0260641|T033|HT|V37|ICD9CM|Other multiple birth (three or more), unspecified whether mates liveborn or stillborn|Other multiple birth (three or more), unspecified whether mates liveborn or stillborn
C0260642|T033|HT|V37.0|ICD9CM|Other multiple, unspecified, born in hospital|Other multiple, unspecified, born in hospital
C0260643|T033|AB|V37.00|ICD9CM|Mult brth NOS-hos w/o cs|Mult brth NOS-hos w/o cs
C0260644|T033|AB|V37.01|ICD9CM|Mult birth NOS-hosp w cs|Mult birth NOS-hosp w cs
C0260645|T033|AB|V37.1|ICD9CM|Mult brth NOS-before adm|Mult brth NOS-before adm
C0260646|T033|AB|V37.2|ICD9CM|Mult birth NOS-nonhosp|Mult birth NOS-nonhosp
C0260647|T033|HT|V39|ICD9CM|Liveborn, unspecified whether single, twin, or multiple|Liveborn, unspecified whether single, twin, or multiple
C0260648|T033|HT|V39.0|ICD9CM|Other liveborn, unspecified, born in hospital|Other liveborn, unspecified, born in hospital
C0260649|T033|AB|V39.00|ICD9CM|Liveborn NOS-hosp w/o cs|Liveborn NOS-hosp w/o cs
C0260650|T033|AB|V39.01|ICD9CM|Liveborn NOS-hosp w cs|Liveborn NOS-hosp w cs
C0260651|T033|AB|V39.1|ICD9CM|Liveborn NOS-before adm|Liveborn NOS-before adm
C0260651|T033|PT|V39.1|ICD9CM|Liveborn, unspecified whether single, twin or multiple, born before admission to hospital|Liveborn, unspecified whether single, twin or multiple, born before admission to hospital
C0260652|T033|AB|V39.2|ICD9CM|Liveborn NOS-nonhosp|Liveborn NOS-nonhosp
C0260652|T033|PT|V39.2|ICD9CM|Liveborn, unspecified whether single, twin or multiple, born outside hospital and not hospitalized|Liveborn, unspecified whether single, twin or multiple, born outside hospital and not hospitalized
C0260658|T033|HT|V40|ICD9CM|Mental and behavioral problems|Mental and behavioral problems
C0260654|T033|PT|V40.0|ICD9CM|Mental and behavioral problems with learning|Mental and behavioral problems with learning
C0260654|T033|AB|V40.0|ICD9CM|Problems with learning|Problems with learning
C0260655|T048|PT|V40.1|ICD9CM|Mental and behavioral problems with communication [including speech]|Mental and behavioral problems with communication [including speech]
C0260655|T048|AB|V40.1|ICD9CM|Prob with communication|Prob with communication
C0260656|T033|AB|V40.2|ICD9CM|Mental problems NEC|Mental problems NEC
C0260656|T033|PT|V40.2|ICD9CM|Other mental problems|Other mental problems
C0260657|T033|HT|V40.3|ICD9CM|Other behavioral problems|Other behavioral problems
C3161151|T033|PT|V40.31|ICD9CM|Wandering in diseases classified elsewhere|Wandering in diseases classified elsewhere
C3161151|T033|AB|V40.31|ICD9CM|Wandering-dis elsewhere|Wandering-dis elsewhere
C3161152|T048|AB|V40.39|ICD9CM|Oth spc behavior problem|Oth spc behavior problem
C3161152|T048|PT|V40.39|ICD9CM|Other specified behavioral problem|Other specified behavioral problem
C0260658|T033|AB|V40.9|ICD9CM|Mental/behavior prob NOS|Mental/behavior prob NOS
C0260658|T033|PT|V40.9|ICD9CM|Unspecified mental or behavioral problem|Unspecified mental or behavioral problem
C0260659|T033|HT|V41|ICD9CM|Problems with special senses and other special functions|Problems with special senses and other special functions
C0728984|T033|AB|V41.0|ICD9CM|Problems with sight|Problems with sight
C0728984|T033|PT|V41.0|ICD9CM|Problems with sight|Problems with sight
C0260661|T033|AB|V41.1|ICD9CM|Eye problems NEC|Eye problems NEC
C0260661|T033|PT|V41.1|ICD9CM|Other eye problems|Other eye problems
C0438989|T033|AB|V41.2|ICD9CM|Problems with hearing|Problems with hearing
C0438989|T033|PT|V41.2|ICD9CM|Problems with hearing|Problems with hearing
C0260663|T033|AB|V41.3|ICD9CM|Ear problems NEC|Ear problems NEC
C0260663|T033|PT|V41.3|ICD9CM|Other ear problems|Other ear problems
C0260664|T033|PT|V41.4|ICD9CM|Problems with voice production|Problems with voice production
C0260664|T033|AB|V41.4|ICD9CM|Voice production problem|Voice production problem
C0260665|T033|PT|V41.5|ICD9CM|Problems with smell and taste|Problems with smell and taste
C0260665|T033|AB|V41.5|ICD9CM|Smell and taste problem|Smell and taste problem
C0481706|T033|AB|V41.6|ICD9CM|Problem w swallowing|Problem w swallowing
C0481706|T033|PT|V41.6|ICD9CM|Problems with swallowing and mastication|Problems with swallowing and mastication
C0260667|T033|PT|V41.7|ICD9CM|Problems with sexual function|Problems with sexual function
C0260667|T033|AB|V41.7|ICD9CM|Sexual function problem|Sexual function problem
C0260668|T033|PT|V41.8|ICD9CM|Other problems with special functions|Other problems with special functions
C0260668|T033|AB|V41.8|ICD9CM|Probl w special func NEC|Probl w special func NEC
C0260669|T033|AB|V41.9|ICD9CM|Probl w special func NOS|Probl w special func NOS
C0260669|T033|PT|V41.9|ICD9CM|Unspecified problem with special functions|Unspecified problem with special functions
C0041866|T033|HT|V42|ICD9CM|Organ or tissue replaced by transplant|Organ or tissue replaced by transplant
C0677491|T033|PT|V42.0|ICD9CM|Kidney replaced by transplant|Kidney replaced by transplant
C0677491|T033|AB|V42.0|ICD9CM|Kidney transplant status|Kidney transplant status
C0018812|T033|PT|V42.1|ICD9CM|Heart replaced by transplant|Heart replaced by transplant
C0018812|T033|AB|V42.1|ICD9CM|Heart transplant status|Heart transplant status
C0677631|T033|PT|V42.2|ICD9CM|Heart valve replaced by transplant|Heart valve replaced by transplant
C0677631|T033|AB|V42.2|ICD9CM|Heart valve transplant|Heart valve transplant
C0392099|T033|PT|V42.3|ICD9CM|Skin replaced by transplant|Skin replaced by transplant
C0392099|T033|AB|V42.3|ICD9CM|Skin transplant status|Skin transplant status
C0040750|T033|PT|V42.4|ICD9CM|Bone replaced by transplant|Bone replaced by transplant
C0040750|T033|AB|V42.4|ICD9CM|Bone transplant status|Bone transplant status
C1384683|T033|PT|V42.5|ICD9CM|Cornea replaced by transplant|Cornea replaced by transplant
C1384683|T033|AB|V42.5|ICD9CM|Cornea transplant status|Cornea transplant status
C0392098|T033|PT|V42.6|ICD9CM|Lung replaced by transplant|Lung replaced by transplant
C0392098|T033|AB|V42.6|ICD9CM|Lung transplant status|Lung transplant status
C0023908|T033|PT|V42.7|ICD9CM|Liver replaced by transplant|Liver replaced by transplant
C0023908|T033|AB|V42.7|ICD9CM|Liver transplant status|Liver transplant status
C0490023|T033|HT|V42.8|ICD9CM|Other specified organ or tissue replaced by transplant|Other specified organ or tissue replaced by transplant
C0740179|T033|PT|V42.81|ICD9CM|Bone marrow replaced by transplant|Bone marrow replaced by transplant
C0740179|T033|AB|V42.81|ICD9CM|Trnspl status-bne marrow|Trnspl status-bne marrow
C0490022|T033|PT|V42.82|ICD9CM|Peripheral stem cells replaced by transplant|Peripheral stem cells replaced by transplant
C0490022|T033|AB|V42.82|ICD9CM|Trspl sts-perip stm cell|Trspl sts-perip stm cell
C0684250|T033|PT|V42.83|ICD9CM|Pancreas replaced by transplant|Pancreas replaced by transplant
C0684250|T033|AB|V42.83|ICD9CM|Trnspl status-pancreas|Trnspl status-pancreas
C0728908|T033|PT|V42.84|ICD9CM|Organ or tissue replaced by transplant, intestines|Organ or tissue replaced by transplant, intestines
C0728908|T033|AB|V42.84|ICD9CM|Trnspl status-intestines|Trnspl status-intestines
C0490023|T033|PT|V42.89|ICD9CM|Other specified organ or tissue replaced by transplant|Other specified organ or tissue replaced by transplant
C0490023|T033|AB|V42.89|ICD9CM|Trnspl status organ NEC|Trnspl status organ NEC
C0041866|T033|AB|V42.9|ICD9CM|Transplant status NOS|Transplant status NOS
C0041866|T033|PT|V42.9|ICD9CM|Unspecified organ or tissue replaced by transplant|Unspecified organ or tissue replaced by transplant
C0260672|T033|HT|V43|ICD9CM|Organ or tissue replaced by other means|Organ or tissue replaced by other means
C0260673|T033|PT|V43.0|ICD9CM|Eye globe replaced by other means|Eye globe replaced by other means
C0260673|T033|AB|V43.0|ICD9CM|Eye replacement NEC|Eye replacement NEC
C0033825|T033|PT|V43.1|ICD9CM|Lens replaced by other means|Lens replaced by other means
C0033825|T033|AB|V43.1|ICD9CM|Lens replacement NEC|Lens replacement NEC
C0260674|T033|HT|V43.2|ICD9CM|Heart replaced by other means|Heart replaced by other means
C1260458|T033|AB|V43.22|ICD9CM|Artficial heart replace|Artficial heart replace
C1260458|T033|PT|V43.22|ICD9CM|Organ or tissue replaced by other means, fully implantable artificial heart|Organ or tissue replaced by other means, fully implantable artificial heart
C0260675|T033|AB|V43.3|ICD9CM|Heart valve replac NEC|Heart valve replac NEC
C0260675|T033|PT|V43.3|ICD9CM|Heart valve replaced by other means|Heart valve replaced by other means
C0260676|T033|AB|V43.4|ICD9CM|Blood vessel replac NEC|Blood vessel replac NEC
C0260676|T033|PT|V43.4|ICD9CM|Blood vessel replaced by other means|Blood vessel replaced by other means
C0481487|T033|PT|V43.5|ICD9CM|Bladder replaced by other means|Bladder replaced by other means
C0481487|T033|AB|V43.5|ICD9CM|Bladder replacement NEC|Bladder replacement NEC
C0260678|T033|HT|V43.6|ICD9CM|Joint replaced by other means|Joint replaced by other means
C0375836|T033|AB|V43.60|ICD9CM|Joint replaced unspcf|Joint replaced unspcf
C0375836|T033|PT|V43.60|ICD9CM|Unspecified joint replacement|Unspecified joint replacement
C2186390|T033|AB|V43.61|ICD9CM|Joint replaced shoulder|Joint replaced shoulder
C2186390|T033|PT|V43.61|ICD9CM|Shoulder joint replacement|Shoulder joint replacement
C0375838|T033|PT|V43.62|ICD9CM|Elbow joint replacement|Elbow joint replacement
C0375838|T033|AB|V43.62|ICD9CM|Joint replaced elbow|Joint replaced elbow
C0375839|T033|AB|V43.63|ICD9CM|Joint replaced wrist|Joint replaced wrist
C0375839|T033|PT|V43.63|ICD9CM|Wrist joint replacement|Wrist joint replacement
C0850128|T033|PT|V43.64|ICD9CM|Hip joint replacement|Hip joint replacement
C0850128|T033|AB|V43.64|ICD9CM|Joint replaced hip|Joint replaced hip
C0375841|T033|AB|V43.65|ICD9CM|Joint replaced knee|Joint replaced knee
C0375841|T033|PT|V43.65|ICD9CM|Knee joint replacement|Knee joint replacement
C0375842|T033|PT|V43.66|ICD9CM|Ankle joint replacement|Ankle joint replacement
C0375842|T033|AB|V43.66|ICD9CM|Joint replaced ankle|Joint replaced ankle
C0375843|T033|AB|V43.69|ICD9CM|Oth spcf joint replaced|Oth spcf joint replaced
C0375843|T033|PT|V43.69|ICD9CM|Other joint replacement|Other joint replacement
C0260679|T033|PT|V43.7|ICD9CM|Limb replaced by other means|Limb replaced by other means
C0260679|T033|AB|V43.7|ICD9CM|Limb replacement NEC|Limb replacement NEC
C0260680|T033|HT|V43.8|ICD9CM|Other organ or tissue replaced by other means|Other organ or tissue replaced by other means
C0375844|T033|AB|V43.81|ICD9CM|Larynx replacement|Larynx replacement
C0375844|T033|PT|V43.81|ICD9CM|Larynx replacement|Larynx replacement
C0375845|T033|AB|V43.82|ICD9CM|Breast replacement|Breast replacement
C0375845|T033|PT|V43.82|ICD9CM|Breast replacement|Breast replacement
C0695273|T033|AB|V43.83|ICD9CM|Artific skin repl status|Artific skin repl status
C0695273|T033|PT|V43.83|ICD9CM|Artificial skin replacement|Artificial skin replacement
C0260680|T033|AB|V43.89|ICD9CM|Organ/tiss replacmnt NEC|Organ/tiss replacmnt NEC
C0260680|T033|PT|V43.89|ICD9CM|Other organ or tissue replaced by other means|Other organ or tissue replaced by other means
C0260691|T033|HT|V44|ICD9CM|Artificial opening status|Artificial opening status
C0260682|T033|AB|V44.0|ICD9CM|Tracheostomy status|Tracheostomy status
C0260682|T033|PT|V44.0|ICD9CM|Tracheostomy status|Tracheostomy status
C0260683|T033|AB|V44.1|ICD9CM|Gastrostomy status|Gastrostomy status
C0260683|T033|PT|V44.1|ICD9CM|Gastrostomy status|Gastrostomy status
C0260684|T033|AB|V44.2|ICD9CM|Ileostomy status|Ileostomy status
C0260684|T033|PT|V44.2|ICD9CM|Ileostomy status|Ileostomy status
C0260685|T033|AB|V44.3|ICD9CM|Colostomy status|Colostomy status
C0260685|T033|PT|V44.3|ICD9CM|Colostomy status|Colostomy status
C0260686|T033|AB|V44.4|ICD9CM|Enterostomy status NEC|Enterostomy status NEC
C0260686|T033|PT|V44.4|ICD9CM|Status of other artificial opening of gastrointestinal tract|Status of other artificial opening of gastrointestinal tract
C0260687|T033|HT|V44.5|ICD9CM|Cystostomy status|Cystostomy status
C0260687|T033|AB|V44.50|ICD9CM|Cystostomy status NOS|Cystostomy status NOS
C0260687|T033|PT|V44.50|ICD9CM|Cystostomy, unspecified|Cystostomy, unspecified
C2911489|T033|AB|V44.51|ICD9CM|Cutaneous-vesicos status|Cutaneous-vesicos status
C2911489|T033|PT|V44.51|ICD9CM|Cutaneous-vesicostomy|Cutaneous-vesicostomy
C2911490|T033|AB|V44.52|ICD9CM|Appendico-vesicos status|Appendico-vesicos status
C2911490|T033|PT|V44.52|ICD9CM|Appendico-vesicostomy|Appendico-vesicostomy
C2911491|T033|AB|V44.59|ICD9CM|Cystostomy status NEC|Cystostomy status NEC
C2911491|T033|PT|V44.59|ICD9CM|Other cystostomy|Other cystostomy
C0260688|T033|PT|V44.6|ICD9CM|Other artificial opening of urinary tract status|Other artificial opening of urinary tract status
C0260688|T033|AB|V44.6|ICD9CM|Urinostomy status NEC|Urinostomy status NEC
C0260689|T033|AB|V44.7|ICD9CM|Artificial vagina status|Artificial vagina status
C0260689|T033|PT|V44.7|ICD9CM|Artificial vagina status|Artificial vagina status
C0260690|T033|AB|V44.8|ICD9CM|Artif open status NEC|Artif open status NEC
C0260690|T033|PT|V44.8|ICD9CM|Other artificial opening status|Other artificial opening status
C0260691|T033|AB|V44.9|ICD9CM|Artif open status NOS|Artif open status NOS
C0260691|T033|PT|V44.9|ICD9CM|Unspecified artificial opening status|Unspecified artificial opening status
C0260698|T033|HT|V45|ICD9CM|Other postprocedural states|Other postprocedural states
C2712998|T033|HT|V45.0|ICD9CM|Cardiac pacemaker in situ|Cardiac pacemaker in situ
C0375846|T033|AB|V45.00|ICD9CM|Status cardc dvce unspcf|Status cardc dvce unspcf
C0375846|T033|PT|V45.00|ICD9CM|Unspecified cardiac device in situ|Unspecified cardiac device in situ
C2240369|T033|PT|V45.01|ICD9CM|Cardiac pacemaker in situ|Cardiac pacemaker in situ
C2240369|T033|AB|V45.01|ICD9CM|Status cardiac pacemaker|Status cardiac pacemaker
C2911500|T033|PT|V45.02|ICD9CM|Automatic implantable cardiac defibrillator in situ|Automatic implantable cardiac defibrillator in situ
C2911500|T033|AB|V45.02|ICD9CM|Status autm crd dfbrltr|Status autm crd dfbrltr
C0375848|T033|PT|V45.09|ICD9CM|Other specified cardiac device in situ|Other specified cardiac device in situ
C0375848|T033|AB|V45.09|ICD9CM|Status oth spcf crdc dvc|Status oth spcf crdc dvc
C0260694|T033|HT|V45.1|ICD9CM|Postsurgical renal dialysis status|Postsurgical renal dialysis status
C0481496|T033|AB|V45.11|ICD9CM|Renal dialysis status|Renal dialysis status
C0481496|T033|PT|V45.11|ICD9CM|Renal dialysis status|Renal dialysis status
C2349872|T033|AB|V45.12|ICD9CM|Noncmplnt w renal dialys|Noncmplnt w renal dialys
C2349872|T033|PT|V45.12|ICD9CM|Noncompliance with renal dialysis|Noncompliance with renal dialysis
C0496750|T033|PT|V45.2|ICD9CM|Presence of cerebrospinal fluid drainage device|Presence of cerebrospinal fluid drainage device
C0496750|T033|AB|V45.2|ICD9CM|Ventricular shunt status|Ventricular shunt status
C1401143|T033|PT|V45.3|ICD9CM|Intestinal bypass or anastomosis status|Intestinal bypass or anastomosis status
C1401143|T033|AB|V45.3|ICD9CM|Intestinal bypass status|Intestinal bypass status
C0391994|T033|AB|V45.4|ICD9CM|Arthrodesis status|Arthrodesis status
C0391994|T033|PT|V45.4|ICD9CM|Arthrodesis status|Arthrodesis status
C0375849|T033|HT|V45.5|ICD9CM|Presence of contraceptive device|Presence of contraceptive device
C0344225|T033|PT|V45.51|ICD9CM|Presence of intrauterine contraceptive device|Presence of intrauterine contraceptive device
C0344225|T033|AB|V45.51|ICD9CM|Prsc ntrutr cntrcptv dvc|Prsc ntrutr cntrcptv dvc
C0375850|T033|PT|V45.52|ICD9CM|Presence of subdermal contraceptive implant|Presence of subdermal contraceptive implant
C0375850|T033|AB|V45.52|ICD9CM|Prsc sbdrml cntrcp mplnt|Prsc sbdrml cntrcp mplnt
C0375851|T033|PT|V45.59|ICD9CM|Presence of other contraceptive device|Presence of other contraceptive device
C0375851|T033|AB|V45.59|ICD9CM|Prsc other cntrcptv dvc|Prsc other cntrcptv dvc
C0490025|T033|HT|V45.6|ICD9CM|States following surgery of eye and adnexa|States following surgery of eye and adnexa
C0490024|T033|AB|V45.61|ICD9CM|Cataract extract status|Cataract extract status
C0490024|T033|PT|V45.61|ICD9CM|Cataract extraction status|Cataract extraction status
C0490025|T033|PT|V45.69|ICD9CM|Other states following surgery of eye and adnexa|Other states following surgery of eye and adnexa
C0490025|T033|AB|V45.69|ICD9CM|Post-proc st eye/adn NEC|Post-proc st eye/adn NEC
C0476700|T033|HT|V45.7|ICD9CM|Acquired absence of organ|Acquired absence of organ
C2349873|T033|AB|V45.71|ICD9CM|Acq absnce breast/nipple|Acq absnce breast/nipple
C2349873|T033|PT|V45.71|ICD9CM|Acquired absence of breast and nipple|Acquired absence of breast and nipple
C0490027|T033|AB|V45.72|ICD9CM|Acquire absnce intestine|Acquire absnce intestine
C0490027|T033|PT|V45.72|ICD9CM|Acquired absence of intestine (large) (small)|Acquired absence of intestine (large) (small)
C0476705|T033|AB|V45.73|ICD9CM|Acquired absence kidney|Acquired absence kidney
C0476705|T033|PT|V45.73|ICD9CM|Acquired absence of kidney|Acquired absence of kidney
C0878725|T033|AB|V45.74|ICD9CM|Acq absence urinary trct|Acq absence urinary trct
C0878725|T033|PT|V45.74|ICD9CM|Acquired absence of organ, other parts of urinary tract|Acquired absence of organ, other parts of urinary tract
C0878726|T033|AB|V45.75|ICD9CM|Acq absence of stomach|Acq absence of stomach
C0878726|T033|PT|V45.75|ICD9CM|Acquired absence of organ, stomach|Acquired absence of organ, stomach
C0878727|T033|AB|V45.76|ICD9CM|Acq absence of lung|Acq absence of lung
C0878727|T033|PT|V45.76|ICD9CM|Acquired absence of organ, lung|Acquired absence of organ, lung
C0476706|T033|AB|V45.77|ICD9CM|Acq absnce genital organ|Acq absnce genital organ
C0476706|T033|PT|V45.77|ICD9CM|Acquired absence of organ, genital organs|Acquired absence of organ, genital organs
C0917922|T033|AB|V45.78|ICD9CM|Acquired absence of eye|Acquired absence of eye
C0917922|T033|PT|V45.78|ICD9CM|Acquired absence of organ, eye|Acquired absence of organ, eye
C0886366|T033|AB|V45.79|ICD9CM|Acq absence of organ NEC|Acq absence of organ NEC
C0886366|T033|PT|V45.79|ICD9CM|Other acquired absence of organ|Other acquired absence of organ
C0260698|T033|HT|V45.8|ICD9CM|Other postprocedural status|Other postprocedural status
C0032811|T033|AB|V45.81|ICD9CM|Aortocoronary bypass|Aortocoronary bypass
C0032811|T033|PT|V45.81|ICD9CM|Aortocoronary bypass status|Aortocoronary bypass status
C0375852|T033|PT|V45.82|ICD9CM|Percutaneous transluminal coronary angioplasty status|Percutaneous transluminal coronary angioplasty status
C0375852|T033|AB|V45.82|ICD9CM|Status-post ptca|Status-post ptca
C0375853|T033|AB|V45.83|ICD9CM|Breast impl remov status|Breast impl remov status
C0375853|T033|PT|V45.83|ICD9CM|Breast implant removal status|Breast implant removal status
C2911565|T033|PT|V45.84|ICD9CM|Dental restoration status|Dental restoration status
C2911565|T033|AB|V45.84|ICD9CM|Dental restoratn status|Dental restoratn status
C1260459|T033|AB|V45.85|ICD9CM|Insulin pump status|Insulin pump status
C1260459|T033|PT|V45.85|ICD9CM|Insulin pump status|Insulin pump status
C1719686|T033|PT|V45.86|ICD9CM|Bariatric surgery status|Bariatric surgery status
C1719686|T033|AB|V45.86|ICD9CM|Bariatric surgery status|Bariatric surgery status
C2349874|T033|PT|V45.87|ICD9CM|Transplanted organ removal status|Transplanted organ removal status
C2349874|T033|AB|V45.87|ICD9CM|Trnsplnt orgn rem status|Trnsplnt orgn rem status
C2349876|T033|AB|V45.88|ICD9CM|TPA adm status 24 hr pta|TPA adm status 24 hr pta
C0260698|T033|PT|V45.89|ICD9CM|Other postprocedural status|Other postprocedural status
C0260698|T033|AB|V45.89|ICD9CM|Post-proc states NEC|Post-proc states NEC
C2349878|T033|HT|V46|ICD9CM|Other dependence on machines and devices|Other dependence on machines and devices
C0260700|T033|AB|V46.0|ICD9CM|Dependence on aspirator|Dependence on aspirator
C0260700|T033|PT|V46.0|ICD9CM|Dependence on aspirator|Dependence on aspirator
C1321831|T033|HT|V46.1|ICD9CM|Dependence on respirator [Ventilator]|Dependence on respirator [Ventilator]
C1455974|T033|PT|V46.11|ICD9CM|Dependence on respirator, status|Dependence on respirator, status
C1455974|T033|AB|V46.11|ICD9CM|Respirator depend status|Respirator depend status
C1455975|T033|PT|V46.12|ICD9CM|Encounter for respirator dependence during power failure|Encounter for respirator dependence during power failure
C1455975|T033|AB|V46.12|ICD9CM|Resp depend-powr failure|Resp depend-powr failure
C1561673|T033|PT|V46.13|ICD9CM|Encounter for weaning from respirator [ventilator]|Encounter for weaning from respirator [ventilator]
C1561673|T033|AB|V46.13|ICD9CM|Weaning from respirator|Weaning from respirator
C1561674|T033|AB|V46.14|ICD9CM|Mech comp respirator|Mech comp respirator
C1561674|T033|PT|V46.14|ICD9CM|Mechanical complication of respirator [ventilator]|Mechanical complication of respirator [ventilator]
C2363337|T033|AB|V46.2|ICD9CM|Depend-supplement oxygen|Depend-supplement oxygen
C2363337|T033|PT|V46.2|ICD9CM|Other dependence on machines, supplemental oxygen|Other dependence on machines, supplemental oxygen
C0476582|T033|AB|V46.3|ICD9CM|Wheelchair dependence|Wheelchair dependence
C0476582|T033|PT|V46.3|ICD9CM|Wheelchair dependence|Wheelchair dependence
C0260702|T033|PT|V46.8|ICD9CM|Dependence on other enabling machines|Dependence on other enabling machines
C0260702|T033|AB|V46.8|ICD9CM|Machine dependence NEC|Machine dependence NEC
C0260703|T033|AB|V46.9|ICD9CM|Machine dependence NOS|Machine dependence NOS
C0260703|T033|PT|V46.9|ICD9CM|Unspecified machine dependence|Unspecified machine dependence
C0260704|T033|HT|V47|ICD9CM|Other problems with internal organs|Other problems with internal organs
C0260705|T033|PT|V47.0|ICD9CM|Deficiencies of internal organs|Deficiencies of internal organs
C0260705|T033|AB|V47.0|ICD9CM|Intern organ deficiency|Intern organ deficiency
C0260706|T033|AB|V47.1|ICD9CM|Mech prob w internal org|Mech prob w internal org
C0260706|T033|PT|V47.1|ICD9CM|Mechanical and motor problems with internal organs|Mechanical and motor problems with internal organs
C0260707|T033|AB|V47.2|ICD9CM|Cardiorespirat probl NEC|Cardiorespirat probl NEC
C0260707|T033|PT|V47.2|ICD9CM|Other cardiorespiratory problems|Other cardiorespiratory problems
C0260708|T033|AB|V47.3|ICD9CM|Digestive problems NEC|Digestive problems NEC
C0260708|T033|PT|V47.3|ICD9CM|Other digestive problems|Other digestive problems
C0260709|T033|PT|V47.4|ICD9CM|Other urinary problems|Other urinary problems
C0260709|T033|AB|V47.4|ICD9CM|Urinary problems NEC|Urinary problems NEC
C0260710|T033|AB|V47.5|ICD9CM|Genital problems NEC|Genital problems NEC
C0260710|T033|PT|V47.5|ICD9CM|Other genital problems|Other genital problems
C0260711|T033|AB|V47.9|ICD9CM|Probl w internal org NOS|Probl w internal org NOS
C0260711|T033|PT|V47.9|ICD9CM|Unspecified problems with internal organs|Unspecified problems with internal organs
C0260712|T033|HT|V48|ICD9CM|Problems with head, neck, and trunk|Problems with head, neck, and trunk
C0260713|T033|AB|V48.0|ICD9CM|Deficiencies of head|Deficiencies of head
C0260713|T033|PT|V48.0|ICD9CM|Deficiencies of head|Deficiencies of head
C0260714|T033|AB|V48.1|ICD9CM|Deficiencies neck/trunk|Deficiencies neck/trunk
C0260714|T033|PT|V48.1|ICD9CM|Deficiencies of neck and trunk|Deficiencies of neck and trunk
C0260715|T033|PT|V48.2|ICD9CM|Mechanical and motor problems with head|Mechanical and motor problems with head
C0260715|T033|AB|V48.2|ICD9CM|Mechanical prob w head|Mechanical prob w head
C0260716|T033|AB|V48.3|ICD9CM|Mech prob w neck & trunk|Mech prob w neck & trunk
C0260716|T033|PT|V48.3|ICD9CM|Mechanical and motor problems with neck and trunk|Mechanical and motor problems with neck and trunk
C0260717|T033|AB|V48.4|ICD9CM|Sensory problem w head|Sensory problem w head
C0260717|T033|PT|V48.4|ICD9CM|Sensory problem with head|Sensory problem with head
C0260718|T033|AB|V48.5|ICD9CM|Sensor prob w neck/trunk|Sensor prob w neck/trunk
C0260718|T033|PT|V48.5|ICD9CM|Sensory problem with neck and trunk|Sensory problem with neck and trunk
C0260719|T033|AB|V48.6|ICD9CM|Disfigurements of head|Disfigurements of head
C0260719|T033|PT|V48.6|ICD9CM|Disfigurements of head|Disfigurements of head
C0260720|T033|AB|V48.7|ICD9CM|Disfigurement neck/trunk|Disfigurement neck/trunk
C0260720|T033|PT|V48.7|ICD9CM|Disfigurements of neck and trunk|Disfigurements of neck and trunk
C0260721|T033|PT|V48.8|ICD9CM|Other problems with head, neck, and trunk|Other problems with head, neck, and trunk
C0260721|T033|AB|V48.8|ICD9CM|Prob-head/neck/trunk NEC|Prob-head/neck/trunk NEC
C0260722|T033|AB|V48.9|ICD9CM|Prob-head/neck/trunk NOS|Prob-head/neck/trunk NOS
C0260722|T033|PT|V48.9|ICD9CM|Unspecified problem with head, neck, or trunk|Unspecified problem with head, neck, or trunk
C0878755|T033|HT|V49|ICD9CM|Other conditions influencing health status|Other conditions influencing health status
C0260724|T033|AB|V49.0|ICD9CM|Deficiencies of limbs|Deficiencies of limbs
C0260724|T033|PT|V49.0|ICD9CM|Deficiencies of limbs|Deficiencies of limbs
C0260725|T033|AB|V49.1|ICD9CM|Mechanical prob w limbs|Mechanical prob w limbs
C0260725|T033|PT|V49.1|ICD9CM|Mechanical problems with limbs|Mechanical problems with limbs
C0260726|T033|AB|V49.2|ICD9CM|Motor problems w limbs|Motor problems w limbs
C0260726|T033|PT|V49.2|ICD9CM|Motor problems with limbs|Motor problems with limbs
C0260727|T033|AB|V49.3|ICD9CM|Sensory problems w limbs|Sensory problems w limbs
C0260727|T033|PT|V49.3|ICD9CM|Sensory problems with limbs|Sensory problems with limbs
C0260728|T033|AB|V49.4|ICD9CM|Disfigurements of limbs|Disfigurements of limbs
C0260728|T033|PT|V49.4|ICD9CM|Disfigurements of limbs|Disfigurements of limbs
C2586328|T033|AB|V49.5|ICD9CM|Limb problems NEC|Limb problems NEC
C2586328|T033|PT|V49.5|ICD9CM|Other problems of limbs|Other problems of limbs
C0376137|T033|HT|V49.6|ICD9CM|Status post amputation of upper limb|Status post amputation of upper limb
C0376138|T033|AB|V49.60|ICD9CM|Status amput up lmb NOS|Status amput up lmb NOS
C0376138|T033|PT|V49.60|ICD9CM|Unspecified level upper limb amputation status|Unspecified level upper limb amputation status
C0376139|T033|AB|V49.61|ICD9CM|Status amput thumb|Status amput thumb
C0376139|T033|PT|V49.61|ICD9CM|Thumb amputation status|Thumb amputation status
C0375854|T033|PT|V49.62|ICD9CM|Other finger(s) amputation status|Other finger(s) amputation status
C0375854|T033|AB|V49.62|ICD9CM|Status amput oth fingers|Status amput oth fingers
C0376140|T033|PT|V49.63|ICD9CM|Hand amputation status|Hand amputation status
C0376140|T033|AB|V49.63|ICD9CM|Status amput hand|Status amput hand
C0376141|T033|AB|V49.64|ICD9CM|Status amput wrist|Status amput wrist
C0376141|T033|PT|V49.64|ICD9CM|Wrist amputation status|Wrist amputation status
C0376142|T033|PT|V49.65|ICD9CM|Below elbow amputation status|Below elbow amputation status
C0376142|T033|AB|V49.65|ICD9CM|Status amput below elbow|Status amput below elbow
C0376143|T033|PT|V49.66|ICD9CM|Above elbow amputation status|Above elbow amputation status
C0376143|T033|AB|V49.66|ICD9CM|Status amput above elbow|Status amput above elbow
C0376144|T033|PT|V49.67|ICD9CM|Shoulder amputation status|Shoulder amputation status
C0376144|T033|AB|V49.67|ICD9CM|Status amput shoulder|Status amput shoulder
C1955601|T033|HT|V49.7|ICD9CM|Lower limb amputation status|Lower limb amputation status
C1955592|T033|AB|V49.70|ICD9CM|Status amput lwr lmb NOS|Status amput lwr lmb NOS
C1955592|T033|PT|V49.70|ICD9CM|Unspecified level lower limb amputation status|Unspecified level lower limb amputation status
C1955593|T033|PT|V49.71|ICD9CM|Great toe amputation status|Great toe amputation status
C1955593|T033|AB|V49.71|ICD9CM|Status amput great toe|Status amput great toe
C1955594|T033|PT|V49.72|ICD9CM|Other toe(s) amputation status|Other toe(s) amputation status
C1955594|T033|AB|V49.72|ICD9CM|Status amput othr toe(s)|Status amput othr toe(s)
C1955595|T033|PT|V49.73|ICD9CM|Foot amputation status|Foot amputation status
C1955595|T033|AB|V49.73|ICD9CM|Status amput foot|Status amput foot
C1955596|T033|PT|V49.74|ICD9CM|Ankle amputation status|Ankle amputation status
C1955596|T033|AB|V49.74|ICD9CM|Status amput ankle|Status amput ankle
C0376124|T033|PT|V49.75|ICD9CM|Below knee amputation status|Below knee amputation status
C0376124|T033|AB|V49.75|ICD9CM|Status amput below knee|Status amput below knee
C0376125|T033|PT|V49.76|ICD9CM|Above knee amputation status|Above knee amputation status
C0376125|T033|AB|V49.76|ICD9CM|Status amput above knee|Status amput above knee
C1955599|T033|PT|V49.77|ICD9CM|Hip amputation status|Hip amputation status
C1955599|T033|AB|V49.77|ICD9CM|Status amput hip|Status amput hip
C0878729|T033|HT|V49.8|ICD9CM|Other specified conditions influencing health status|Other specified conditions influencing health status
C1135338|T033|AB|V49.81|ICD9CM|Asympt postmeno status|Asympt postmeno status
C1135338|T033|PT|V49.81|ICD9CM|Asymptomatic postmenopausal status (age-related) (natural)|Asymptomatic postmenopausal status (age-related) (natural)
C0949155|T033|AB|V49.82|ICD9CM|Dental sealant status|Dental sealant status
C0949155|T033|PT|V49.82|ICD9CM|Dental sealant status|Dental sealant status
C1455976|T033|AB|V49.83|ICD9CM|Await organ transplnt st|Await organ transplnt st
C1455976|T033|PT|V49.83|ICD9CM|Awaiting organ transplant status|Awaiting organ transplant status
C1561676|T033|AB|V49.84|ICD9CM|Bed confinement status|Bed confinement status
C1561676|T033|PT|V49.84|ICD9CM|Bed confinement status|Bed confinement status
C1955602|T033|PT|V49.85|ICD9CM|Dual sensory impairment|Dual sensory impairment
C1955602|T033|AB|V49.85|ICD9CM|Dual sensory impairment|Dual sensory impairment
C0582114|T033|PT|V49.86|ICD9CM|Do not resuscitate status|Do not resuscitate status
C0582114|T033|AB|V49.86|ICD9CM|Do not resusctate status|Do not resusctate status
C2921308|T033|AB|V49.87|ICD9CM|Physical restrain status|Physical restrain status
C2921308|T033|PT|V49.87|ICD9CM|Physical restraints status|Physical restraints status
C0878729|T033|AB|V49.89|ICD9CM|Conditn influ health NEC|Conditn influ health NEC
C0878729|T033|PT|V49.89|ICD9CM|Other specified conditions influencing health status|Other specified conditions influencing health status
C0260729|T033|AB|V49.9|ICD9CM|Probl influ health NOS|Probl influ health NOS
C0260729|T033|PT|V49.9|ICD9CM|Unspecified problems with limbs and other problems|Unspecified problems with limbs and other problems
C0260731|T033|HT|V50|ICD9CM|Elective surgery for purposes other than remedying health states|Elective surgery for purposes other than remedying health states
C0740181|T033|PT|V50.0|ICD9CM|Elective hair transplant for purposes other than remedying health states|Elective hair transplant for purposes other than remedying health states
C0740181|T033|AB|V50.0|ICD9CM|Hair transplant|Hair transplant
C0029711|T033|PT|V50.1|ICD9CM|Other plastic surgery for unacceptable cosmetic appearance|Other plastic surgery for unacceptable cosmetic appearance
C0029711|T033|AB|V50.1|ICD9CM|Plastic surgery NEC|Plastic surgery NEC
C1971613|T033|AB|V50.2|ICD9CM|Routine circumcision|Routine circumcision
C1971613|T033|PT|V50.2|ICD9CM|Routine or ritual circumcision|Routine or ritual circumcision
C0700645|T033|AB|V50.3|ICD9CM|Ear piercing|Ear piercing
C0700645|T033|PT|V50.3|ICD9CM|Ear piercing|Ear piercing
C2910787|T033|PT|V50.41|ICD9CM|Prophylactic breast removal|Prophylactic breast removal
C2910787|T033|AB|V50.41|ICD9CM|Prphylct orgn rmvl brst|Prphylct orgn rmvl brst
C2910788|T033|PT|V50.42|ICD9CM|Prophylactic ovary removal|Prophylactic ovary removal
C2910788|T033|AB|V50.42|ICD9CM|Prphylct orgn rmvl ovary|Prphylct orgn rmvl ovary
C2910789|T033|PT|V50.49|ICD9CM|Other prophylactic gland removal|Other prophylactic gland removal
C2910789|T033|AB|V50.49|ICD9CM|Prphylct orgn rmvl other|Prphylct orgn rmvl other
C0260734|T033|AB|V50.8|ICD9CM|Elective surgery NEC|Elective surgery NEC
C0260734|T033|PT|V50.8|ICD9CM|Other elective surgery for purposes other than remedying health states|Other elective surgery for purposes other than remedying health states
C0260735|T033|AB|V50.9|ICD9CM|Elective surgery NOS|Elective surgery NOS
C0260735|T033|PT|V50.9|ICD9CM|Unspecified elective surgery for purposes other than remedying health states|Unspecified elective surgery for purposes other than remedying health states
C0260736|T033|HT|V51|ICD9CM|Aftercare involving the use of plastic surgery|Aftercare involving the use of plastic surgery
C2349879|T033|AB|V51.0|ICD9CM|Brst reconst fol mastect|Brst reconst fol mastect
C2349879|T033|PT|V51.0|ICD9CM|Encounter for breast reconstruction following mastectomy|Encounter for breast reconstruction following mastectomy
C2349880|T033|AB|V51.8|ICD9CM|Aftercre plastc surg NEC|Aftercre plastc surg NEC
C2349880|T033|PT|V51.8|ICD9CM|Other aftercare involving the use of plastic surgery|Other aftercare involving the use of plastic surgery
C0375859|T033|HT|V52|ICD9CM|Fitting and adjustment of prosthetic device and implant|Fitting and adjustment of prosthetic device and implant
C0260738|T033|PT|V52.0|ICD9CM|Fitting and adjustment of artificial arm (complete) (partial)|Fitting and adjustment of artificial arm (complete) (partial)
C0260738|T033|AB|V52.0|ICD9CM|Fitting artificial arm|Fitting artificial arm
C0260739|T033|PT|V52.1|ICD9CM|Fitting and adjustment of artificial leg (complete) (partial)|Fitting and adjustment of artificial leg (complete) (partial)
C0260739|T033|AB|V52.1|ICD9CM|Fitting artificial leg|Fitting artificial leg
C1971617|T033|PT|V52.2|ICD9CM|Fitting and adjustment of artificial eye|Fitting and adjustment of artificial eye
C1971617|T033|AB|V52.2|ICD9CM|Fitting artificial eye|Fitting artificial eye
C0481749|T033|PT|V52.3|ICD9CM|Fitting and adjustment of dental prosthetic device|Fitting and adjustment of dental prosthetic device
C0481749|T033|AB|V52.3|ICD9CM|Fitting dental prosthes|Fitting dental prosthes
C0375860|T033|AB|V52.4|ICD9CM|Fit/adj breast pros/impl|Fit/adj breast pros/impl
C0375860|T033|PT|V52.4|ICD9CM|Fitting and adjustment of breast prosthesis and implant|Fitting and adjustment of breast prosthesis and implant
C0260743|T033|PT|V52.8|ICD9CM|Fitting and adjustment of other specified prosthetic device|Fitting and adjustment of other specified prosthetic device
C0260743|T033|AB|V52.8|ICD9CM|Fitting prosthesis NEC|Fitting prosthesis NEC
C0260744|T033|PT|V52.9|ICD9CM|Fitting and adjustment of unspecified prosthetic device|Fitting and adjustment of unspecified prosthetic device
C0260744|T033|AB|V52.9|ICD9CM|Fitting prosthesis NOS|Fitting prosthesis NOS
C0260746|T033|HT|V53.0|ICD9CM|Fitting and adjustment of devices related to nervous system and special senses|Fitting and adjustment of devices related to nervous system and special senses
C0490028|T033|AB|V53.01|ICD9CM|Adj cerebral vent shunt|Adj cerebral vent shunt
C0490028|T033|PT|V53.01|ICD9CM|Fitting and adjustment of cerebral ventricular (communicating) shunt|Fitting and adjustment of cerebral ventricular (communicating) shunt
C0490029|T033|AB|V53.02|ICD9CM|Adjust neuropacemaker|Adjust neuropacemaker
C0490029|T033|PT|V53.02|ICD9CM|Fitting and adjustment of neuropacemaker (brain) (peripheral nerve) (spinal cord)|Fitting and adjustment of neuropacemaker (brain) (peripheral nerve) (spinal cord)
C0478576|T033|AB|V53.09|ICD9CM|Adj nerv syst device NEC|Adj nerv syst device NEC
C0478576|T033|PT|V53.09|ICD9CM|Fitting and adjustment of other devices related to nervous system and special senses|Fitting and adjustment of other devices related to nervous system and special senses
C0260747|T033|AB|V53.1|ICD9CM|Fit contact lens/glasses|Fit contact lens/glasses
C0260747|T033|PT|V53.1|ICD9CM|Fitting and adjustment of spectacles and contact lenses|Fitting and adjustment of spectacles and contact lenses
C0260748|T033|AB|V53.2|ICD9CM|Adjustment hearing aid|Adjustment hearing aid
C0260748|T033|PT|V53.2|ICD9CM|Fitting and adjustment of hearing aid|Fitting and adjustment of hearing aid
C0260749|T033|HT|V53.3|ICD9CM|Fitting and adjustment of cardiac pacemaker|Fitting and adjustment of cardiac pacemaker
C0260749|T033|PT|V53.31|ICD9CM|Fitting and adjustment of cardiac pacemaker|Fitting and adjustment of cardiac pacemaker
C0260749|T033|AB|V53.31|ICD9CM|Ftng cardiac pacemaker|Ftng cardiac pacemaker
C0375861|T033|PT|V53.32|ICD9CM|Fitting and adjustment of automatic implantable cardiac defibrillator|Fitting and adjustment of automatic implantable cardiac defibrillator
C0375861|T033|AB|V53.32|ICD9CM|Ftng autmtc dfibrillator|Ftng autmtc dfibrillator
C0375862|T033|PT|V53.39|ICD9CM|Fitting and adjustment of other cardiac device|Fitting and adjustment of other cardiac device
C0375862|T033|AB|V53.39|ICD9CM|Ftng oth cardiac device|Ftng oth cardiac device
C0260750|T033|AB|V53.4|ICD9CM|Fit orthodontic device|Fit orthodontic device
C0260750|T033|PT|V53.4|ICD9CM|Fitting and adjustment of orthodontic devices|Fitting and adjustment of orthodontic devices
C2712802|T033|HT|V53.5|ICD9CM|Fitting and adjustment of other gastrointestinal appliance and device|Fitting and adjustment of other gastrointestinal appliance and device
C2712549|T033|AB|V53.50|ICD9CM|Fit/adjust intestinl dev|Fit/adjust intestinl dev
C2712549|T033|PT|V53.50|ICD9CM|Fitting and adjustment of intestinal appliance and device|Fitting and adjustment of intestinal appliance and device
C2910897|T033|AB|V53.51|ICD9CM|Fit/adj gastric lap band|Fit/adj gastric lap band
C2910897|T033|PT|V53.51|ICD9CM|Fitting and adjustment of gastric lap band|Fitting and adjustment of gastric lap band
C2712802|T033|AB|V53.59|ICD9CM|Fit/adjust gi app-device|Fit/adjust gi app-device
C2712802|T033|PT|V53.59|ICD9CM|Fitting and adjustment of other gastrointestinal appliance and device|Fitting and adjustment of other gastrointestinal appliance and device
C0260752|T033|PT|V53.6|ICD9CM|Fitting and adjustment of urinary devices|Fitting and adjustment of urinary devices
C0260752|T033|AB|V53.6|ICD9CM|Fitting urinary devices|Fitting urinary devices
C0481768|T033|AB|V53.8|ICD9CM|Adjustment of wheelchair|Adjustment of wheelchair
C0481768|T033|PT|V53.8|ICD9CM|Fitting and adjustment of wheelchair|Fitting and adjustment of wheelchair
C0260755|T033|HT|V53.9|ICD9CM|Fitting and adjustment of other and unspecified device|Fitting and adjustment of other and unspecified device
C0496668|T033|AB|V53.90|ICD9CM|Fit/adjust device NOS|Fit/adjust device NOS
C0496668|T033|PT|V53.90|ICD9CM|Fitting and adjustment, unspecified device|Fitting and adjustment, unspecified device
C0260756|T033|HT|V54|ICD9CM|Other orthopedic aftercare|Other orthopedic aftercare
C0260757|T033|HT|V54.0|ICD9CM|Aftercare involving internal fixation device|Aftercare involving internal fixation device
C1260461|T033|PT|V54.01|ICD9CM|Encounter for removal of internal fixation device|Encounter for removal of internal fixation device
C1260461|T033|AB|V54.01|ICD9CM|Removal int fixation dev|Removal int fixation dev
C1135277|T033|HT|V54.1|ICD9CM|Aftercare for healing traumatic fracture|Aftercare for healing traumatic fracture
C1135278|T033|PT|V54.10|ICD9CM|Aftercare for healing traumatic fracture of arm, unspecified|Aftercare for healing traumatic fracture of arm, unspecified
C1135278|T033|AB|V54.10|ICD9CM|Aftrcre traum fx arm NOS|Aftrcre traum fx arm NOS
C1135279|T033|PT|V54.11|ICD9CM|Aftercare for healing traumatic fracture of upper arm|Aftercare for healing traumatic fracture of upper arm
C1135279|T033|AB|V54.11|ICD9CM|Aftrcare traum fx up arm|Aftrcare traum fx up arm
C1135280|T033|PT|V54.12|ICD9CM|Aftercare for healing traumatic fracture of lower arm|Aftercare for healing traumatic fracture of lower arm
C1135280|T033|AB|V54.12|ICD9CM|Aftrcre traum fx low arm|Aftrcre traum fx low arm
C1135281|T033|PT|V54.13|ICD9CM|Aftercare for healing traumatic fracture of hip|Aftercare for healing traumatic fracture of hip
C1135281|T033|AB|V54.13|ICD9CM|Aftrcre traumatic fx hip|Aftrcre traumatic fx hip
C1135282|T033|PT|V54.14|ICD9CM|Aftercare for healing traumatic fracture of leg, unspecified|Aftercare for healing traumatic fracture of leg, unspecified
C1135282|T033|AB|V54.14|ICD9CM|Aftrcre traum fx leg NOS|Aftrcre traum fx leg NOS
C1135283|T033|PT|V54.15|ICD9CM|Aftercare for healing traumatic fracture of upper leg|Aftercare for healing traumatic fracture of upper leg
C1135283|T033|AB|V54.15|ICD9CM|Aftrcare traum fx up leg|Aftrcare traum fx up leg
C1135284|T033|PT|V54.16|ICD9CM|Aftercare for healing traumatic fracture of lower leg|Aftercare for healing traumatic fracture of lower leg
C1135284|T033|AB|V54.16|ICD9CM|Aftrcre traum fx low leg|Aftrcre traum fx low leg
C1135285|T033|PT|V54.17|ICD9CM|Aftercare for healing traumatic fracture of vertebrae|Aftercare for healing traumatic fracture of vertebrae
C1135285|T033|AB|V54.17|ICD9CM|Aftrcre traum fx vertebr|Aftrcre traum fx vertebr
C1135286|T033|PT|V54.19|ICD9CM|Aftercare for healing traumatic fracture of other bone|Aftercare for healing traumatic fracture of other bone
C1135286|T033|AB|V54.19|ICD9CM|Aftrce traum fx bone NEC|Aftrce traum fx bone NEC
C1135287|T033|HT|V54.2|ICD9CM|Aftercare for healing pathologic fracture|Aftercare for healing pathologic fracture
C1135288|T033|PT|V54.20|ICD9CM|Aftercare for healing pathologic fracture of arm, unspecified|Aftercare for healing pathologic fracture of arm, unspecified
C1135288|T033|AB|V54.20|ICD9CM|Aftrcare path fx arm NOS|Aftrcare path fx arm NOS
C1135289|T033|PT|V54.21|ICD9CM|Aftercare for healing pathologic fracture of upper arm|Aftercare for healing pathologic fracture of upper arm
C1135289|T033|AB|V54.21|ICD9CM|Aftercare path fx up arm|Aftercare path fx up arm
C1135290|T033|PT|V54.22|ICD9CM|Aftercare for healing pathologic fracture of lower arm|Aftercare for healing pathologic fracture of lower arm
C1135290|T033|AB|V54.22|ICD9CM|Aftrcare path fx low arm|Aftrcare path fx low arm
C1135291|T033|PT|V54.23|ICD9CM|Aftercare for healing pathologic fracture of hip|Aftercare for healing pathologic fracture of hip
C1135291|T033|AB|V54.23|ICD9CM|Aftercare path fx hip|Aftercare path fx hip
C1135292|T033|PT|V54.24|ICD9CM|Aftercare for healing pathologic fracture of leg, unspecified|Aftercare for healing pathologic fracture of leg, unspecified
C1135292|T033|AB|V54.24|ICD9CM|Aftrcare path fx leg NOS|Aftrcare path fx leg NOS
C1135293|T033|PT|V54.25|ICD9CM|Aftercare for healing pathologic fracture of upper leg|Aftercare for healing pathologic fracture of upper leg
C1135293|T033|AB|V54.25|ICD9CM|Aftrcare path fx up leg|Aftrcare path fx up leg
C1135294|T033|PT|V54.26|ICD9CM|Aftercare for healing pathologic fracture of lower leg|Aftercare for healing pathologic fracture of lower leg
C1135294|T033|AB|V54.26|ICD9CM|Aftrcare path fx low leg|Aftrcare path fx low leg
C1135295|T033|PT|V54.27|ICD9CM|Aftercare for healing pathologic fracture of vertebrae|Aftercare for healing pathologic fracture of vertebrae
C1135295|T033|AB|V54.27|ICD9CM|Aftrcare path fx vertebr|Aftrcare path fx vertebr
C1135296|T033|PT|V54.29|ICD9CM|Aftercare for healing pathologic fracture of other bone|Aftercare for healing pathologic fracture of other bone
C1135296|T033|AB|V54.29|ICD9CM|Aftrcre path fx bone NEC|Aftrcre path fx bone NEC
C0260756|T033|HT|V54.8|ICD9CM|Other orthopedic aftercare|Other orthopedic aftercare
C1135297|T033|PT|V54.81|ICD9CM|Aftercare following joint replacement|Aftercare following joint replacement
C1135297|T033|AB|V54.81|ICD9CM|Aftercare joint replace|Aftercare joint replace
C3161153|T033|AB|V54.82|ICD9CM|Aftcr explantatn jt pros|Aftcr explantatn jt pros
C3161153|T033|PT|V54.82|ICD9CM|Aftercare following explantation of joint prosthesis|Aftercare following explantation of joint prosthesis
C0260756|T033|AB|V54.89|ICD9CM|Orthopedic aftercare NEC|Orthopedic aftercare NEC
C0260756|T033|PT|V54.89|ICD9CM|Other orthopedic aftercare|Other orthopedic aftercare
C0260758|T033|AB|V54.9|ICD9CM|Orthopedic aftercare NOS|Orthopedic aftercare NOS
C0260758|T033|PT|V54.9|ICD9CM|Unspecified orthopedic aftercare|Unspecified orthopedic aftercare
C0740203|T033|HT|V55|ICD9CM|Attention to artificial openings|Attention to artificial openings
C0260760|T033|AB|V55.0|ICD9CM|Atten to tracheostomy|Atten to tracheostomy
C0260760|T033|PT|V55.0|ICD9CM|Attention to tracheostomy|Attention to tracheostomy
C0260761|T033|AB|V55.1|ICD9CM|Atten to gastrostomy|Atten to gastrostomy
C0260761|T033|PT|V55.1|ICD9CM|Attention to gastrostomy|Attention to gastrostomy
C0260762|T033|AB|V55.2|ICD9CM|Atten to ileostomy|Atten to ileostomy
C0260762|T033|PT|V55.2|ICD9CM|Attention to ileostomy|Attention to ileostomy
C0260763|T033|AB|V55.3|ICD9CM|Atten to colostomy|Atten to colostomy
C0260763|T033|PT|V55.3|ICD9CM|Attention to colostomy|Attention to colostomy
C0260764|T033|AB|V55.4|ICD9CM|Atten to enterostomy NEC|Atten to enterostomy NEC
C0260764|T033|PT|V55.4|ICD9CM|Attention to other artificial opening of digestive tract|Attention to other artificial opening of digestive tract
C0260765|T033|AB|V55.5|ICD9CM|Atten to cystostomy|Atten to cystostomy
C0260765|T033|PT|V55.5|ICD9CM|Attention to cystostomy|Attention to cystostomy
C0260766|T033|AB|V55.6|ICD9CM|Atten to urinostomy NEC|Atten to urinostomy NEC
C0260766|T033|PT|V55.6|ICD9CM|Attention to other artificial opening of urinary tract|Attention to other artificial opening of urinary tract
C0260767|T033|AB|V55.7|ICD9CM|Atten artificial vagina|Atten artificial vagina
C0260767|T033|PT|V55.7|ICD9CM|Attention to artificial vagina|Attention to artificial vagina
C0260768|T033|PT|V55.8|ICD9CM|Attention to other specified artificial opening|Attention to other specified artificial opening
C0260768|T033|AB|V55.8|ICD9CM|Attn to artif open NEC|Attn to artif open NEC
C0740203|T033|PT|V55.9|ICD9CM|Attention to unspecified artificial opening|Attention to unspecified artificial opening
C0740203|T033|AB|V55.9|ICD9CM|Attn to artif open NOS|Attn to artif open NOS
C0375864|T033|HT|V56|ICD9CM|Encounter for dialysis and dialysis catheter care|Encounter for dialysis and dialysis catheter care
C0260771|T033|PT|V56.0|ICD9CM|Encounter for extracorporeal dialysis|Encounter for extracorporeal dialysis
C0260771|T033|AB|V56.0|ICD9CM|Renal dialysis encounter|Renal dialysis encounter
C2910939|T033|PT|V56.1|ICD9CM|Fitting and adjustment of extracorporeal dialysis catheter|Fitting and adjustment of extracorporeal dialysis catheter
C2910939|T033|AB|V56.1|ICD9CM|Ft/adj xtrcorp dial cath|Ft/adj xtrcorp dial cath
C2910940|T033|AB|V56.2|ICD9CM|Fit/adj perit dial cath|Fit/adj perit dial cath
C2910940|T033|PT|V56.2|ICD9CM|Fitting and adjustment of peritoneal dialysis catheter|Fitting and adjustment of peritoneal dialysis catheter
C0878730|T033|HT|V56.3|ICD9CM|Encounter for adequacy testing for dialysis|Encounter for adequacy testing for dialysis
C0878731|T033|PT|V56.31|ICD9CM|Encounter for adequacy testing for hemodialysis|Encounter for adequacy testing for hemodialysis
C0878731|T033|AB|V56.31|ICD9CM|Hemodialysis testing|Hemodialysis testing
C0878732|T033|PT|V56.32|ICD9CM|Encounter for adequacy testing for peritoneal dialysis|Encounter for adequacy testing for peritoneal dialysis
C0878732|T033|AB|V56.32|ICD9CM|Peritoneal dialysis test|Peritoneal dialysis test
C0478581|T033|AB|V56.8|ICD9CM|Dialysis encounter, NEC|Dialysis encounter, NEC
C0478581|T033|PT|V56.8|ICD9CM|Encounter for other dialysis|Encounter for other dialysis
C0007237|T033|HT|V57|ICD9CM|Care involving use of rehabilitation procedures|Care involving use of rehabilitation procedures
C0007233|T033|AB|V57.0|ICD9CM|Breathing exercises|Breathing exercises
C0007233|T033|PT|V57.0|ICD9CM|Care involving breathing exercises|Care involving breathing exercises
C0007235|T033|PT|V57.1|ICD9CM|Care involving other physical therapy|Care involving other physical therapy
C0007235|T033|AB|V57.1|ICD9CM|Physical therapy NEC|Physical therapy NEC
C0007234|T033|HT|V57.2|ICD9CM|Care involving occupational therapy and vocational rehabilitation|Care involving occupational therapy and vocational rehabilitation
C1971612|T033|AB|V57.21|ICD9CM|Encntr occupatnal thrpy|Encntr occupatnal thrpy
C1971612|T033|PT|V57.21|ICD9CM|Encounter for occupational therapy|Encounter for occupational therapy
C0375866|T033|AB|V57.22|ICD9CM|Encntr vocational thrpy|Encntr vocational thrpy
C0375866|T033|PT|V57.22|ICD9CM|Encounter for vocational therapy|Encounter for vocational therapy
C0260774|T033|PT|V57.4|ICD9CM|Care involving orthoptic training|Care involving orthoptic training
C0260774|T033|AB|V57.4|ICD9CM|Orthoptic training|Orthoptic training
C0260775|T033|HT|V57.8|ICD9CM|Care involving other specified rehabilitation procedure|Care involving other specified rehabilitation procedure
C0260776|T033|PT|V57.81|ICD9CM|Care involving orthotic training|Care involving orthotic training
C0260776|T033|AB|V57.81|ICD9CM|Orthotic training|Orthotic training
C0260775|T033|PT|V57.89|ICD9CM|Care involving other specified rehabilitation procedure|Care involving other specified rehabilitation procedure
C0260775|T033|AB|V57.89|ICD9CM|Rehabilitation proc NEC|Rehabilitation proc NEC
C0007237|T033|PT|V57.9|ICD9CM|Care involving unspecified rehabilitation procedure|Care involving unspecified rehabilitation procedure
C0007237|T033|AB|V57.9|ICD9CM|Rehabilitation proc NOS|Rehabilitation proc NOS
C0260777|T033|HT|V58|ICD9CM|Encounter for other and unspecified procedures and aftercare|Encounter for other and unspecified procedures and aftercare
C0260778|T033|PT|V58.0|ICD9CM|Encounter for radiotherapy|Encounter for radiotherapy
C0260778|T033|AB|V58.0|ICD9CM|Radiotherapy encounter|Radiotherapy encounter
C0476658|T033|HT|V58.1|ICD9CM|Encounter for antineoplastic chemotherapy and immunotherapy|Encounter for antineoplastic chemotherapy and immunotherapy
C1561677|T033|AB|V58.11|ICD9CM|Antineoplastic chemo enc|Antineoplastic chemo enc
C1561677|T033|PT|V58.11|ICD9CM|Encounter for antineoplastic chemotherapy|Encounter for antineoplastic chemotherapy
C1561678|T033|PT|V58.12|ICD9CM|Encounter for antineoplastic immunotherapy|Encounter for antineoplastic immunotherapy
C1561678|T033|AB|V58.12|ICD9CM|Immunotherapy encounter|Immunotherapy encounter
C0260780|T033|AB|V58.2|ICD9CM|Blood transfusion, no dx|Blood transfusion, no dx
C0260780|T033|PT|V58.2|ICD9CM|Blood transfusion, without reported diagnosis|Blood transfusion, without reported diagnosis
C1719694|T033|HT|V58.3|ICD9CM|Attention to dressings and sutures|Attention to dressings and sutures
C1719690|T033|AB|V58.30|ICD9CM|Attn rem nonsurg dressng|Attn rem nonsurg dressng
C1719690|T033|PT|V58.30|ICD9CM|Encounter for change or removal of nonsurgical wound dressing|Encounter for change or removal of nonsurgical wound dressing
C1719692|T033|AB|V58.31|ICD9CM|Attn rem surg dressing|Attn rem surg dressing
C1719692|T033|PT|V58.31|ICD9CM|Encounter for change or removal of surgical wound dressing|Encounter for change or removal of surgical wound dressing
C1719693|T033|AB|V58.32|ICD9CM|Attn removal of sutures|Attn removal of sutures
C1719693|T033|PT|V58.32|ICD9CM|Encounter for removal of sutures|Encounter for removal of sutures
C0260782|T033|HT|V58.4|ICD9CM|Other aftercare following surgery|Other aftercare following surgery
C0375867|T033|AB|V58.41|ICD9CM|Encntr plnd po wnd clsr|Encntr plnd po wnd clsr
C0375867|T033|PT|V58.41|ICD9CM|Encounter for planned post-operative wound closure|Encounter for planned post-operative wound closure
C1135298|T033|PT|V58.42|ICD9CM|Aftercare following surgery for neoplasm|Aftercare following surgery for neoplasm
C1135298|T033|AB|V58.42|ICD9CM|Aftercare neoplasm surg|Aftercare neoplasm surg
C1135299|T033|PT|V58.43|ICD9CM|Aftercare following surgery for injury and trauma|Aftercare following surgery for injury and trauma
C1135299|T033|AB|V58.43|ICD9CM|Aftrcare inj/trauma surg|Aftrcare inj/trauma surg
C0375868|T033|PT|V58.49|ICD9CM|Other specified aftercare following surgery|Other specified aftercare following surgery
C0375868|T033|AB|V58.49|ICD9CM|Postop oth specfd aftrcr|Postop oth specfd aftrcr
C0029336|T033|AB|V58.5|ICD9CM|Orthodontics aftercare|Orthodontics aftercare
C0029336|T033|PT|V58.5|ICD9CM|Orthodontics aftercare|Orthodontics aftercare
C0375869|T033|HT|V58.6|ICD9CM|Encounter for long-term (current) drug use|Encounter for long-term (current) drug use
C2911178|T033|PT|V58.61|ICD9CM|Long-term (current) use of anticoagulants|Long-term (current) use of anticoagulants
C2911178|T033|AB|V58.61|ICD9CM|Long-term use anticoagul|Long-term use anticoagul
C2911181|T033|PT|V58.62|ICD9CM|Long-term (current) use of antibiotics|Long-term (current) use of antibiotics
C2911181|T033|AB|V58.62|ICD9CM|Long-term use antibiotic|Long-term use antibiotic
C2911179|T033|AB|V58.63|ICD9CM|Lng use antiplte/thrmbtc|Lng use antiplte/thrmbtc
C2911179|T033|PT|V58.63|ICD9CM|Long-term (current) use of antiplatelet/antithrombotic|Long-term (current) use of antiplatelet/antithrombotic
C2911180|T033|PT|V58.64|ICD9CM|Long-term (current) use of non-steroidal anti-inflammatories (NSAID)|Long-term (current) use of non-steroidal anti-inflammatories (NSAID)
C2911180|T033|AB|V58.64|ICD9CM|Long-term anti-inflamtry|Long-term anti-inflamtry
C1260466|T033|PT|V58.65|ICD9CM|Long-term (current) use of steroids|Long-term (current) use of steroids
C1260466|T033|AB|V58.65|ICD9CM|Long-term use steroids|Long-term use steroids
C2911205|T033|PT|V58.66|ICD9CM|Long-term (current) use of aspirin|Long-term (current) use of aspirin
C2911205|T033|AB|V58.66|ICD9CM|Long-term use of aspirin|Long-term use of aspirin
C1455979|T033|PT|V58.67|ICD9CM|Long-term (current) use of insulin|Long-term (current) use of insulin
C1455979|T033|AB|V58.67|ICD9CM|Long-term use of insulin|Long-term use of insulin
C3161154|T033|AB|V58.68|ICD9CM|Lng term bisphosphonates|Lng term bisphosphonates
C3161154|T033|PT|V58.68|ICD9CM|Long term (current) use of bisphosphonates|Long term (current) use of bisphosphonates
C0375871|T033|PT|V58.69|ICD9CM|Long-term (current) use of other medications|Long-term (current) use of other medications
C0375871|T033|AB|V58.69|ICD9CM|Long-term use meds NEC|Long-term use meds NEC
C1135300|T033|HT|V58.7|ICD9CM|Aftercare following surgery to specified body systems, not elsewhere classified|Aftercare following surgery to specified body systems, not elsewhere classified
C1135301|T033|AB|V58.71|ICD9CM|Aft surg sense org NEC|Aft surg sense org NEC
C1135301|T033|PT|V58.71|ICD9CM|Aftercare following surgery of the sense organs, NEC|Aftercare following surgery of the sense organs, NEC
C1135302|T033|AB|V58.72|ICD9CM|Aftcre surg nerv sys NEC|Aftcre surg nerv sys NEC
C1135302|T033|PT|V58.72|ICD9CM|Aftercare following surgery of the nervous system, NEC|Aftercare following surgery of the nervous system, NEC
C1135303|T033|AB|V58.73|ICD9CM|Aft surg circ syst NEC|Aft surg circ syst NEC
C1135303|T033|PT|V58.73|ICD9CM|Aftercare following surgery of the circulatory system, NEC|Aftercare following surgery of the circulatory system, NEC
C1135304|T033|PT|V58.74|ICD9CM|Aftercare following surgery of the respiratory system, NEC|Aftercare following surgery of the respiratory system, NEC
C1135304|T033|AB|V58.74|ICD9CM|Aftrcre surg respsys NEC|Aftrcre surg respsys NEC
C1135305|T033|AB|V58.75|ICD9CM|Aft oral cav/dig sys NEC|Aft oral cav/dig sys NEC
C1135305|T033|PT|V58.75|ICD9CM|Aftercare following surgery of the teeth, oral cavity and digestive system, NEC|Aftercare following surgery of the teeth, oral cavity and digestive system, NEC
C1135306|T033|PT|V58.76|ICD9CM|Aftercare following surgery of the genitourinary system, NEC|Aftercare following surgery of the genitourinary system, NEC
C1135306|T033|AB|V58.76|ICD9CM|Aftrcre surg GU syst NEC|Aftrcre surg GU syst NEC
C1135307|T033|AB|V58.77|ICD9CM|Aft surg skin/subcu NEC|Aft surg skin/subcu NEC
C1135307|T033|PT|V58.77|ICD9CM|Aftercare following surgery of the skin and subcutaneous tissue, NEC|Aftercare following surgery of the skin and subcutaneous tissue, NEC
C1135308|T033|PT|V58.78|ICD9CM|Aftercare following surgery of the musculoskeletal system, NEC|Aftercare following surgery of the musculoskeletal system, NEC
C1135308|T033|AB|V58.78|ICD9CM|Aftrcre surg MS syst NEC|Aftrcre surg MS syst NEC
C0375872|T033|HT|V58.8|ICD9CM|Encounter for other specified procedures and aftercare|Encounter for other specified procedures and aftercare
C0375873|T033|AB|V58.81|ICD9CM|Fit/adj vascular cathetr|Fit/adj vascular cathetr
C0375873|T033|PT|V58.81|ICD9CM|Fitting and adjustment of vascular catheter|Fitting and adjustment of vascular catheter
C0375874|T033|AB|V58.82|ICD9CM|Fit/adj non-vsc cath NEC|Fit/adj non-vsc cath NEC
C0375874|T033|PT|V58.82|ICD9CM|Fitting and adjustment of nonvascular catheter, NEC|Fitting and adjustment of nonvascular catheter, NEC
C2910943|T033|PT|V58.83|ICD9CM|Encounter for therapeutic drug monitoring|Encounter for therapeutic drug monitoring
C2910943|T033|AB|V58.83|ICD9CM|Therapeutic drug monitor|Therapeutic drug monitor
C0260783|T033|AB|V58.89|ICD9CM|Other specfied aftercare|Other specfied aftercare
C0260783|T033|PT|V58.89|ICD9CM|Other specified aftercare|Other specified aftercare
C0260784|T033|AB|V58.9|ICD9CM|Aftercare NOS|Aftercare NOS
C0260784|T033|PT|V58.9|ICD9CM|Unspecified aftercare|Unspecified aftercare
C1527169|T033|HT|V59|ICD9CM|Donors|Donors
C1313951|T033|HT|V59.0|ICD9CM|Blood donors|Blood donors
C2830121|T033|AB|V59.01|ICD9CM|Blood donor-whole blood|Blood donor-whole blood
C2830121|T033|PT|V59.01|ICD9CM|Blood donors, whole blood|Blood donors, whole blood
C2830119|T033|AB|V59.02|ICD9CM|Blood donor-stem cells|Blood donor-stem cells
C2830119|T033|PT|V59.02|ICD9CM|Blood donors, stem cells|Blood donors, stem cells
C0375878|T033|AB|V59.09|ICD9CM|Blood donor NEC|Blood donor NEC
C0375878|T033|PT|V59.09|ICD9CM|Other blood donors|Other blood donors
C0260785|T033|AB|V59.1|ICD9CM|Skin donor|Skin donor
C0260785|T033|PT|V59.1|ICD9CM|Skin donors|Skin donors
C1313933|T033|AB|V59.2|ICD9CM|Bone donor|Bone donor
C1313933|T033|PT|V59.2|ICD9CM|Bone donors|Bone donors
C1313934|T033|AB|V59.3|ICD9CM|Bone marrow donor|Bone marrow donor
C1313934|T033|PT|V59.3|ICD9CM|Bone marrow donors|Bone marrow donors
C1313935|T033|AB|V59.4|ICD9CM|Kidney donor|Kidney donor
C1313935|T033|PT|V59.4|ICD9CM|Kidney donors|Kidney donors
C0260789|T033|AB|V59.5|ICD9CM|Cornea donor|Cornea donor
C0260789|T033|PT|V59.5|ICD9CM|Cornea donors|Cornea donors
C2830120|T033|AB|V59.6|ICD9CM|Liver donor|Liver donor
C2830120|T033|PT|V59.6|ICD9CM|Liver donors|Liver donors
C1561686|T033|HT|V59.7|ICD9CM|Egg (oocyte) (ovum)|Egg (oocyte) (ovum)
C2910967|T033|PT|V59.70|ICD9CM|Egg (oocyte) (ovum) donor, unspecified|Egg (oocyte) (ovum) donor, unspecified
C2910967|T033|AB|V59.70|ICD9CM|Egg donor NEC|Egg donor NEC
C1561680|T033|PT|V59.71|ICD9CM|Egg (oocyte) (ovum) donor, under age 35, anonymous recipient|Egg (oocyte) (ovum) donor, under age 35, anonymous recipient
C1561680|T033|AB|V59.71|ICD9CM|Egg donor age <35 anon|Egg donor age <35 anon
C2910964|T033|PT|V59.72|ICD9CM|Egg (oocyte) (ovum) donor, under age 35, designated recipient|Egg (oocyte) (ovum) donor, under age 35, designated recipient
C2910964|T033|AB|V59.72|ICD9CM|Egg donor age <35 desig|Egg donor age <35 desig
C1561683|T033|PT|V59.73|ICD9CM|Egg (oocyte) (ovum) donor, age 35 and over, anonymous recipient|Egg (oocyte) (ovum) donor, age 35 and over, anonymous recipient
C1561683|T033|AB|V59.73|ICD9CM|Egg donor age 35+ anon|Egg donor age 35+ anon
C2910966|T033|PT|V59.74|ICD9CM|Egg (oocyte) (ovum) donor, age 35 and over, designated recipient|Egg (oocyte) (ovum) donor, age 35 and over, designated recipient
C2910966|T033|AB|V59.74|ICD9CM|Egg donor age 35+ desig|Egg donor age 35+ desig
C0260790|T033|PT|V59.8|ICD9CM|Donors of other specified organ or tissue|Donors of other specified organ or tissue
C0260790|T033|AB|V59.8|ICD9CM|Org or tissue donor NEC|Org or tissue donor NEC
C0013019|T033|PT|V59.9|ICD9CM|Donors of unspecified organ or tissue|Donors of unspecified organ or tissue
C0013019|T033|AB|V59.9|ICD9CM|Org or tissue donor NOS|Org or tissue donor NOS
C0260791|T033|HT|V60|ICD9CM|Housing, household, and economic circumstances|Housing, household, and economic circumstances
C0178343|T033|HT|V60-V69.99|ICD9CM|PERSONS ENCOUNTERING HEALTH SERVICES IN OTHER CIRCUMSTANCES|PERSONS ENCOUNTERING HEALTH SERVICES IN OTHER CIRCUMSTANCES
C0687129|T033|AB|V60.0|ICD9CM|Lack of housing|Lack of housing
C0687129|T033|PT|V60.0|ICD9CM|Lack of housing|Lack of housing
C0260793|T033|AB|V60.1|ICD9CM|Inadequate housing|Inadequate housing
C0260793|T033|PT|V60.1|ICD9CM|Inadequate housing|Inadequate housing
C0021138|T033|AB|V60.2|ICD9CM|Economic problem|Economic problem
C0021138|T033|PT|V60.2|ICD9CM|Inadequate material resources|Inadequate material resources
C0260794|T033|AB|V60.3|ICD9CM|Person living alone|Person living alone
C0260794|T033|PT|V60.3|ICD9CM|Person living alone|Person living alone
C0260795|T033|AB|V60.4|ICD9CM|No family able to care|No family able to care
C0260795|T033|PT|V60.4|ICD9CM|No other household member able to render care|No other household member able to render care
C0260796|T033|AB|V60.5|ICD9CM|Holiday relief care|Holiday relief care
C0260796|T033|PT|V60.5|ICD9CM|Holiday relief care|Holiday relief care
C0260797|T033|AB|V60.6|ICD9CM|Person in resident inst|Person in resident inst
C0260797|T033|PT|V60.6|ICD9CM|Person living in residential institution|Person living in residential institution
C0260798|T033|HT|V60.8|ICD9CM|Other specified housing or economic circumstances|Other specified housing or economic circumstances
C2712551|T033|AB|V60.81|ICD9CM|Foster care (status)|Foster care (status)
C2712551|T033|PT|V60.81|ICD9CM|Foster care (status)|Foster care (status)
C2712997|T033|AB|V60.89|ICD9CM|Housing/econo circum NEC|Housing/econo circum NEC
C2712997|T033|PT|V60.89|ICD9CM|Other specified housing or economic circumstances|Other specified housing or economic circumstances
C0260799|T033|AB|V60.9|ICD9CM|Housing/econo circum NOS|Housing/econo circum NOS
C0260799|T033|PT|V60.9|ICD9CM|Unspecified housing or economic circumstance|Unspecified housing or economic circumstance
C0481797|T033|HT|V61|ICD9CM|Other family circumstances|Other family circumstances
C0481798|T033|HT|V61.0|ICD9CM|Family disruption|Family disruption
C2349886|T033|PT|V61.01|ICD9CM|Family disruption due to family member on military deployment|Family disruption due to family member on military deployment
C2349886|T033|AB|V61.01|ICD9CM|Fmily dsrpt-fam military|Fmily dsrpt-fam military
C2349888|T033|PT|V61.02|ICD9CM|Family disruption due to return of family member from military deployment|Family disruption due to return of family member from military deployment
C2349888|T033|AB|V61.02|ICD9CM|Fmily dsrpt-ret military|Fmily dsrpt-ret military
C2349890|T033|PT|V61.03|ICD9CM|Family disruption due to divorce or legal separation|Family disruption due to divorce or legal separation
C2349890|T033|AB|V61.03|ICD9CM|Fmily dsrpt- divorce/sep|Fmily dsrpt- divorce/sep
C2349891|T033|PT|V61.04|ICD9CM|Family disruption due to parent-child estrangement|Family disruption due to parent-child estrangement
C2349891|T033|AB|V61.04|ICD9CM|Family dsrpt-estrangmemt|Family dsrpt-estrangmemt
C2349892|T033|PT|V61.05|ICD9CM|Family disruption due to child in welfare custody|Family disruption due to child in welfare custody
C2349892|T033|AB|V61.05|ICD9CM|Famly dsrpt-chld custody|Famly dsrpt-chld custody
C2349893|T033|PT|V61.06|ICD9CM|Family disruption due to child in foster care or in care of non-parental family member|Family disruption due to child in foster care or in care of non-parental family member
C2349893|T033|AB|V61.06|ICD9CM|Family dsrpt-foster care|Family dsrpt-foster care
C2712552|T033|PT|V61.07|ICD9CM|Family disruption due to death of family member|Family disruption due to death of family member
C2712552|T033|AB|V61.07|ICD9CM|Family dsrpt-death membr|Family dsrpt-death membr
C2712553|T033|PT|V61.08|ICD9CM|Family disruption due to other extended absence of family member|Family disruption due to other extended absence of family member
C2712553|T033|AB|V61.08|ICD9CM|Fmly dsrp-fam absnce NEC|Fmly dsrp-fam absnce NEC
C2349894|T033|AB|V61.09|ICD9CM|Family disruption NEC|Family disruption NEC
C2349894|T033|PT|V61.09|ICD9CM|Other family disruption|Other family disruption
C0375879|T033|HT|V61.1|ICD9CM|Counseling for marital and partner problems|Counseling for marital and partner problems
C0375880|T033|AB|V61.10|ICD9CM|Consl partner prob|Consl partner prob
C0375880|T033|PT|V61.10|ICD9CM|Counseling for marital and partner problems, unspecified|Counseling for marital and partner problems, unspecified
C2911077|T033|AB|V61.11|ICD9CM|Cnsl victm partner abuse|Cnsl victm partner abuse
C2911077|T033|PT|V61.11|ICD9CM|Counseling for victim of spousal and partner abuse|Counseling for victim of spousal and partner abuse
C0795786|T033|AB|V61.12|ICD9CM|Cnsl perp partner abuse|Cnsl perp partner abuse
C0795786|T033|PT|V61.12|ICD9CM|Counseling for perpetrator of spousal and partner abuse|Counseling for perpetrator of spousal and partner abuse
C0700498|T033|HT|V61.2|ICD9CM|Parent-child problems|Parent-child problems
C0375882|T033|AB|V61.20|ICD9CM|Cnsl prnt-chld prob NOS|Cnsl prnt-chld prob NOS
C0375882|T033|PT|V61.20|ICD9CM|Counseling for parent-child problem, unspecified|Counseling for parent-child problem, unspecified
C0375883|T033|AB|V61.21|ICD9CM|Cnsl victim child abuse|Cnsl victim child abuse
C0375883|T033|PT|V61.21|ICD9CM|Counseling for victim of child abuse|Counseling for victim of child abuse
C0795786|T033|AB|V61.22|ICD9CM|Cnsl perp parent chld ab|Cnsl perp parent chld ab
C0795786|T033|PT|V61.22|ICD9CM|Counseling for perpetrator of spousal and partner abuse|Counseling for perpetrator of spousal and partner abuse
C2712554|T033|AB|V61.23|ICD9CM|Cnsl prnt-biol chld prob|Cnsl prnt-biol chld prob
C2712554|T033|PT|V61.23|ICD9CM|Counseling for parent-biological child problem|Counseling for parent-biological child problem
C2712555|T033|AB|V61.24|ICD9CM|Cnsl prnt-adpt chld prob|Cnsl prnt-adpt chld prob
C2712555|T033|PT|V61.24|ICD9CM|Counseling for parent-adopted child problem|Counseling for parent-adopted child problem
C2712556|T033|AB|V61.25|ICD9CM|Cnsl prnt-fstr chld prob|Cnsl prnt-fstr chld prob
C2712556|T033|PT|V61.25|ICD9CM|Counseling for parent (guardian)-foster child problem|Counseling for parent (guardian)-foster child problem
C0029699|T033|AB|V61.29|ICD9CM|Oth parent-child problem|Oth parent-child problem
C0029699|T033|PT|V61.29|ICD9CM|Other parent-child problems|Other parent-child problems
C0260801|T033|AB|V61.3|ICD9CM|Problem w aged parent|Problem w aged parent
C0260801|T033|PT|V61.3|ICD9CM|Problems with aged parents or in-laws|Problems with aged parents or in-laws
C0481514|T033|HT|V61.4|ICD9CM|Health problems within family|Health problems within family
C0476560|T033|AB|V61.41|ICD9CM|Alcoholism in family|Alcoholism in family
C0476560|T033|PT|V61.41|ICD9CM|Alcoholism in family|Alcoholism in family
C2712557|T033|PT|V61.42|ICD9CM|Substance abuse in family|Substance abuse in family
C2712557|T033|AB|V61.42|ICD9CM|Substance abuse-family|Substance abuse-family
C0260804|T033|AB|V61.49|ICD9CM|Family health probl NEC|Family health probl NEC
C0260804|T033|PT|V61.49|ICD9CM|Other health problems within the family|Other health problems within the family
C0700322|T033|AB|V61.5|ICD9CM|Multiparity|Multiparity
C0700322|T033|PT|V61.5|ICD9CM|Multiparity|Multiparity
C1313860|T033|PT|V61.6|ICD9CM|Illegitimacy or illegitimate pregnancy|Illegitimacy or illegitimate pregnancy
C1313860|T033|AB|V61.6|ICD9CM|Illegitimate pregnancy|Illegitimate pregnancy
C0029865|T033|PT|V61.7|ICD9CM|Other unwanted pregnancy|Other unwanted pregnancy
C0029865|T033|AB|V61.7|ICD9CM|Unwanted pregnancy NEC|Unwanted pregnancy NEC
C0481799|T033|AB|V61.8|ICD9CM|Family circumstances NEC|Family circumstances NEC
C0481799|T033|PT|V61.8|ICD9CM|Other specified family circumstances|Other specified family circumstances
C0029795|T033|AB|V61.9|ICD9CM|Family circumstance NOS|Family circumstance NOS
C0029795|T033|PT|V61.9|ICD9CM|Unspecified family circumstance|Unspecified family circumstance
C0260805|T033|HT|V62|ICD9CM|Other psychosocial circumstances|Other psychosocial circumstances
C0496682|T033|AB|V62.0|ICD9CM|Unemployment|Unemployment
C0496682|T033|PT|V62.0|ICD9CM|Unemployment|Unemployment
C0260806|T033|AB|V62.1|ICD9CM|Adverse eff-work environ|Adverse eff-work environ
C0260806|T033|PT|V62.1|ICD9CM|Adverse effects of work environment|Adverse effects of work environment
C0029680|T033|HT|V62.2|ICD9CM|Other occupational circumstances or maladjustment|Other occupational circumstances or maladjustment
C2349895|T033|AB|V62.21|ICD9CM|Hx military deployment|Hx military deployment
C2349895|T033|PT|V62.21|ICD9CM|Personal current military deployment status|Personal current military deployment status
C2349897|T033|AB|V62.22|ICD9CM|Hx retrn military deploy|Hx retrn military deploy
C2349897|T033|PT|V62.22|ICD9CM|Personal history of return from military deployment|Personal history of return from military deployment
C0029680|T033|AB|V62.29|ICD9CM|Occupationl circumst NEC|Occupationl circumst NEC
C0029680|T033|PT|V62.29|ICD9CM|Other occupational circumstances or maladjustment|Other occupational circumstances or maladjustment
C0013654|T033|AB|V62.3|ICD9CM|Educational circumstance|Educational circumstance
C0013654|T033|PT|V62.3|ICD9CM|Educational circumstances|Educational circumstances
C0677639|T033|AB|V62.4|ICD9CM|Social maladjustment|Social maladjustment
C0677639|T033|PT|V62.4|ICD9CM|Social maladjustment|Social maladjustment
C0260807|T033|AB|V62.5|ICD9CM|Legal circumstances|Legal circumstances
C0260807|T033|PT|V62.5|ICD9CM|Legal circumstances|Legal circumstances
C0080099|T033|AB|V62.6|ICD9CM|Refusal of treatment|Refusal of treatment
C0080099|T033|PT|V62.6|ICD9CM|Refusal of treatment for reasons of religion or conscience|Refusal of treatment for reasons of religion or conscience
C0302431|T033|HT|V62.8|ICD9CM|Other psychological or physical stress, not elsewhere classified|Other psychological or physical stress, not elsewhere classified
C0869289|T033|AB|V62.81|ICD9CM|Interpersonal probl NEC|Interpersonal probl NEC
C0869289|T033|PT|V62.81|ICD9CM|Interpersonal problems, not elsewhere classified|Interpersonal problems, not elsewhere classified
C0684255|T033|AB|V62.82|ICD9CM|Bereavement, uncomplicat|Bereavement, uncomplicat
C0684255|T033|PT|V62.82|ICD9CM|Bereavement, uncomplicated|Bereavement, uncomplicated
C0375885|T033|AB|V62.83|ICD9CM|Cnsl perp phys/sex abuse|Cnsl perp phys/sex abuse
C0375885|T033|PT|V62.83|ICD9CM|Counseling for perpetrator of physical/sexual abuse|Counseling for perpetrator of physical/sexual abuse
C0424000|T033|AB|V62.84|ICD9CM|Suicidal ideation|Suicidal ideation
C0424000|T033|PT|V62.84|ICD9CM|Suicidal ideation|Suicidal ideation
C0455204|T033|AB|V62.85|ICD9CM|Homicidal ideation|Homicidal ideation
C0455204|T033|PT|V62.85|ICD9CM|Homicidal ideation|Homicidal ideation
C0302431|T033|PT|V62.89|ICD9CM|Other psychological or physical stress, not elsewhere classified|Other psychological or physical stress, not elsewhere classified
C0302431|T033|AB|V62.89|ICD9CM|Psychological stress NEC|Psychological stress NEC
C0260808|T033|AB|V62.9|ICD9CM|Psychosocial circum NOS|Psychosocial circum NOS
C0260808|T033|PT|V62.9|ICD9CM|Unspecified psychosocial circumstance|Unspecified psychosocial circumstance
C0260809|T033|HT|V63|ICD9CM|Unavailability of other medical facilities for care|Unavailability of other medical facilities for care
C0260810|T033|AB|V63.0|ICD9CM|Home remote from hospitl|Home remote from hospitl
C0260810|T033|PT|V63.0|ICD9CM|Residence remote from hospital or other health care facility|Residence remote from hospital or other health care facility
C0420585|T033|PT|V63.1|ICD9CM|Medical services in home not available|Medical services in home not available
C0420585|T033|AB|V63.1|ICD9CM|No medical serv in home|No medical serv in home
C0260812|T033|PT|V63.2|ICD9CM|Person awaiting admission to adequate facility elsewhere|Person awaiting admission to adequate facility elsewhere
C0260812|T033|AB|V63.2|ICD9CM|Wait adm to oth facility|Wait adm to oth facility
C0260813|T033|AB|V63.8|ICD9CM|No med facilities NEC|No med facilities NEC
C0260813|T033|PT|V63.8|ICD9CM|Other specified reasons for unavailability of medical facilities|Other specified reasons for unavailability of medical facilities
C0260814|T033|AB|V63.9|ICD9CM|No med facilities NOS|No med facilities NOS
C0260814|T033|PT|V63.9|ICD9CM|Unspecified reason for unavailability of medical facilities|Unspecified reason for unavailability of medical facilities
C0260815|T033|HT|V64|ICD9CM|Persons encountering health services for specific procedures, not carried out|Persons encountering health services for specific procedures, not carried out
C2919035|T033|HT|V64.0|ICD9CM|Vaccination not carried out|Vaccination not carried out
C0476665|T033|AB|V64.00|ICD9CM|No vaccination NOS|No vaccination NOS
C0476665|T033|PT|V64.00|ICD9CM|Vaccination not carried out, unspecified reason|Vaccination not carried out, unspecified reason
C2910670|T033|AB|V64.01|ICD9CM|No vaccin-acute illness|No vaccin-acute illness
C2910670|T033|PT|V64.01|ICD9CM|Vaccination not carried out because of acute illness|Vaccination not carried out because of acute illness
C2910671|T033|AB|V64.02|ICD9CM|No vaccin-chronc illness|No vaccin-chronc illness
C2910671|T033|PT|V64.02|ICD9CM|Vaccination not carried out because of chronic illness or condition|Vaccination not carried out because of chronic illness or condition
C2910672|T033|AB|V64.03|ICD9CM|No vaccin-immune comp|No vaccin-immune comp
C2910672|T033|PT|V64.03|ICD9CM|Vaccination not carried out because of immune compromised state|Vaccination not carried out because of immune compromised state
C1561694|T033|AB|V64.04|ICD9CM|No vaccin-allergy to vac|No vaccin-allergy to vac
C1561694|T033|PT|V64.04|ICD9CM|Vaccination not carried out because of allergy to vaccine or component|Vaccination not carried out because of allergy to vaccine or component
C1561695|T033|AB|V64.05|ICD9CM|No vaccin-caregiv refuse|No vaccin-caregiv refuse
C1561695|T033|PT|V64.05|ICD9CM|Vaccination not carried out because of caregiver refusal|Vaccination not carried out because of caregiver refusal
C1561696|T033|AB|V64.06|ICD9CM|No vaccination-pt refuse|No vaccination-pt refuse
C1561696|T033|PT|V64.06|ICD9CM|Vaccination not carried out because of patient refusal|Vaccination not carried out because of patient refusal
C1561697|T033|AB|V64.07|ICD9CM|No vaccination-religion|No vaccination-religion
C1561697|T033|PT|V64.07|ICD9CM|Vaccination not carried out for religious reasons|Vaccination not carried out for religious reasons
C1561698|T033|AB|V64.08|ICD9CM|No vaccin-prev disease|No vaccin-prev disease
C1561698|T033|PT|V64.08|ICD9CM|Vaccination not carried out because patient had disease being vaccinated against|Vaccination not carried out because patient had disease being vaccinated against
C0476664|T033|AB|V64.09|ICD9CM|No vaccination NEC|No vaccination NEC
C0476664|T033|PT|V64.09|ICD9CM|Vaccination not carried out for other reason|Vaccination not carried out for other reason
C0260817|T033|AB|V64.1|ICD9CM|No proc/contraindication|No proc/contraindication
C0260817|T033|PT|V64.1|ICD9CM|Surgical or other procedure not carried out because of contraindication|Surgical or other procedure not carried out because of contraindication
C0260818|T033|AB|V64.2|ICD9CM|No proc/patient decision|No proc/patient decision
C0260818|T033|PT|V64.2|ICD9CM|Surgical or other procedure not carried out because of patient's decision|Surgical or other procedure not carried out because of patient's decision
C0260819|T033|AB|V64.3|ICD9CM|No proc for reasons NEC|No proc for reasons NEC
C0260819|T033|PT|V64.3|ICD9CM|Procedure not carried out for other reasons|Procedure not carried out for other reasons
C0490030|T033|HT|V64.4|ICD9CM|Closed surgical procedure converted to open procedure|Closed surgical procedure converted to open procedure
C1260467|T033|AB|V64.41|ICD9CM|Lap surg convert to open|Lap surg convert to open
C1260467|T033|PT|V64.41|ICD9CM|Laparoscopic surgical procedure converted to open procedure|Laparoscopic surgical procedure converted to open procedure
C1260468|T033|AB|V64.42|ICD9CM|Thoracoscop conv to open|Thoracoscop conv to open
C1260468|T033|PT|V64.42|ICD9CM|Thoracoscopic surgical procedure converted to open procedure|Thoracoscopic surgical procedure converted to open procedure
C1260469|T033|AB|V64.43|ICD9CM|Arthroscopc conv to open|Arthroscopc conv to open
C1260469|T033|PT|V64.43|ICD9CM|Arthroscopic surgical procedure converted to open procedure|Arthroscopic surgical procedure converted to open procedure
C0260820|T033|HT|V65|ICD9CM|Other persons seeking consultation|Other persons seeking consultation
C0260821|T033|PT|V65.0|ICD9CM|Healthy person accompanying sick person|Healthy person accompanying sick person
C0260821|T033|AB|V65.0|ICD9CM|Healthy person w sick|Healthy person w sick
C0260822|T033|HT|V65.1|ICD9CM|Person consulting on behalf of another person|Person consulting on behalf of another person
C2911138|T033|AB|V65.11|ICD9CM|Ped pre-brth vst-parent|Ped pre-brth vst-parent
C2911138|T033|PT|V65.11|ICD9CM|Pediatric pre-birth visit for expectant parent(s)|Pediatric pre-birth visit for expectant parent(s)
C0496703|T033|AB|V65.2|ICD9CM|Person feigning illness|Person feigning illness
C0496703|T033|PT|V65.2|ICD9CM|Person feigning illness|Person feigning illness
C0260823|T033|AB|V65.3|ICD9CM|Dietary surveil/counsel|Dietary surveil/counsel
C0260823|T033|PT|V65.3|ICD9CM|Dietary surveillance and counseling|Dietary surveillance and counseling
C0869481|T033|HT|V65.4|ICD9CM|Other counseling, not elsewhere classified|Other counseling, not elsewhere classified
C0740209|T033|AB|V65.40|ICD9CM|Counseling NOS|Counseling NOS
C0740209|T033|PT|V65.40|ICD9CM|Counseling NOS|Counseling NOS
C0375886|T033|AB|V65.41|ICD9CM|Exercise counseling|Exercise counseling
C0375886|T033|PT|V65.41|ICD9CM|Exercise counseling|Exercise counseling
C0375888|T033|AB|V65.43|ICD9CM|Counseling injry prevent|Counseling injry prevent
C0375888|T033|PT|V65.43|ICD9CM|Counseling on injury prevention|Counseling on injury prevention
C0476681|T033|AB|V65.44|ICD9CM|Hiv counseling|Hiv counseling
C0476681|T033|PT|V65.44|ICD9CM|Human immunodeficiency virus (HIV) counseling|Human immunodeficiency virus (HIV) counseling
C0375890|T033|AB|V65.45|ICD9CM|Consln ot sex trnsmt dis|Consln ot sex trnsmt dis
C0375890|T033|PT|V65.45|ICD9CM|Counseling on other sexually transmitted diseases|Counseling on other sexually transmitted diseases
C0348773|T033|AB|V65.49|ICD9CM|Other specfd counseling|Other specfd counseling
C0348773|T033|PT|V65.49|ICD9CM|Other specified counseling|Other specified counseling
C0851311|T033|AB|V65.5|ICD9CM|Persn w feared complaint|Persn w feared complaint
C0851311|T033|PT|V65.5|ICD9CM|Person with feared complaint in whom no diagnosis was made|Person with feared complaint in whom no diagnosis was made
C0260825|T033|PT|V65.8|ICD9CM|Other reasons for seeking consultation|Other reasons for seeking consultation
C0260825|T033|AB|V65.8|ICD9CM|Reason for consult NEC|Reason for consult NEC
C0041880|T033|AB|V65.9|ICD9CM|Reason for consult NOS|Reason for consult NOS
C0041880|T033|PT|V65.9|ICD9CM|Unspecified reason for consultation|Unspecified reason for consultation
C0375891|T033|HT|V66|ICD9CM|Convalescence and palliative care|Convalescence and palliative care
C0260826|T033|PT|V66.0|ICD9CM|Convalescence following surgery|Convalescence following surgery
C0260826|T033|AB|V66.0|ICD9CM|Surgical convalescence|Surgical convalescence
C0260827|T033|PT|V66.1|ICD9CM|Convalescence following radiotherapy|Convalescence following radiotherapy
C0260827|T033|AB|V66.1|ICD9CM|Radiotherapy convalescen|Radiotherapy convalescen
C0260828|T033|AB|V66.2|ICD9CM|Chemotherapy convalescen|Chemotherapy convalescen
C0260828|T033|PT|V66.2|ICD9CM|Convalescence following chemotherapy|Convalescence following chemotherapy
C0481522|T033|PT|V66.3|ICD9CM|Convalescence following psychotherapy and other treatment for mental disorder|Convalescence following psychotherapy and other treatment for mental disorder
C0481522|T033|AB|V66.3|ICD9CM|Mental dis convalescence|Mental dis convalescence
C0260830|T033|PT|V66.4|ICD9CM|Convalescence following treatment of fracture|Convalescence following treatment of fracture
C0260830|T033|AB|V66.4|ICD9CM|Fracture treatmnt conval|Fracture treatmnt conval
C0009941|T033|PT|V66.5|ICD9CM|Convalescence following other treatment|Convalescence following other treatment
C0009941|T033|AB|V66.5|ICD9CM|Convalescence NEC|Convalescence NEC
C0375892|T033|PT|V66.7|ICD9CM|Encounter for palliative care|Encounter for palliative care
C0375892|T033|AB|V66.7|ICD9CM|Encountr palliative care|Encountr palliative care
C0677614|T033|AB|V66.9|ICD9CM|Convalescence NOS|Convalescence NOS
C0677614|T033|PT|V66.9|ICD9CM|Unspecified convalescence|Unspecified convalescence
C0260832|T033|HT|V67|ICD9CM|Follow-up examination|Follow-up examination
C0260833|T033|HT|V67.0|ICD9CM|Follow-up examination following surgery|Follow-up examination following surgery
C0878734|T033|PT|V67.00|ICD9CM|Follow-up examination, following surgery, unspecified|Follow-up examination, following surgery, unspecified
C0878734|T033|AB|V67.00|ICD9CM|Follow-up surgery NOS|Follow-up surgery NOS
C0878735|T033|AB|V67.01|ICD9CM|Follow-up vag pap smear|Follow-up vag pap smear
C0878735|T033|PT|V67.01|ICD9CM|Following surgery, follow-up vaginal pap smear|Following surgery, follow-up vaginal pap smear
C0878736|T033|PT|V67.09|ICD9CM|Follow-up examination, following other surgery|Follow-up examination, following other surgery
C0878736|T033|AB|V67.09|ICD9CM|Follow-up surgery NEC|Follow-up surgery NEC
C0260834|T033|PT|V67.1|ICD9CM|Follow-up examination, following radiotherapy|Follow-up examination, following radiotherapy
C0260834|T033|AB|V67.1|ICD9CM|Radiotherapy follow-up|Radiotherapy follow-up
C1261324|T033|AB|V67.2|ICD9CM|Chemotherapy follow-up|Chemotherapy follow-up
C1261324|T033|PT|V67.2|ICD9CM|Follow-up examination, following chemotherapy|Follow-up examination, following chemotherapy
C0260836|T033|PT|V67.3|ICD9CM|Follow-up examination, following psychotherapy and other treatment for mental disorder|Follow-up examination, following psychotherapy and other treatment for mental disorder
C0260836|T033|AB|V67.3|ICD9CM|Psychiatric follow-up|Psychiatric follow-up
C0481525|T033|PT|V67.4|ICD9CM|Follow-up examination, following treatment of healed fracture|Follow-up examination, following treatment of healed fracture
C0481525|T033|AB|V67.4|ICD9CM|FU exam treatd healed fx|FU exam treatd healed fx
C0260838|T033|HT|V67.5|ICD9CM|Follow-up examination following other treatment|Follow-up examination following other treatment
C0302433|T033|AB|V67.51|ICD9CM|High-risk rx NEC exam|High-risk rx NEC exam
C0260840|T033|AB|V67.59|ICD9CM|Follow-up exam NEC|Follow-up exam NEC
C0260840|T033|PT|V67.59|ICD9CM|Other follow-up examination|Other follow-up examination
C0260841|T033|AB|V67.6|ICD9CM|Comb treatment follow-up|Comb treatment follow-up
C0260841|T033|PT|V67.6|ICD9CM|Follow-up examination, following combined treatment|Follow-up examination, following combined treatment
C0260832|T033|AB|V67.9|ICD9CM|Follow-up exam NOS|Follow-up exam NOS
C0260832|T033|PT|V67.9|ICD9CM|Unspecified follow-up examination|Unspecified follow-up examination
C0260843|T033|HT|V68|ICD9CM|Encounters for administrative purposes|Encounters for administrative purposes
C0260844|T033|HT|V68.0|ICD9CM|Issue of medical certificates|Issue of medical certificates
C1955613|T033|AB|V68.01|ICD9CM|Disability examination|Disability examination
C1955613|T033|PT|V68.01|ICD9CM|Disability examination|Disability examination
C2910517|T033|AB|V68.09|ICD9CM|Issue of med certif NEC|Issue of med certif NEC
C2910517|T033|PT|V68.09|ICD9CM|Other issue of medical certificates|Other issue of medical certificates
C0260845|T033|PT|V68.1|ICD9CM|Issue of repeat prescriptions|Issue of repeat prescriptions
C0260845|T033|AB|V68.1|ICD9CM|Issue repeat prescript|Issue repeat prescript
C0260846|T033|AB|V68.2|ICD9CM|Request expert evidence|Request expert evidence
C0260846|T033|PT|V68.2|ICD9CM|Request for expert evidence|Request for expert evidence
C0260847|T033|HT|V68.8|ICD9CM|Encounters for other specified administrative purpose|Encounters for other specified administrative purpose
C0260848|T033|PT|V68.81|ICD9CM|Referral of patient without examination or treatment|Referral of patient without examination or treatment
C0260848|T033|AB|V68.81|ICD9CM|Referral-no exam/treat|Referral-no exam/treat
C0260847|T033|AB|V68.89|ICD9CM|Administrtve encount NEC|Administrtve encount NEC
C0260847|T033|PT|V68.89|ICD9CM|Encounters for other specified administrative purpose|Encounters for other specified administrative purpose
C0260849|T033|AB|V68.9|ICD9CM|Administrtve encount NOS|Administrtve encount NOS
C0260849|T033|PT|V68.9|ICD9CM|Encounters for unspecified administrative purpose|Encounters for unspecified administrative purpose
C0348087|T033|HT|V69|ICD9CM|Problems related to lifestyle|Problems related to lifestyle
C1306891|T033|PT|V69.0|ICD9CM|Lack of physical exercise|Lack of physical exercise
C1306891|T033|AB|V69.0|ICD9CM|Lack of physical exercse|Lack of physical exercse
C3537062|T033|PT|V69.1|ICD9CM|Inappropriate diet and eating habits|Inappropriate diet and eating habits
C3537062|T033|AB|V69.1|ICD9CM|Inapprt diet eat habits|Inapprt diet eat habits
C0348089|T033|PT|V69.2|ICD9CM|High-risk sexual behavior|High-risk sexual behavior
C0348089|T033|AB|V69.2|ICD9CM|High-risk sexual behavr|High-risk sexual behavr
C0348090|T033|AB|V69.3|ICD9CM|Gambling and betting|Gambling and betting
C0348090|T033|PT|V69.3|ICD9CM|Gambling and betting|Gambling and betting
C1455980|T033|AB|V69.4|ICD9CM|Lack of adequate sleep|Lack of adequate sleep
C1455980|T033|PT|V69.4|ICD9CM|Lack of adequate sleep|Lack of adequate sleep
C4317290|T033|AB|V69.5|ICD9CM|Behav insomnia-childhood|Behav insomnia-childhood
C4317290|T033|PT|V69.5|ICD9CM|Behavioral insomnia of childhood|Behavioral insomnia of childhood
C0348774|T033|AB|V69.8|ICD9CM|Oth prblms rltd lfstyle|Oth prblms rltd lfstyle
C0348774|T033|PT|V69.8|ICD9CM|Other problems related to lifestyle|Other problems related to lifestyle
C0348775|T033|AB|V69.9|ICD9CM|Prblm rltd lfstyle NOS|Prblm rltd lfstyle NOS
C0348775|T033|PT|V69.9|ICD9CM|Unspecified problem related to lifestyle|Unspecified problem related to lifestyle
C0260860|T033|HT|V70|ICD9CM|General medical examination|General medical examination
C0260851|T033|PT|V70.0|ICD9CM|Routine general medical examination at a health care facility|Routine general medical examination at a health care facility
C0260851|T033|AB|V70.0|ICD9CM|Routine medical exam|Routine medical exam
C0260852|T033|PT|V70.1|ICD9CM|General psychiatric examination, requested by the authority|General psychiatric examination, requested by the authority
C0260852|T033|AB|V70.1|ICD9CM|Psych exam-authority req|Psych exam-authority req
C0302434|T033|AB|V70.2|ICD9CM|Gen psychiatric exam NEC|Gen psychiatric exam NEC
C0302434|T033|PT|V70.2|ICD9CM|General psychiatric examination, other and unspecified|General psychiatric examination, other and unspecified
C0481845|T033|AB|V70.3|ICD9CM|Med exam NEC-admin purp|Med exam NEC-admin purp
C0481845|T033|PT|V70.3|ICD9CM|Other general medical examination for administrative purposes|Other general medical examination for administrative purposes
C0260855|T033|AB|V70.4|ICD9CM|Exam-medicolegal reasons|Exam-medicolegal reasons
C0260855|T033|PT|V70.4|ICD9CM|Examination for medicolegal reasons|Examination for medicolegal reasons
C0260857|T033|AB|V70.6|ICD9CM|Health exam-pop survey|Health exam-pop survey
C0260857|T033|PT|V70.6|ICD9CM|Health examination in population surveys|Health examination in population surveys
C0260859|T033|AB|V70.8|ICD9CM|General medical exam NEC|General medical exam NEC
C0260859|T033|PT|V70.8|ICD9CM|Other specified general medical examinations|Other specified general medical examinations
C0260860|T033|AB|V70.9|ICD9CM|General medical exam NOS|General medical exam NOS
C0260860|T033|PT|V70.9|ICD9CM|Unspecified general medical examination|Unspecified general medical examination
C0375893|T033|HT|V71|ICD9CM|Observation and evaluation for suspected conditions not found|Observation and evaluation for suspected conditions not found
C0260862|T033|HT|V71.0|ICD9CM|Observation for suspected mental condition|Observation for suspected mental condition
C0260863|T033|PT|V71.01|ICD9CM|Observation for adult antisocial behavior|Observation for adult antisocial behavior
C0260863|T033|AB|V71.01|ICD9CM|Obsv-adult antisoc behav|Obsv-adult antisoc behav
C0260864|T033|PT|V71.02|ICD9CM|Observation for childhood or adolescent antisocial behavior|Observation for childhood or adolescent antisocial behavior
C0260864|T033|AB|V71.02|ICD9CM|Obsv-adolesc antisoc beh|Obsv-adolesc antisoc beh
C0260865|T033|AB|V71.09|ICD9CM|Observ-mental cond NEC|Observ-mental cond NEC
C0260865|T033|PT|V71.09|ICD9CM|Observation for other suspected mental condition|Observation for other suspected mental condition
C0260866|T033|PT|V71.1|ICD9CM|Observation for suspected malignant neoplasm|Observation for suspected malignant neoplasm
C0260866|T033|AB|V71.1|ICD9CM|Obsv-suspct mal neoplasm|Obsv-suspct mal neoplasm
C0260867|T033|AB|V71.2|ICD9CM|Observ-suspect TB|Observ-suspect TB
C0260867|T033|PT|V71.2|ICD9CM|Observation for suspected tuberculosis|Observation for suspected tuberculosis
C0260868|T033|AB|V71.3|ICD9CM|Observ-work accident|Observ-work accident
C0260868|T033|PT|V71.3|ICD9CM|Observation following accident at work|Observation following accident at work
C0260869|T033|AB|V71.4|ICD9CM|Observ-accident NEC|Observ-accident NEC
C0260869|T033|PT|V71.4|ICD9CM|Observation following other accident|Observation following other accident
C0260870|T033|AB|V71.5|ICD9CM|Observ following rape|Observ following rape
C0260870|T033|PT|V71.5|ICD9CM|Observation following alleged rape or seduction|Observation following alleged rape or seduction
C0260871|T033|AB|V71.6|ICD9CM|Observ-inflicted inj NEC|Observ-inflicted inj NEC
C0260871|T033|PT|V71.6|ICD9CM|Observation following other inflicted injury|Observation following other inflicted injury
C0260872|T033|AB|V71.7|ICD9CM|Obs-susp cardiovasc dis|Obs-susp cardiovasc dis
C0260872|T033|PT|V71.7|ICD9CM|Observation for suspected cardiovascular disease|Observation for suspected cardiovascular disease
C0481850|T033|HT|V71.8|ICD9CM|Observation and evaluation for other specified suspected conditions|Observation and evaluation for other specified suspected conditions
C1135309|T033|AB|V71.82|ICD9CM|Obs/eval sus exp anthrax|Obs/eval sus exp anthrax
C1135309|T033|PT|V71.82|ICD9CM|Observation and evaluation for suspected exposure to anthrax|Observation and evaluation for suspected exposure to anthrax
C1135310|T033|AB|V71.83|ICD9CM|Obs/eval exp biol NEC|Obs/eval exp biol NEC
C1135310|T033|PT|V71.83|ICD9CM|Observation and evaluation for suspected exposure to other biological agent|Observation and evaluation for suspected exposure to other biological agent
C0481850|T033|AB|V71.89|ICD9CM|Observ-suspect cond NEC|Observ-suspect cond NEC
C0481850|T033|PT|V71.89|ICD9CM|Observation and evaluation for other specified suspected conditions|Observation and evaluation for other specified suspected conditions
C0490065|T033|AB|V71.9|ICD9CM|Observ-suspect cond NOS|Observ-suspect cond NOS
C0490065|T033|PT|V71.9|ICD9CM|Observation for unspecified suspected condition|Observation for unspecified suspected condition
C0260875|T033|HT|V72|ICD9CM|Special investigations and examinations|Special investigations and examinations
C1961134|T033|PT|V72.0|ICD9CM|Examination of eyes and vision|Examination of eyes and vision
C1961134|T033|AB|V72.0|ICD9CM|Eye & vision examination|Eye & vision examination
C0015222|T033|HT|V72.1|ICD9CM|Examination of ears and hearing|Examination of ears and hearing
C1719698|T033|PT|V72.11|ICD9CM|Encounter for hearing examination following failed hearing screening|Encounter for hearing examination following failed hearing screening
C1719698|T033|AB|V72.11|ICD9CM|Hearing exam-fail screen|Hearing exam-fail screen
C1955615|T033|PT|V72.12|ICD9CM|Encounter for hearing conservation and treatment|Encounter for hearing conservation and treatment
C1955615|T033|AB|V72.12|ICD9CM|Hearing conservatn/trtmt|Hearing conservatn/trtmt
C0490066|T033|AB|V72.2|ICD9CM|Dental examination|Dental examination
C0490066|T033|PT|V72.2|ICD9CM|Dental examination|Dental examination
C1455986|T033|HT|V72.3|ICD9CM|Special investigations and examinations - Gynecological examination|Special investigations and examinations - Gynecological examination
C1455982|T033|AB|V72.31|ICD9CM|Routine gyn examination|Routine gyn examination
C1455982|T033|PT|V72.31|ICD9CM|Routine gynecological examination|Routine gynecological examination
C1455985|T033|AB|V72.32|ICD9CM|Pap smear confirmation|Pap smear confirmation
C0260876|T033|PT|V72.40|ICD9CM|Pregnancy examination or test, pregnancy unconfirmed|Pregnancy examination or test, pregnancy unconfirmed
C0260876|T033|AB|V72.40|ICD9CM|Pregnancy test unconfirm|Pregnancy test unconfirm
C1455988|T033|PT|V72.41|ICD9CM|Pregnancy examination or test, negative result|Pregnancy examination or test, negative result
C1455988|T033|AB|V72.41|ICD9CM|Pregnancy test negative|Pregnancy test negative
C0869291|T033|AB|V72.5|ICD9CM|Radiological exam NEC|Radiological exam NEC
C0869291|T033|PT|V72.5|ICD9CM|Radiological examination, not elsewhere classified|Radiological examination, not elsewhere classified
C0260877|T033|HT|V72.6|ICD9CM|Laboratory examination|Laboratory examination
C2712559|T033|AB|V72.60|ICD9CM|Laboratory exam NOS|Laboratory exam NOS
C2712559|T033|PT|V72.60|ICD9CM|Laboratory examination, unspecified|Laboratory examination, unspecified
C2712560|T033|AB|V72.61|ICD9CM|Antibody response exam|Antibody response exam
C2712560|T033|PT|V72.61|ICD9CM|Antibody response examination|Antibody response examination
C2712561|T033|PT|V72.62|ICD9CM|Laboratory examination ordered as part of a routine general medical examination|Laboratory examination ordered as part of a routine general medical examination
C2712561|T033|AB|V72.62|ICD9CM|Routine physicl lab exam|Routine physicl lab exam
C2712562|T033|PT|V72.63|ICD9CM|Pre-procedural laboratory examination|Pre-procedural laboratory examination
C2712562|T033|AB|V72.63|ICD9CM|Pre-procedure lab exam|Pre-procedure lab exam
C2712563|T033|AB|V72.69|ICD9CM|Laboratory exam NEC|Laboratory exam NEC
C2712563|T033|PT|V72.69|ICD9CM|Other laboratory examination|Other laboratory examination
C0362085|T033|PT|V72.7|ICD9CM|Diagnostic skin and sensitization tests|Diagnostic skin and sensitization tests
C0362085|T033|AB|V72.7|ICD9CM|Skin/sensitization tests|Skin/sensitization tests
C0260879|T033|HT|V72.8|ICD9CM|Other specified examinations|Other specified examinations
C0375894|T033|PT|V72.81|ICD9CM|Pre-operative cardiovascular examination|Pre-operative cardiovascular examination
C0375894|T033|AB|V72.81|ICD9CM|Preop cardiovsclr exam|Preop cardiovsclr exam
C0375895|T033|PT|V72.82|ICD9CM|Pre-operative respiratory examination|Pre-operative respiratory examination
C0375895|T033|AB|V72.82|ICD9CM|Preop respiratory exam|Preop respiratory exam
C0375896|T033|AB|V72.83|ICD9CM|Oth spcf preop exam|Oth spcf preop exam
C0375896|T033|PT|V72.83|ICD9CM|Other specified pre-operative examination|Other specified pre-operative examination
C0375897|T033|PT|V72.84|ICD9CM|Pre-operative examination, unspecified|Pre-operative examination, unspecified
C0375897|T033|AB|V72.84|ICD9CM|Preop exam unspcf|Preop exam unspcf
C0260879|T033|AB|V72.85|ICD9CM|Oth specified exam|Oth specified exam
C0260879|T033|PT|V72.85|ICD9CM|Other specified examination|Other specified examination
C1561709|T033|AB|V72.86|ICD9CM|Blood typing encounter|Blood typing encounter
C1561709|T033|PT|V72.86|ICD9CM|Encounter for blood typing|Encounter for blood typing
C0260880|T033|AB|V72.9|ICD9CM|Examination NOS|Examination NOS
C0260880|T033|PT|V72.9|ICD9CM|Unspecified examination|Unspecified examination
C0375898|T033|HT|V73|ICD9CM|Special screening examination for viral and chlamydial diseases|Special screening examination for viral and chlamydial diseases
C0260882|T033|PT|V73.0|ICD9CM|Screening examination for poliomyelitis|Screening examination for poliomyelitis
C0260882|T033|AB|V73.0|ICD9CM|Screening-poliomyelitis|Screening-poliomyelitis
C0260883|T033|PT|V73.1|ICD9CM|Screening examination for smallpox|Screening examination for smallpox
C0260883|T033|AB|V73.1|ICD9CM|Screening for smallpox|Screening for smallpox
C0260884|T033|PT|V73.2|ICD9CM|Screening examination for measles|Screening examination for measles
C0260884|T033|AB|V73.2|ICD9CM|Screening for measles|Screening for measles
C0419585|T033|PT|V73.3|ICD9CM|Screening examination for rubella|Screening examination for rubella
C0419585|T033|AB|V73.3|ICD9CM|Screening for rubella|Screening for rubella
C1313924|T033|PT|V73.4|ICD9CM|Screening examination for yellow fever|Screening examination for yellow fever
C1313924|T033|AB|V73.4|ICD9CM|Screening-yellow fever|Screening-yellow fever
C0260887|T033|PT|V73.5|ICD9CM|Screening examination for other arthropod-borne viral diseases|Screening examination for other arthropod-borne viral diseases
C0260887|T033|AB|V73.5|ICD9CM|Screening-arbovirus dis|Screening-arbovirus dis
C0455701|T033|PT|V73.6|ICD9CM|Screening examination for trachoma|Screening examination for trachoma
C0455701|T033|AB|V73.6|ICD9CM|Screening for trachoma|Screening for trachoma
C1955616|T033|HT|V73.8|ICD9CM|Screening examination for other specified viral and chlamydial diseases|Screening examination for other specified viral and chlamydial diseases
C1959639|T033|AB|V73.81|ICD9CM|Special screen exam HPV|Special screen exam HPV
C1959639|T033|PT|V73.81|ICD9CM|Special screening examination for Human papillomavirus (HPV)|Special screening examination for Human papillomavirus (HPV)
C0375899|T033|AB|V73.88|ICD9CM|Scrn oth spcf chlmyd dis|Scrn oth spcf chlmyd dis
C0375899|T033|PT|V73.88|ICD9CM|Special screening examination for other specified chlamydial diseases|Special screening examination for other specified chlamydial diseases
C0260889|T033|AB|V73.89|ICD9CM|Scrn oth spcf viral dis|Scrn oth spcf viral dis
C0260889|T033|PT|V73.89|ICD9CM|Special screening examination for other specified viral diseases|Special screening examination for other specified viral diseases
C0700433|T033|HT|V73.9|ICD9CM|Screening examination for unspecified viral disease|Screening examination for unspecified viral disease
C0375900|T033|AB|V73.98|ICD9CM|Scrn unspcf chlmyd dis|Scrn unspcf chlmyd dis
C0375900|T033|PT|V73.98|ICD9CM|Special screening examination for unspecified chlamydial disease|Special screening examination for unspecified chlamydial disease
C0700433|T033|AB|V73.99|ICD9CM|Scrn unspcf viral dis|Scrn unspcf viral dis
C0700433|T033|PT|V73.99|ICD9CM|Special screening examination for unspecified viral disease|Special screening examination for unspecified viral disease
C0260899|T033|HT|V74|ICD9CM|Special screening examination for bacterial and spirochetal diseases|Special screening examination for bacterial and spirochetal diseases
C0260892|T033|PT|V74.0|ICD9CM|Screening examination for cholera|Screening examination for cholera
C0260892|T033|AB|V74.0|ICD9CM|Screening for cholera|Screening for cholera
C2910575|T033|PT|V74.1|ICD9CM|Screening examination for pulmonary tuberculosis|Screening examination for pulmonary tuberculosis
C2910575|T033|AB|V74.1|ICD9CM|Screening-pulmonary TB|Screening-pulmonary TB
C0420007|T033|PT|V74.2|ICD9CM|Screening examination for leprosy (Hansen's disease)|Screening examination for leprosy (Hansen's disease)
C0420007|T033|AB|V74.2|ICD9CM|Screening for leprosy|Screening for leprosy
C0260894|T033|PT|V74.3|ICD9CM|Screening examination for diphtheria|Screening examination for diphtheria
C0260894|T033|AB|V74.3|ICD9CM|Screening for diphtheria|Screening for diphtheria
C0260895|T033|AB|V74.4|ICD9CM|Screen-bact conjunctivit|Screen-bact conjunctivit
C0260895|T033|PT|V74.4|ICD9CM|Screening examination for bacterial conjunctivitis|Screening examination for bacterial conjunctivitis
C1961127|T033|AB|V74.5|ICD9CM|Screen for veneral dis|Screen for veneral dis
C1961127|T033|PT|V74.5|ICD9CM|Screening examination for venereal disease|Screening examination for venereal disease
C0260897|T033|PT|V74.6|ICD9CM|Screening examination for yaws|Screening examination for yaws
C0260897|T033|AB|V74.6|ICD9CM|Screening for yaws|Screening for yaws
C0260898|T033|AB|V74.8|ICD9CM|Screen-bacterial dis NEC|Screen-bacterial dis NEC
C0260898|T033|PT|V74.8|ICD9CM|Screening examination for other specified bacterial and spirochetal diseases|Screening examination for other specified bacterial and spirochetal diseases
C0260899|T033|AB|V74.9|ICD9CM|Screen-bacterial dis NOS|Screen-bacterial dis NOS
C0260899|T033|PT|V74.9|ICD9CM|Screening examination for unspecified bacterial and spirochetal diseases|Screening examination for unspecified bacterial and spirochetal diseases
C0260900|T033|HT|V75|ICD9CM|Special screening examination for other infectious diseases|Special screening examination for other infectious diseases
C0260901|T033|AB|V75.0|ICD9CM|Screen-rickettsial dis|Screen-rickettsial dis
C0260901|T033|PT|V75.0|ICD9CM|Screening examination for rickettsial diseases|Screening examination for rickettsial diseases
C0260902|T033|PT|V75.1|ICD9CM|Screening examination for malaria|Screening examination for malaria
C0260902|T033|AB|V75.1|ICD9CM|Screening for malaria|Screening for malaria
C0420015|T033|AB|V75.2|ICD9CM|Screen for leishmaniasis|Screen for leishmaniasis
C0420015|T033|PT|V75.2|ICD9CM|Screening examination for leishmaniasis|Screening examination for leishmaniasis
C0481870|T033|AB|V75.3|ICD9CM|Screen-trypanosomiasis|Screen-trypanosomiasis
C0481870|T033|PT|V75.3|ICD9CM|Screening examination for trypanosomiasis|Screening examination for trypanosomiasis
C0260905|T033|AB|V75.4|ICD9CM|Screen-mycotic infect|Screen-mycotic infect
C0260905|T033|PT|V75.4|ICD9CM|Screening examination for mycotic infections|Screening examination for mycotic infections
C0260906|T033|AB|V75.5|ICD9CM|Screen-schistosomiasis|Screen-schistosomiasis
C0260906|T033|PT|V75.5|ICD9CM|Screening examination for schistosomiasis|Screening examination for schistosomiasis
C0260907|T033|AB|V75.6|ICD9CM|Screen for filariasis|Screen for filariasis
C0260907|T033|PT|V75.6|ICD9CM|Screening examination for filariasis|Screening examination for filariasis
C1399262|T033|AB|V75.7|ICD9CM|Screen for helminthiasis|Screen for helminthiasis
C1399262|T033|PT|V75.7|ICD9CM|Screening examination for intestinal helminthiasis|Screening examination for intestinal helminthiasis
C0260909|T033|AB|V75.8|ICD9CM|Screen-parasitic dis NEC|Screen-parasitic dis NEC
C0260909|T033|PT|V75.8|ICD9CM|Screening examination for other specified parasitic infections|Screening examination for other specified parasitic infections
C0260910|T033|AB|V75.9|ICD9CM|Screen for infec dis NOS|Screen for infec dis NOS
C0260910|T033|PT|V75.9|ICD9CM|Screening examination for unspecified infectious disease|Screening examination for unspecified infectious disease
C0260922|T033|HT|V76|ICD9CM|Special screening for malignant neoplasms|Special screening for malignant neoplasms
C0481873|T033|AB|V76.0|ICD9CM|Screen mal neop-resp org|Screen mal neop-resp org
C0481873|T033|PT|V76.0|ICD9CM|Special screening for malignant neoplasms of respiratory organs|Special screening for malignant neoplasms of respiratory organs
C2921311|T033|HT|V76.1|ICD9CM|Screening examination for malignant neoplasms of the breast|Screening examination for malignant neoplasms of the breast
C0490031|T033|PT|V76.10|ICD9CM|Breast screening, unspecified|Breast screening, unspecified
C0490031|T033|AB|V76.10|ICD9CM|Scrn mal neo breast NOS|Scrn mal neo breast NOS
C0490033|T033|PT|V76.12|ICD9CM|Other screening mammogram|Other screening mammogram
C0490033|T033|AB|V76.12|ICD9CM|Screen mammogram NEC|Screen mammogram NEC
C0490034|T033|PT|V76.19|ICD9CM|Other screening breast examination|Other screening breast examination
C0490034|T033|AB|V76.19|ICD9CM|Scrn mal neo breast NEC|Scrn mal neo breast NEC
C0260914|T033|AB|V76.2|ICD9CM|Screen mal neop-cervix|Screen mal neop-cervix
C0260914|T033|PT|V76.2|ICD9CM|Screening for malignant neoplasms of cervix|Screening for malignant neoplasms of cervix
C0260915|T033|AB|V76.3|ICD9CM|Screen mal neop-bladder|Screen mal neop-bladder
C0260915|T033|PT|V76.3|ICD9CM|Screening for malignant neoplasms of bladder|Screening for malignant neoplasms of bladder
C0877843|T033|HT|V76.4|ICD9CM|Screening for malignant neoplasms of other sites|Screening for malignant neoplasms of other sites
C0260917|T033|AB|V76.41|ICD9CM|Screen mal neop-rectum|Screen mal neop-rectum
C0260917|T033|PT|V76.41|ICD9CM|Screening for malignant neoplasms of rectum|Screening for malignant neoplasms of rectum
C0260918|T033|AB|V76.42|ICD9CM|Screen mal neop-oral cav|Screen mal neop-oral cav
C0260918|T033|PT|V76.42|ICD9CM|Screening for malignant neoplasms of oral cavity|Screening for malignant neoplasms of oral cavity
C0260919|T033|AB|V76.43|ICD9CM|Screen mal neop-skin|Screen mal neop-skin
C0260919|T033|PT|V76.43|ICD9CM|Screening for malignant neoplasms of skin|Screening for malignant neoplasms of skin
C0699916|T033|PT|V76.44|ICD9CM|Screening for malignant neoplasms of prostate|Screening for malignant neoplasms of prostate
C0699916|T033|AB|V76.44|ICD9CM|Scrn malig neop-prostate|Scrn malig neop-prostate
C2910598|T033|AB|V76.45|ICD9CM|Screen malig neop-testis|Screen malig neop-testis
C2910598|T033|PT|V76.45|ICD9CM|Screening for malignant neoplasms of testis|Screening for malignant neoplasms of testis
C0878739|T033|AB|V76.47|ICD9CM|Screen malig neop-vagina|Screen malig neop-vagina
C0878739|T033|PT|V76.47|ICD9CM|Special screening for malignant neoplasms of vagina|Special screening for malignant neoplasms of vagina
C0877843|T033|AB|V76.49|ICD9CM|Screen mal neop oth site|Screen mal neop oth site
C0877843|T033|PT|V76.49|ICD9CM|Special screening for malignant neoplasms of other sites|Special screening for malignant neoplasms of other sites
C0878740|T033|HT|V76.5|ICD9CM|Screening for malignant neoplasms of intestine|Screening for malignant neoplasms of intestine
C0878741|T033|AB|V76.50|ICD9CM|Scrn malig neo-intes NOS|Scrn malig neo-intes NOS
C0878741|T033|PT|V76.50|ICD9CM|Special screening for malignant neoplasms for intestine, unspecified|Special screening for malignant neoplasms for intestine, unspecified
C0878742|T033|AB|V76.51|ICD9CM|Screen malig neop-colon|Screen malig neop-colon
C0878742|T033|PT|V76.51|ICD9CM|Special screening for malignant neoplasms of colon|Special screening for malignant neoplasms of colon
C2910590|T033|AB|V76.52|ICD9CM|Scrn mal neo-small intes|Scrn mal neo-small intes
C2910590|T033|PT|V76.52|ICD9CM|Special screening for malignant neoplasms of small intestine|Special screening for malignant neoplasms of small intestine
C0877844|T033|HT|V76.8|ICD9CM|Screening for other malignant neoplasms|Screening for other malignant neoplasms
C2910603|T033|AB|V76.81|ICD9CM|Screen neop-nervous syst|Screen neop-nervous syst
C2910603|T033|PT|V76.81|ICD9CM|Special screening for malignant neoplasms of nervous system|Special screening for malignant neoplasms of nervous system
C0260922|T033|AB|V76.9|ICD9CM|Screen-neoplasm NOS|Screen-neoplasm NOS
C0260922|T033|PT|V76.9|ICD9CM|Special screening for unspecified malignant neoplasms|Special screening for unspecified malignant neoplasms
C0260923|T033|HT|V77|ICD9CM|Special screening for endocrine, nutritional, metabolic, and immunity disorders|Special screening for endocrine, nutritional, metabolic, and immunity disorders
C0260924|T033|AB|V77.0|ICD9CM|Screen-thyroid disorder|Screen-thyroid disorder
C0260924|T033|PT|V77.0|ICD9CM|Screening for thyroid disorders|Screening for thyroid disorders
C0260925|T033|AB|V77.1|ICD9CM|Screen-diabetes mellitus|Screen-diabetes mellitus
C0260925|T033|PT|V77.1|ICD9CM|Screening for diabetes mellitus|Screening for diabetes mellitus
C0260926|T033|AB|V77.2|ICD9CM|Screen for malnutrition|Screen for malnutrition
C0260926|T033|PT|V77.2|ICD9CM|Screening for malnutrition|Screening for malnutrition
C0260927|T033|AB|V77.3|ICD9CM|Screen-phenylketonuria|Screen-phenylketonuria
C0260927|T033|PT|V77.3|ICD9CM|Screening for phenylketonuria (PKU)|Screening for phenylketonuria (PKU)
C0260928|T033|AB|V77.4|ICD9CM|Screen for galactosemia|Screen for galactosemia
C0260928|T033|PT|V77.4|ICD9CM|Screening for galactosemia|Screening for galactosemia
C0260929|T033|AB|V77.5|ICD9CM|Screening for gout|Screening for gout
C0260929|T033|PT|V77.5|ICD9CM|Screening for gout|Screening for gout
C0260930|T033|AB|V77.6|ICD9CM|Screen-cystic fibrosis|Screen-cystic fibrosis
C0260930|T033|PT|V77.6|ICD9CM|Screening for cystic fibrosis|Screening for cystic fibrosis
C0260931|T033|AB|V77.7|ICD9CM|Screen-inborn err metab|Screen-inborn err metab
C0260931|T033|PT|V77.7|ICD9CM|Screening for other inborn errors of metabolism|Screening for other inborn errors of metabolism
C0260932|T033|AB|V77.8|ICD9CM|Screening for obesity|Screening for obesity
C0260932|T033|PT|V77.8|ICD9CM|Screening for obesity|Screening for obesity
C0877845|T033|HT|V77.9|ICD9CM|Screening for other and unspecified endocrine, nutritional, metabolic and immunity disorders|Screening for other and unspecified endocrine, nutritional, metabolic and immunity disorders
C2910614|T033|AB|V77.91|ICD9CM|Screen lipoid disorders|Screen lipoid disorders
C2910614|T033|PT|V77.91|ICD9CM|Screening for lipoid disorders|Screening for lipoid disorders
C0877845|T033|AB|V77.99|ICD9CM|Screen-endoc/nut/met NEC|Screen-endoc/nut/met NEC
C0877845|T033|PT|V77.99|ICD9CM|Screening for other and unspecified endocrine, nutritional, metabolic, and immunity disorders|Screening for other and unspecified endocrine, nutritional, metabolic, and immunity disorders
C0260934|T033|HT|V78|ICD9CM|Special screening for disorders of blood and blood-forming organs|Special screening for disorders of blood and blood-forming organs
C0260935|T033|AB|V78.0|ICD9CM|Screen-iron defic anemia|Screen-iron defic anemia
C0260935|T033|PT|V78.0|ICD9CM|Screening for iron deficiency anemia|Screening for iron deficiency anemia
C0260936|T033|AB|V78.1|ICD9CM|Screen-defic anemia NEC|Screen-defic anemia NEC
C0260936|T033|PT|V78.1|ICD9CM|Screening for other and unspecified deficiency anemia|Screening for other and unspecified deficiency anemia
C0260937|T033|AB|V78.2|ICD9CM|Screen-sickle cell dis|Screen-sickle cell dis
C0260937|T033|PT|V78.2|ICD9CM|Screening for sickle-cell disease or trait|Screening for sickle-cell disease or trait
C2586327|T033|PT|V78.3|ICD9CM|Screening for other hemoglobinopathies|Screening for other hemoglobinopathies
C2586327|T033|AB|V78.3|ICD9CM|Scrn-hemoglobinopath NEC|Scrn-hemoglobinopath NEC
C0260939|T033|AB|V78.8|ICD9CM|Screen-blood dis NEC|Screen-blood dis NEC
C0260939|T033|PT|V78.8|ICD9CM|Screening for other disorders of blood and blood-forming organs|Screening for other disorders of blood and blood-forming organs
C0260940|T033|AB|V78.9|ICD9CM|Screen-blood dis NOS|Screen-blood dis NOS
C0260940|T033|PT|V78.9|ICD9CM|Screening for unspecified disorder of blood and blood-forming organs|Screening for unspecified disorder of blood and blood-forming organs
C0260941|T033|HT|V79|ICD9CM|Special screening for mental disorders and developmental handicaps|Special screening for mental disorders and developmental handicaps
C0260942|T033|AB|V79.0|ICD9CM|Screening for depression|Screening for depression
C0260942|T033|PT|V79.0|ICD9CM|Screening for depression|Screening for depression
C0260943|T033|AB|V79.1|ICD9CM|Screening for alcoholism|Screening for alcoholism
C0260943|T033|PT|V79.1|ICD9CM|Screening for alcoholism|Screening for alcoholism
C0260944|T033|AB|V79.2|ICD9CM|Scrn intellect disabilty|Scrn intellect disabilty
C0260944|T033|PT|V79.2|ICD9CM|Special screening for intellectual disabilities|Special screening for intellectual disabilities
C0260945|T033|AB|V79.3|ICD9CM|Screen-development prob|Screen-development prob
C0260945|T033|PT|V79.3|ICD9CM|Screening for developmental handicaps in early childhood|Screening for developmental handicaps in early childhood
C0260946|T033|AB|V79.8|ICD9CM|Screen-mental dis NEC|Screen-mental dis NEC
C0260946|T033|PT|V79.8|ICD9CM|Screening for other specified mental disorders and developmental handicaps|Screening for other specified mental disorders and developmental handicaps
C0600027|T033|AB|V79.9|ICD9CM|Screen-mental dis NOS|Screen-mental dis NOS
C0600027|T033|PT|V79.9|ICD9CM|Screening for unspecified mental disorder and developmental handicap|Screening for unspecified mental disorder and developmental handicap
C0260948|T033|HT|V80|ICD9CM|Special screening for neurological, eye, and ear diseases|Special screening for neurological, eye, and ear diseases
C0260949|T033|HT|V80.0|ICD9CM|Screening for neurological conditions|Screening for neurological conditions
C2921402|T033|AB|V80.01|ICD9CM|Screen-traumtc brain inj|Screen-traumtc brain inj
C2921402|T033|PT|V80.01|ICD9CM|Special screening for traumatic brain injury|Special screening for traumatic brain injury
C2712564|T033|AB|V80.09|ICD9CM|Screen-neuro condition|Screen-neuro condition
C2712564|T033|PT|V80.09|ICD9CM|Special screening for other neurological conditions|Special screening for other neurological conditions
C0260950|T033|AB|V80.1|ICD9CM|Screening for glaucoma|Screening for glaucoma
C0260950|T033|PT|V80.1|ICD9CM|Screening for glaucoma|Screening for glaucoma
C0260951|T033|PT|V80.2|ICD9CM|Screening for other eye conditions|Screening for other eye conditions
C0260951|T033|AB|V80.2|ICD9CM|Screening-eye cond NEC|Screening-eye cond NEC
C0260952|T033|AB|V80.3|ICD9CM|Screening for ear dis|Screening for ear dis
C0260952|T033|PT|V80.3|ICD9CM|Screening for ear diseases|Screening for ear diseases
C0260953|T033|HT|V81|ICD9CM|Special screening for cardiovascular, respiratory, and genitourinary diseases|Special screening for cardiovascular, respiratory, and genitourinary diseases
C0260954|T033|PT|V81.0|ICD9CM|Screening for ischemic heart disease|Screening for ischemic heart disease
C0260954|T033|AB|V81.0|ICD9CM|Scrn-ischemic heart dis|Scrn-ischemic heart dis
C0260955|T033|AB|V81.1|ICD9CM|Screen for hypertension|Screen for hypertension
C0260955|T033|PT|V81.1|ICD9CM|Screening for hypertension|Screening for hypertension
C0260956|T033|AB|V81.2|ICD9CM|Screen-cardiovasc NEC|Screen-cardiovasc NEC
C0260956|T033|PT|V81.2|ICD9CM|Screening for other and unspecified cardiovascular conditions|Screening for other and unspecified cardiovascular conditions
C0260957|T033|AB|V81.3|ICD9CM|Screen-bronch/emphysema|Screen-bronch/emphysema
C0260957|T033|PT|V81.3|ICD9CM|Screening for chronic bronchitis and emphysema|Screening for chronic bronchitis and emphysema
C0260958|T033|AB|V81.4|ICD9CM|Screen-respir cond NEC|Screen-respir cond NEC
C0260958|T033|PT|V81.4|ICD9CM|Screening for other and unspecified respiratory conditions|Screening for other and unspecified respiratory conditions
C0260959|T033|AB|V81.5|ICD9CM|Screen for nephropathy|Screen for nephropathy
C0260959|T033|PT|V81.5|ICD9CM|Screening for nephropathy|Screening for nephropathy
C0260960|T033|AB|V81.6|ICD9CM|Screen for gu cond NEC|Screen for gu cond NEC
C0260960|T033|PT|V81.6|ICD9CM|Screening for other and unspecified genitourinary conditions|Screening for other and unspecified genitourinary conditions
C0260961|T033|HT|V82|ICD9CM|Special screening for other conditions|Special screening for other conditions
C0260962|T033|AB|V82.0|ICD9CM|Screen for skin cond|Screen for skin cond
C0260962|T033|PT|V82.0|ICD9CM|Screening for skin conditions|Screening for skin conditions
C0260963|T033|AB|V82.1|ICD9CM|Screen-rheumatoid arthr|Screen-rheumatoid arthr
C0260963|T033|PT|V82.1|ICD9CM|Screening for rheumatoid arthritis|Screening for rheumatoid arthritis
C0260964|T033|AB|V82.2|ICD9CM|Screen-rheumat dis NEC|Screen-rheumat dis NEC
C0260964|T033|PT|V82.2|ICD9CM|Screening for other rheumatic disorders|Screening for other rheumatic disorders
C0260965|T033|AB|V82.3|ICD9CM|Screen-cong hip dislocat|Screen-cong hip dislocat
C0260965|T033|PT|V82.3|ICD9CM|Screening for congenital dislocation of hip|Screening for congenital dislocation of hip
C0695272|T033|AB|V82.4|ICD9CM|Mat pstntl scr-chrm anom|Mat pstntl scr-chrm anom
C0695272|T033|PT|V82.4|ICD9CM|Maternal postnatal screening for chromosomal anomalies|Maternal postnatal screening for chromosomal anomalies
C0260967|T033|AB|V82.5|ICD9CM|Screen-contamination NEC|Screen-contamination NEC
C0260967|T033|PT|V82.5|ICD9CM|Screening for chemical poisoning and other contamination|Screening for chemical poisoning and other contamination
C0740225|T033|AB|V82.6|ICD9CM|Multiphasic screening|Multiphasic screening
C0740225|T033|PT|V82.6|ICD9CM|Multiphasic screening|Multiphasic screening
C0017394|T033|HT|V82.7|ICD9CM|Genetic screening|Genetic screening
C0017394|T033|AB|V82.79|ICD9CM|Genetic screening NEC|Genetic screening NEC
C0017394|T033|PT|V82.79|ICD9CM|Other genetic screening|Other genetic screening
C0036464|T033|HT|V82.8|ICD9CM|Screening for other specified conditions|Screening for other specified conditions
C2910630|T033|AB|V82.81|ICD9CM|Screen - osteoporosis|Screen - osteoporosis
C2910630|T033|PT|V82.81|ICD9CM|Special screening for osteoporosis|Special screening for osteoporosis
C0036464|T033|AB|V82.89|ICD9CM|Screen for condition NEC|Screen for condition NEC
C0036464|T033|PT|V82.89|ICD9CM|Special screening for other specified conditions|Special screening for other specified conditions
C0949156|T033|HT|V83|ICD9CM|Genetic carrier status|Genetic carrier status
C2919122|T033|HT|V83.0|ICD9CM|Hemophilia A carrier|Hemophilia A carrier
C2911654|T033|AB|V83.01|ICD9CM|Asympt hemoph a carrier|Asympt hemoph a carrier
C2911654|T033|PT|V83.01|ICD9CM|Asymptomatic hemophilia A carrier|Asymptomatic hemophilia A carrier
C2911655|T033|AB|V83.02|ICD9CM|Sympt hemophil a carrier|Sympt hemophil a carrier
C2911655|T033|PT|V83.02|ICD9CM|Symptomatic hemophilia A carrier|Symptomatic hemophilia A carrier
C1135312|T033|HT|V83.8|ICD9CM|Other genetic carrier status|Other genetic carrier status
C2711060|T033|AB|V83.81|ICD9CM|Cystic fibrosis gene car|Cystic fibrosis gene car
C2711060|T033|PT|V83.81|ICD9CM|Cystic fibrosis gene carrier|Cystic fibrosis gene carrier
C1135312|T033|AB|V83.89|ICD9CM|Genetic carrier stat NEC|Genetic carrier stat NEC
C1135312|T033|PT|V83.89|ICD9CM|Other genetic carrier status|Other genetic carrier status
C2919134|T033|HT|V84|ICD9CM|Genetic susceptibility to disease|Genetic susceptibility to disease
C1455995|T033|HT|V84.0|ICD9CM|Genetic susceptibility to malignant neoplasm|Genetic susceptibility to malignant neoplasm
C1455990|T033|AB|V84.01|ICD9CM|Genetc sus mal neo brest|Genetc sus mal neo brest
C1455990|T033|PT|V84.01|ICD9CM|Genetic susceptibility to malignant neoplasm of breast|Genetic susceptibility to malignant neoplasm of breast
C1455991|T033|AB|V84.02|ICD9CM|Genetc sus mal neo ovary|Genetc sus mal neo ovary
C1455991|T033|PT|V84.02|ICD9CM|Genetic susceptibility to malignant neoplasm of ovary|Genetic susceptibility to malignant neoplasm of ovary
C1455992|T033|AB|V84.03|ICD9CM|Genetc sus mal neo prost|Genetc sus mal neo prost
C1455992|T033|PT|V84.03|ICD9CM|Genetic susceptibility to malignant neoplasm of prostate|Genetic susceptibility to malignant neoplasm of prostate
C1455993|T033|AB|V84.04|ICD9CM|Genetc susc mal neo endo|Genetc susc mal neo endo
C1455993|T033|PT|V84.04|ICD9CM|Genetic susceptibility to malignant neoplasm of endometrium|Genetic susceptibility to malignant neoplasm of endometrium
C1455994|T033|AB|V84.09|ICD9CM|Genetic susc mal neo NEC|Genetic susc mal neo NEC
C1455994|T033|PT|V84.09|ICD9CM|Genetic susceptibility to other malignant neoplasm|Genetic susceptibility to other malignant neoplasm
C1455996|T033|HT|V84.8|ICD9CM|Genetic susceptibility to other disease|Genetic susceptibility to other disease
C1955618|T033|AB|V84.81|ICD9CM|Genetc sus mult endo neo|Genetc sus mult endo neo
C1955618|T033|PT|V84.81|ICD9CM|Genetic susceptibility to multiple endocrine neoplasia [MEN]|Genetic susceptibility to multiple endocrine neoplasia [MEN]
C1455996|T033|AB|V84.89|ICD9CM|Genetic suscept dis NEC|Genetic suscept dis NEC
C1455996|T033|PT|V84.89|ICD9CM|Genetic susceptibility to other disease|Genetic susceptibility to other disease
C2240399|T033|HT|V85|ICD9CM|Body mass index [BMI]|Body mass index [BMI]
C2240399|T033|HT|V85-V85.99|ICD9CM|BODY MASS INDEX|BODY MASS INDEX
C1561710|T033|AB|V85.0|ICD9CM|BMI less than 19,adult|BMI less than 19,adult
C1561710|T033|PT|V85.0|ICD9CM|Body Mass Index less than 19, adult|Body Mass Index less than 19, adult
C1561711|T033|AB|V85.1|ICD9CM|BMI between 19-24,adult|BMI between 19-24,adult
C1561711|T033|PT|V85.1|ICD9CM|Body Mass Index between 19-24, adult|Body Mass Index between 19-24, adult
C1561717|T033|HT|V85.2|ICD9CM|Body Mass Index between 25-29, adult|Body Mass Index between 25-29, adult
C2911045|T033|AB|V85.21|ICD9CM|BMI 25.0-25.9,adult|BMI 25.0-25.9,adult
C2911045|T033|PT|V85.21|ICD9CM|Body Mass Index 25.0-25.9, adult|Body Mass Index 25.0-25.9, adult
C2911046|T033|AB|V85.22|ICD9CM|BMI 26.0-26.9,adult|BMI 26.0-26.9,adult
C2911046|T033|PT|V85.22|ICD9CM|Body Mass Index 26.0-26.9, adult|Body Mass Index 26.0-26.9, adult
C2911047|T033|AB|V85.23|ICD9CM|BMI 27.0-27.9,adult|BMI 27.0-27.9,adult
C2911047|T033|PT|V85.23|ICD9CM|Body Mass Index 27.0-27.9, adult|Body Mass Index 27.0-27.9, adult
C2911048|T033|AB|V85.24|ICD9CM|BMI 28.0-28.9,adult|BMI 28.0-28.9,adult
C2911048|T033|PT|V85.24|ICD9CM|Body Mass Index 28.0-28.9, adult|Body Mass Index 28.0-28.9, adult
C2911049|T033|AB|V85.25|ICD9CM|BMI 29.0-29.9,adult|BMI 29.0-29.9,adult
C2911049|T033|PT|V85.25|ICD9CM|Body Mass Index 29.0-29.9, adult|Body Mass Index 29.0-29.9, adult
C1561728|T033|HT|V85.3|ICD9CM|Body Mass Index between 30-39, adult|Body Mass Index between 30-39, adult
C2911051|T033|AB|V85.30|ICD9CM|BMI 30.0-30.9,adult|BMI 30.0-30.9,adult
C2911051|T033|PT|V85.30|ICD9CM|Body Mass Index 30.0-30.9, adult|Body Mass Index 30.0-30.9, adult
C2911052|T033|AB|V85.31|ICD9CM|BMI 31.0-31.9,adult|BMI 31.0-31.9,adult
C2911052|T033|PT|V85.31|ICD9CM|Body Mass Index 31.0-31.9, adult|Body Mass Index 31.0-31.9, adult
C2911053|T033|AB|V85.32|ICD9CM|BMI 32.0-32.9,adult|BMI 32.0-32.9,adult
C2911053|T033|PT|V85.32|ICD9CM|Body Mass Index 32.0-32.9, adult|Body Mass Index 32.0-32.9, adult
C2911054|T033|AB|V85.33|ICD9CM|BMI 33.0-33.9,adult|BMI 33.0-33.9,adult
C2911054|T033|PT|V85.33|ICD9CM|Body Mass Index 33.0-33.9, adult|Body Mass Index 33.0-33.9, adult
C2911055|T033|AB|V85.34|ICD9CM|BMI 34.0-34.9,adult|BMI 34.0-34.9,adult
C2911055|T033|PT|V85.34|ICD9CM|Body Mass Index 34.0-34.9, adult|Body Mass Index 34.0-34.9, adult
C2911056|T033|AB|V85.35|ICD9CM|BMI 35.0-35.9,adult|BMI 35.0-35.9,adult
C2911056|T033|PT|V85.35|ICD9CM|Body Mass Index 35.0-35.9, adult|Body Mass Index 35.0-35.9, adult
C2911057|T033|AB|V85.36|ICD9CM|BMI 36.0-36.9,adult|BMI 36.0-36.9,adult
C2911057|T033|PT|V85.36|ICD9CM|Body Mass Index 36.0-36.9, adult|Body Mass Index 36.0-36.9, adult
C2911058|T033|AB|V85.37|ICD9CM|BMI 37.0-37.9,adult|BMI 37.0-37.9,adult
C2911058|T033|PT|V85.37|ICD9CM|Body Mass Index 37.0-37.9, adult|Body Mass Index 37.0-37.9, adult
C2911059|T033|AB|V85.38|ICD9CM|BMI 38.0-38.9,adult|BMI 38.0-38.9,adult
C2911059|T033|PT|V85.38|ICD9CM|Body Mass Index 38.0-38.9, adult|Body Mass Index 38.0-38.9, adult
C2911060|T033|AB|V85.39|ICD9CM|BMI 39.0-39.9,adult|BMI 39.0-39.9,adult
C2911060|T033|PT|V85.39|ICD9CM|Body Mass Index 39.0-39.9, adult|Body Mass Index 39.0-39.9, adult
C1561729|T033|HT|V85.4|ICD9CM|Body Mass Index 40 and over, adult|Body Mass Index 40 and over, adult
C2921312|T033|AB|V85.41|ICD9CM|BMI 40.0-44.9, adult|BMI 40.0-44.9, adult
C2921312|T033|PT|V85.41|ICD9CM|Body Mass Index 40.0-44.9, adult|Body Mass Index 40.0-44.9, adult
C2921313|T033|AB|V85.42|ICD9CM|BMI 45.0-49.9, adult|BMI 45.0-49.9, adult
C2921313|T033|PT|V85.42|ICD9CM|Body Mass Index 45.0-49.9, adult|Body Mass Index 45.0-49.9, adult
C2921314|T033|AB|V85.43|ICD9CM|BMI 50.0-59.9, adult|BMI 50.0-59.9, adult
C2921314|T033|PT|V85.43|ICD9CM|Body Mass Index 50.0-59.9, adult|Body Mass Index 50.0-59.9, adult
C2921315|T033|AB|V85.44|ICD9CM|BMI 60.0-69.9, adult|BMI 60.0-69.9, adult
C2921315|T033|PT|V85.44|ICD9CM|Body Mass Index 60.0-69.9, adult|Body Mass Index 60.0-69.9, adult
C2921316|T033|AB|V85.45|ICD9CM|BMI 70 and over, adult|BMI 70 and over, adult
C2921316|T033|PT|V85.45|ICD9CM|Body Mass Index 70 and over, adult|Body Mass Index 70 and over, adult
C2911062|T033|HT|V85.5|ICD9CM|Body Mass Index, pediatric|Body Mass Index, pediatric
C2911063|T033|AB|V85.51|ICD9CM|BMI,pediatric <5%|BMI,pediatric <5%
C2911063|T033|PT|V85.51|ICD9CM|Body Mass Index, pediatric, less than 5th percentile for age|Body Mass Index, pediatric, less than 5th percentile for age
C2911064|T033|AB|V85.52|ICD9CM|BMI,pediatric 5% - <85%|BMI,pediatric 5% - <85%
C2911064|T033|PT|V85.52|ICD9CM|Body Mass Index, pediatric, 5th percentile to less than 85th percentile for age|Body Mass Index, pediatric, 5th percentile to less than 85th percentile for age
C2911065|T033|AB|V85.53|ICD9CM|BMI,pediatric 85% - <95%|BMI,pediatric 85% - <95%
C2911065|T033|PT|V85.53|ICD9CM|Body Mass Index, pediatric, 85th percentile to less than 95th percentile for age|Body Mass Index, pediatric, 85th percentile to less than 95th percentile for age
C2911066|T033|AB|V85.54|ICD9CM|BMI,pediatric >= 95%|BMI,pediatric >= 95%
C2911066|T033|PT|V85.54|ICD9CM|Body Mass Index, pediatric, greater than or equal to 95th percentile for age|Body Mass Index, pediatric, greater than or equal to 95th percentile for age
C2919114|T033|HT|V86|ICD9CM|Estrogen receptor status|Estrogen receptor status
C2919114|T033|HT|V86-V86.99|ICD9CM|ESTROGEN RECEPTOR STATUS|ESTROGEN RECEPTOR STATUS
C1719706|T033|AB|V86.0|ICD9CM|Estrogen recep pstv stat|Estrogen recep pstv stat
C1719706|T033|PT|V86.0|ICD9CM|Estrogen receptor positive status [ER+]|Estrogen receptor positive status [ER+]
C1719707|T033|AB|V86.1|ICD9CM|Estrogen recep neg stat|Estrogen recep neg stat
C1719707|T033|PT|V86.1|ICD9CM|Estrogen receptor negative status [ER-]|Estrogen receptor negative status [ER-]
C2349917|T047|HT|V87|ICD9CM|Other specified personal exposures and history presenting hazards to health|Other specified personal exposures and history presenting hazards to health
C2349917|T047|HT|V87-V87.99|ICD9CM|OTHER SPECIFIED PERSONAL EXPOSURES AND HISTORY PRESENTING HAZARDS TO HEALTH|OTHER SPECIFIED PERSONAL EXPOSURES AND HISTORY PRESENTING HAZARDS TO HEALTH
C2349903|T033|HT|V87.0|ICD9CM|Contact with and (suspected) exposure to hazardous metals|Contact with and (suspected) exposure to hazardous metals
C2349899|T033|PT|V87.01|ICD9CM|Contact with and (suspected) exposure to arsenic|Contact with and (suspected) exposure to arsenic
C2349899|T033|AB|V87.01|ICD9CM|Contact/exposure arsenic|Contact/exposure arsenic
C3161155|T033|AB|V87.02|ICD9CM|Cont/susp expose uranium|Cont/susp expose uranium
C3161155|T033|PT|V87.02|ICD9CM|Contact with and (suspected) exposure to uranium|Contact with and (suspected) exposure to uranium
C2349900|T033|AB|V87.09|ICD9CM|Cntct/exp hazrd metl NEC|Cntct/exp hazrd metl NEC
C2349900|T033|PT|V87.09|ICD9CM|Contact with and (suspected) exposure to other hazardous metals|Contact with and (suspected) exposure to other hazardous metals
C2349909|T033|HT|V87.1|ICD9CM|Contact with and (suspected) exposure to hazardous aromatic compounds|Contact with and (suspected) exposure to hazardous aromatic compounds
C2349904|T033|AB|V87.11|ICD9CM|Cntct/exp aromatc amines|Cntct/exp aromatc amines
C2349904|T033|PT|V87.11|ICD9CM|Contact with and (suspected) exposure to aromatic amines|Contact with and (suspected) exposure to aromatic amines
C2349905|T033|PT|V87.12|ICD9CM|Contact with and (suspected) exposure to benzene|Contact with and (suspected) exposure to benzene
C2349905|T033|AB|V87.12|ICD9CM|Contact/exposure benzene|Contact/exposure benzene
C2349906|T033|AB|V87.19|ICD9CM|Cont/exp haz aromat NEC|Cont/exp haz aromat NEC
C2349906|T033|PT|V87.19|ICD9CM|Contact with and (suspected) exposure to other hazardous aromatic compounds|Contact with and (suspected) exposure to other hazardous aromatic compounds
C2349910|T033|AB|V87.2|ICD9CM|Cont/exp hazard chem NEC|Cont/exp hazard chem NEC
C2349910|T033|PT|V87.2|ICD9CM|Contact with and (suspected) exposure to other potentially hazardous chemicals|Contact with and (suspected) exposure to other potentially hazardous chemicals
C2349912|T033|HT|V87.3|ICD9CM|Contact with and (suspected ) exposure to other potentially hazardous substances|Contact with and (suspected ) exposure to other potentially hazardous substances
C2362603|T033|PT|V87.31|ICD9CM|Contact with and (suspected) exposure to mold|Contact with and (suspected) exposure to mold
C2362603|T033|AB|V87.31|ICD9CM|Contact/exposure mold|Contact/exposure mold
C2712565|T033|PT|V87.32|ICD9CM|Contact with and (suspected) exposure to algae bloom|Contact with and (suspected) exposure to algae bloom
C2712565|T033|AB|V87.32|ICD9CM|Contact/exp algae bloom|Contact/exp algae bloom
C2349912|T033|AB|V87.39|ICD9CM|Cont/exp hazard sub NEC|Cont/exp hazard sub NEC
C2349912|T033|PT|V87.39|ICD9CM|Contact with and (suspected) exposure to other potentially hazardous substances|Contact with and (suspected) exposure to other potentially hazardous substances
C2349916|T033|HT|V87.4|ICD9CM|Personal history of drug therapy|Personal history of drug therapy
C2349913|T033|AB|V87.41|ICD9CM|Hx antineoplastic chemo|Hx antineoplastic chemo
C2349913|T033|PT|V87.41|ICD9CM|Personal history of antineoplastic chemotherapy|Personal history of antineoplastic chemotherapy
C2349914|T033|AB|V87.42|ICD9CM|Hx monoclonal drug thrpy|Hx monoclonal drug thrpy
C2349914|T033|PT|V87.42|ICD9CM|Personal history of monoclonal drug therapy|Personal history of monoclonal drug therapy
C2712566|T033|AB|V87.43|ICD9CM|Hx estrogen therapy|Hx estrogen therapy
C2712566|T033|PT|V87.43|ICD9CM|Personal history of estrogen therapy|Personal history of estrogen therapy
C2712567|T033|AB|V87.44|ICD9CM|Hx inhaled steroid thrpy|Hx inhaled steroid thrpy
C2712567|T033|PT|V87.44|ICD9CM|Personal history of inhaled steroid therapy|Personal history of inhaled steroid therapy
C2712644|T033|AB|V87.45|ICD9CM|Hx systemc steroid thrpy|Hx systemc steroid thrpy
C2712644|T033|PT|V87.45|ICD9CM|Personal history of systemic steroid therapy|Personal history of systemic steroid therapy
C2911483|T033|AB|V87.46|ICD9CM|Hx immunosuppres thrpy|Hx immunosuppres thrpy
C2911483|T033|PT|V87.46|ICD9CM|Personal history of immunosuppressive therapy|Personal history of immunosuppressive therapy
C2349915|T033|AB|V87.49|ICD9CM|Hx drug therapy NEC|Hx drug therapy NEC
C2349915|T033|PT|V87.49|ICD9CM|Personal history of other drug therapy|Personal history of other drug therapy
C2349918|T033|HT|V88|ICD9CM|Acquired absence of other organs and tissue|Acquired absence of other organs and tissue
C2349918|T033|HT|V88-V88.99|ICD9CM|ACQUIRED ABSENCE OF OTHER ORGANS AND TISSUE|ACQUIRED ABSENCE OF OTHER ORGANS AND TISSUE
C2349925|T020|HT|V88.0|ICD9CM|Acquired absence of cervix and uterus|Acquired absence of cervix and uterus
C2349919|T033|AB|V88.01|ICD9CM|Acq absnce cervix/uterus|Acq absnce cervix/uterus
C2349919|T033|PT|V88.01|ICD9CM|Acquired absence of both cervix and uterus|Acquired absence of both cervix and uterus
C2349922|T033|AB|V88.02|ICD9CM|Acq ab ut remn cerv stmp|Acq ab ut remn cerv stmp
C2349922|T033|PT|V88.02|ICD9CM|Acquired absence of uterus with remaining cervical stump|Acquired absence of uterus with remaining cervical stump
C2349924|T033|AB|V88.03|ICD9CM|Acq absnc cerv/remain ut|Acq absnc cerv/remain ut
C2349924|T033|PT|V88.03|ICD9CM|Acquired absence of cervix with remaining uterus|Acquired absence of cervix with remaining uterus
C1386808|T020|HT|V88.1|ICD9CM|Acquired absence of pancreas|Acquired absence of pancreas
C2921317|T033|AB|V88.11|ICD9CM|Acq total absnc pancreas|Acq total absnc pancreas
C2921317|T033|PT|V88.11|ICD9CM|Acquired total absence of pancreas|Acquired total absence of pancreas
C2921318|T033|AB|V88.12|ICD9CM|Acq part absnce pancreas|Acq part absnce pancreas
C2921318|T033|PT|V88.12|ICD9CM|Acquired partial absence of pancreas|Acquired partial absence of pancreas
C3161260|T020|HT|V88.2|ICD9CM|Acquired absence of joint|Acquired absence of joint
C3161156|T020|AB|V88.21|ICD9CM|Acq absence of hip joint|Acq absence of hip joint
C3161156|T020|PT|V88.21|ICD9CM|Acquired absence of hip joint|Acquired absence of hip joint
C3161157|T020|AB|V88.22|ICD9CM|Acq absence knee joint|Acq absence knee joint
C3161157|T020|PT|V88.22|ICD9CM|Acquired absence of knee joint|Acquired absence of knee joint
C3161158|T020|AB|V88.29|ICD9CM|Acq absence of oth joint|Acq absence of oth joint
C3161158|T020|PT|V88.29|ICD9CM|Acquired absence of other joint|Acquired absence of other joint
C2349935|T047|HT|V89|ICD9CM|Other suspected conditions not found|Other suspected conditions not found
C2349935|T047|HT|V89-V89.99|ICD9CM|OTHER SUSPECTED CONDITIONS NOT FOUND|OTHER SUSPECTED CONDITIONS NOT FOUND
C2349934|T033|HT|V89.0|ICD9CM|Suspected maternal and fetal conditions not found|Suspected maternal and fetal conditions not found
C2349926|T033|AB|V89.01|ICD9CM|Sus amntc cav/mem nt fnd|Sus amntc cav/mem nt fnd
C2349926|T033|PT|V89.01|ICD9CM|Suspected problem with amniotic cavity and membrane not found|Suspected problem with amniotic cavity and membrane not found
C2349929|T033|AB|V89.02|ICD9CM|Sus placentl prob nt fnd|Sus placentl prob nt fnd
C2349929|T033|PT|V89.02|ICD9CM|Suspected placental problem not found|Suspected placental problem not found
C2349930|T033|AB|V89.03|ICD9CM|Sus fetal anomaly nt fnd|Sus fetal anomaly nt fnd
C2349930|T033|PT|V89.03|ICD9CM|Suspected fetal anomaly not found|Suspected fetal anomaly not found
C2349931|T033|AB|V89.04|ICD9CM|Sus fetal growth not fnd|Sus fetal growth not fnd
C2349931|T033|PT|V89.04|ICD9CM|Suspected problem with fetal growth not found|Suspected problem with fetal growth not found
C2349932|T033|AB|V89.05|ICD9CM|Sus cervcl shortn nt fnd|Sus cervcl shortn nt fnd
C2349932|T033|PT|V89.05|ICD9CM|Suspected cervical shortening not found|Suspected cervical shortening not found
C2349933|T033|AB|V89.09|ICD9CM|Oth sus mat/ftl nt fnd|Oth sus mat/ftl nt fnd
C2349933|T033|PT|V89.09|ICD9CM|Other suspected maternal and fetal condition not found|Other suspected maternal and fetal condition not found
C0865505|T037|HT|V90|ICD9CM|Retained foreign body|Retained foreign body
C0865505|T037|HT|V90-V90.99|ICD9CM|RETAINED FOREIGN BODY|RETAINED FOREIGN BODY
C2921322|T033|HT|V90.0|ICD9CM|Retained radioactive fragment|Retained radioactive fragment
C2921323|T033|AB|V90.01|ICD9CM|Retain deplete uran frag|Retain deplete uran frag
C2921323|T033|PT|V90.01|ICD9CM|Retained depleted uranium fragments|Retained depleted uranium fragments
C2921325|T033|PT|V90.09|ICD9CM|Other retained radioactive fragments|Other retained radioactive fragments
C2921325|T033|AB|V90.09|ICD9CM|Retain radioac frag NEC|Retain radioac frag NEC
C2921327|T033|HT|V90.1|ICD9CM|Retained metal fragments|Retained metal fragments
C2921327|T033|AB|V90.10|ICD9CM|Retained metal frag NOS|Retained metal frag NOS
C2921327|T033|PT|V90.10|ICD9CM|Retained metal fragments, unspecified|Retained metal fragments, unspecified
C2921328|T033|AB|V90.11|ICD9CM|Retain magnet metal frag|Retain magnet metal frag
C2921328|T033|PT|V90.11|ICD9CM|Retained magnetic metal fragments|Retained magnetic metal fragments
C2921329|T033|AB|V90.12|ICD9CM|Retain nonmag meta frag|Retain nonmag meta frag
C2921329|T033|PT|V90.12|ICD9CM|Retained nonmagnetic metal fragments|Retained nonmagnetic metal fragments
C2921333|T033|AB|V90.2|ICD9CM|Retain plastic fragments|Retain plastic fragments
C2921333|T033|PT|V90.2|ICD9CM|Retained plastic fragments|Retained plastic fragments
C2921334|T033|HT|V90.3|ICD9CM|Retained organic fragments|Retained organic fragments
C2921335|T033|PT|V90.31|ICD9CM|Retained animal quills or spines|Retained animal quills or spines
C2921335|T033|AB|V90.31|ICD9CM|Retained quills/spines|Retained quills/spines
C4721538|T033|PT|V90.32|ICD9CM|Retained tooth|Retained tooth
C4721538|T033|AB|V90.32|ICD9CM|Retained tooth|Retained tooth
C2921337|T033|PT|V90.33|ICD9CM|Retained wood fragments|Retained wood fragments
C2921337|T033|AB|V90.33|ICD9CM|Retained wood fragments|Retained wood fragments
C2921338|T033|PT|V90.39|ICD9CM|Other retained organic fragments|Other retained organic fragments
C2921338|T033|AB|V90.39|ICD9CM|Retain organic frag NEC|Retain organic frag NEC
C2921339|T033|HT|V90.8|ICD9CM|Other specified retained foreign body|Other specified retained foreign body
C2921340|T033|AB|V90.81|ICD9CM|Retained glass fragments|Retained glass fragments
C2921340|T033|PT|V90.81|ICD9CM|Retained glass fragments|Retained glass fragments
C2921342|T033|AB|V90.83|ICD9CM|Retain stone/crystl frag|Retain stone/crystl frag
C2921342|T033|PT|V90.83|ICD9CM|Retained stone or crystalline fragments|Retained stone or crystalline fragments
C2921339|T033|PT|V90.89|ICD9CM|Other specified retained foreign body|Other specified retained foreign body
C2921339|T033|AB|V90.89|ICD9CM|Retain FB NEC|Retain FB NEC
C2921343|T033|AB|V90.9|ICD9CM|Retain FB, mat NOS|Retain FB, mat NOS
C2921343|T033|PT|V90.9|ICD9CM|Retained foreign body, unspecified material|Retained foreign body, unspecified material
C2921344|T033|HT|V91|ICD9CM|Multiple gestation placenta status|Multiple gestation placenta status
C2921344|T033|HT|V91-V91.99|ICD9CM|MULTIPLE GESTATION PLACENTA STATUS|MULTIPLE GESTATION PLACENTA STATUS
C2921345|T033|HT|V91.0|ICD9CM|Twin gestation placenta status|Twin gestation placenta status
C2921346|T033|AB|V91.00|ICD9CM|Twin gest-plac/sac NOS|Twin gest-plac/sac NOS
C2921346|T033|PT|V91.00|ICD9CM|Twin gestation, unspecified number of placenta, unspecified number of amniotic sacs|Twin gestation, unspecified number of placenta, unspecified number of amniotic sacs
C2921347|T033|AB|V91.01|ICD9CM|Twin gest-monochr/monoam|Twin gest-monochr/monoam
C2921347|T033|PT|V91.01|ICD9CM|Twin gestation, monochorionic/monoamniotic (one placenta, one amniotic sac)|Twin gestation, monochorionic/monoamniotic (one placenta, one amniotic sac)
C2921348|T033|AB|V91.02|ICD9CM|Twin gest-monochr/diamni|Twin gest-monochr/diamni
C2921348|T033|PT|V91.02|ICD9CM|Twin gestation, monochorionic/diamniotic (one placenta, two amniotic sacs)|Twin gestation, monochorionic/diamniotic (one placenta, two amniotic sacs)
C2921349|T033|AB|V91.03|ICD9CM|Twin gest-dich/diamniotc|Twin gest-dich/diamniotc
C2921349|T033|PT|V91.03|ICD9CM|Twin gestation, dichorionic/diamniotic (two placentae, two amniotic sacs)|Twin gestation, dichorionic/diamniotic (two placentae, two amniotic sacs)
C2921350|T033|AB|V91.09|ICD9CM|Twin gest-plac/sac undet|Twin gest-plac/sac undet
C2921350|T033|PT|V91.09|ICD9CM|Twin gestation, unable to determine number of placenta and number of amniotic sacs|Twin gestation, unable to determine number of placenta and number of amniotic sacs
C2921351|T033|HT|V91.1|ICD9CM|Triplet gestation placenta status|Triplet gestation placenta status
C2921352|T033|AB|V91.10|ICD9CM|Tripl gest-plac/sac NOS|Tripl gest-plac/sac NOS
C2921352|T033|PT|V91.10|ICD9CM|Triplet gestation, unspecified number of placenta and unspecified number of amniotic sacs|Triplet gestation, unspecified number of placenta and unspecified number of amniotic sacs
C2921353|T033|AB|V91.11|ICD9CM|Triplet gest 2+ monochor|Triplet gest 2+ monochor
C2921353|T033|PT|V91.11|ICD9CM|Triplet gestation, with two or more monochorionic fetuses|Triplet gestation, with two or more monochorionic fetuses
C2921354|T033|AB|V91.12|ICD9CM|Triplet gest 2+ monoamn|Triplet gest 2+ monoamn
C2921354|T033|PT|V91.12|ICD9CM|Triplet gestation, with two or more monoamniotic fetuses|Triplet gestation, with two or more monoamniotic fetuses
C2921355|T033|AB|V91.19|ICD9CM|Tripl gest-plac/sac und|Tripl gest-plac/sac und
C2921355|T033|PT|V91.19|ICD9CM|Triplet gestation, unable to determine number of placenta and number of amniotic sacs|Triplet gestation, unable to determine number of placenta and number of amniotic sacs
C2921356|T033|HT|V91.2|ICD9CM|Quadruplet gestation placenta status|Quadruplet gestation placenta status
C2921357|T033|AB|V91.20|ICD9CM|Quad gest-plac/sac NOS|Quad gest-plac/sac NOS
C2921357|T033|PT|V91.20|ICD9CM|Quadruplet gestation, unspecified number of placenta and unspecified number of amniotic sacs|Quadruplet gestation, unspecified number of placenta and unspecified number of amniotic sacs
C2921358|T033|AB|V91.21|ICD9CM|Quad gest 2+ monochorion|Quad gest 2+ monochorion
C2921358|T033|PT|V91.21|ICD9CM|Quadruplet gestation, with two or more monochorionic fetuses|Quadruplet gestation, with two or more monochorionic fetuses
C2921359|T033|AB|V91.22|ICD9CM|Quad gest 2+ monoamniotc|Quad gest 2+ monoamniotc
C2921359|T033|PT|V91.22|ICD9CM|Quadruplet gestation, with two or more monoamniotic fetuses|Quadruplet gestation, with two or more monoamniotic fetuses
C2921360|T033|AB|V91.29|ICD9CM|Quad gest-plac/sac undet|Quad gest-plac/sac undet
C2921360|T033|PT|V91.29|ICD9CM|Quadruplet gestation, unable to determine number of placenta and number of amniotic sacs|Quadruplet gestation, unable to determine number of placenta and number of amniotic sacs
C2921361|T033|HT|V91.9|ICD9CM|Other specified multiple gestation placenta status|Other specified multiple gestation placenta status
C2921363|T033|AB|V91.90|ICD9CM|Mult gest-plac/sac NOS|Mult gest-plac/sac NOS
C2921364|T033|AB|V91.91|ICD9CM|Mult gest 2+ monochr NEC|Mult gest 2+ monochr NEC
C2921364|T033|PT|V91.91|ICD9CM|Other specified multiple gestation, with two or more monochorionic fetuses|Other specified multiple gestation, with two or more monochorionic fetuses
C2921365|T033|AB|V91.92|ICD9CM|Mult gest 2+ monoamn NEC|Mult gest 2+ monoamn NEC
C2921365|T033|PT|V91.92|ICD9CM|Other specified multiple gestation, with two or more monoamniotic fetuses|Other specified multiple gestation, with two or more monoamniotic fetuses
C2921366|T033|AB|V91.99|ICD9CM|Mult gest-plac/sac undet|Mult gest-plac/sac undet

C0000737|ICD9CM|HT|789.0|Abdominal pain
C0000737|ICD9CM|PT|789.00|Abdominal pain, unspecified site
C0000737|ICD9CM|AB|789.00|Abdmnal pain unspcf site
C0000768|ICD9CM|HT|740-759.99|CONGENITAL ANOMALIES
C0000768|ICD9CM|AB|759.9|Congenital anomaly NOS
C0000768|ICD9CM|PT|759.9|Congenital anomaly, unspecified
C0000770|ICD9CM|PT|520.2|Abnormalities of size and form of teeth
C0000770|ICD9CM|AB|520.2|Abnormal tooth size/form
C0000774|ICD9CM|PT|251.5|Abnormality of secretion of gastrin
C0000774|ICD9CM|AB|251.5|Abnorm secretion gastrin
C0000786|ICD9CM|HT|634|Spontaneous abortion
C0000804|ICD9CM|HT|636|Illegally induced abortion
C0000814|ICD9CM|AB|632|Missed abortion
C0000814|ICD9CM|PT|632|Missed abortion
C0000821|ICD9CM|HT|640.0|Threatened abortion
C0000821|ICD9CM|PT|640.03|Threatened abortion, antepartum condition or complication
C0000821|ICD9CM|AB|640.03|Threaten abort-antepart
C0000827|ICD9CM|PT|919.0|Abrasion or friction burn of other, multiple, and unspecified sites, without mention of infection
C0000827|ICD9CM|AB|919.0|Abrasion NEC
C0000832|ICD9CM|HT|641.2|Premature separation of placenta
C0000832|ICD9CM|PT|641.20|Premature separation of placenta, unspecified as to episode of care or not applicable
C0000832|ICD9CM|AB|641.20|Prem separ placen-unspec
C0000908|ICD9CM|PT|E924.1|Accident caused by caustic and corrosive substances
C0000908|ICD9CM|AB|E924.1|Accid-caustic substance
C0000909|ICD9CM|PT|E900.0|Accident caused by excessive heat due to weather conditions
C0000909|ICD9CM|AB|E900.0|Excessive heat: weather
C0000912|ICD9CM|PT|E899|Accident caused by unspecified fire
C0000912|ICD9CM|AB|E899|Fire accident NOS
C0000914|ICD9CM|PT|E902.2|Accident due to changes in air pressure due to diving
C0000914|ICD9CM|AB|E902.2|Air press change: diving
C0000915|ICD9CM|PT|E907|Accident due to lightning
C0000915|ICD9CM|AB|E907|Acc due to lightning
C0000916|ICD9CM|PT|E902.0|Accident due to residence or prolonged visit at high altitude
C0000916|ICD9CM|AB|E902.0|High altitude residence
C0000921|ICD9CM|HT|E880-E888.9|ACCIDENTAL FALLS
C0000922|ICD9CM|PT|E913.9|Accidental mechanical suffocation by unspecified means
C0000922|ICD9CM|AB|E913.9|Suffocation NOS
C0000923|ICD9CM|PT|E865.2|Accidental poisoning from other fish
C0000923|ICD9CM|AB|E865.2|Acc poison-fish NEC
C0000926|ICD9CM|PT|E900.9|Accidents due to excessive heat of unspecified origin
C0000926|ICD9CM|AB|E900.9|Excessive heat NOS
C0000929|ICD9CM|PT|E849.0|Home accidents
C0000929|ICD9CM|AB|E849.0|Accident in home
C0001075|ICD9CM|AB|536.0|Achlorhydria
C0001075|ICD9CM|PT|536.0|Achlorhydria
C0001122|ICD9CM|AB|276.2|Acidosis
C0001122|ICD9CM|PT|276.2|Acidosis
C0001163|ICD9CM|PT|388.5|Disorders of acoustic nerve
C0001163|ICD9CM|AB|388.5|Acoustic nerve disorders
C0001169|ICD9CM|PT|286.7|Acquired coagulation factor deficiency
C0001169|ICD9CM|AB|286.7|Acq coagul factor defic
C0001170|ICD9CM|PT|380.32|Acquired deformities of auricle or pinna
C0001170|ICD9CM|AB|380.32|Acq deform auricle/pinna
C0001171|ICD9CM|PT|738.3|Acquired deformity of chest and rib
C0001171|ICD9CM|AB|738.3|Acq chest deformity
C0001261|ICD9CM|AB|039.9|Actinomycosis NOS
C0001261|ICD9CM|PT|039.9|Actinomycotic infection of unspecified site
C0001261|ICD9CM|HT|039|Actinomycotic infections
C0001263|ICD9CM|AB|039.2|Abdominal actinomycosis
C0001263|ICD9CM|PT|039.2|Abdominal actinomycotic infection
C0001264|ICD9CM|PT|039.3|Cervicofacial actinomycotic infection
C0001264|ICD9CM|AB|039.3|Cervicofac actinomycosis
C0001265|ICD9CM|PT|039.8|Actinomycotic infection of other specified sites
C0001265|ICD9CM|AB|039.8|Actinomycosis NEC
C0001301|ICD9CM|AB|99.91|Anesthesia acupuncture
C0001301|ICD9CM|PT|99.91|Acupuncture for anesthesia
C0001306|ICD9CM|PT|571.1|Acute alcoholic hepatitis
C0001306|ICD9CM|AB|571.1|Ac alcoholic hepatitis
C0001308|ICD9CM|PT|570|Acute and subacute necrosis of liver
C0001308|ICD9CM|AB|570|Acute necrosis of liver
C0001309|ICD9CM|PT|372.05|Acute atopic conjunctivitis
C0001309|ICD9CM|AB|372.05|Ac atopic conjunctivitis
C0001311|ICD9CM|HT|466.1|Acute bronchiolitis
C0001317|ICD9CM|HT|207.0|Acute erythremia and erythroleukemia
C0001327|ICD9CM|HT|464.0|Acute laryngitis
C0001339|ICD9CM|AB|577.0|Acute pancreatitis
C0001339|ICD9CM|PT|577.0|Acute pancreatitis
C0001342|ICD9CM|PT|523.33|Acute periodontitis
C0001342|ICD9CM|AB|523.33|Acute periodontitis
C0001342|ICD9CM|HT|523.3|Aggressive and acute periodontitis
C0001344|ICD9CM|AB|462|Acute pharyngitis
C0001344|ICD9CM|PT|462|Acute pharyngitis
C0001360|ICD9CM|AB|245.0|Acute thyroiditis
C0001360|ICD9CM|PT|245.0|Acute thyroiditis
C0001361|ICD9CM|AB|463|Acute tonsillitis
C0001361|ICD9CM|PT|463|Acute tonsillitis
C0001363|ICD9CM|PT|557.0|Acute vascular insufficiency of intestine
C0001363|ICD9CM|AB|557.0|Ac vasc insuff intestine
C0001365|ICD9CM|PT|436|Acute, but ill-defined, cerebrovascular disease
C0001365|ICD9CM|AB|436|Cva
C0001425|ICD9CM|AB|28.6|Adenoidectomy
C0001425|ICD9CM|PT|28.6|Adenoidectomy without tonsillectomy
C0001485|ICD9CM|PT|079.0|Adenovirus infection in conditions classified elsewhere and of unspecified site
C0001485|ICD9CM|AB|079.0|Adenovirus infect NOS
C0001539|ICD9CM|PT|309.0|Adjustment disorder with depressed mood
C0001539|ICD9CM|AB|309.0|Adjustmnt dis w depressn
C0001540|ICD9CM|PT|309.3|Adjustment disorder with disturbance of conduct
C0001540|ICD9CM|AB|309.3|Adjust disor/dis conduct
C0001541|ICD9CM|PT|309.4|Adjustment disorder with mixed disturbance of emotions and conduct
C0001541|ICD9CM|AB|309.4|Adj dis-emotion/conduct
C0001621|ICD9CM|PT|255.9|Unspecified disorder of adrenal glands
C0001621|ICD9CM|AB|255.9|Adrenal disorder NOS
C0001621|ICD9CM|HT|255|Disorders of adrenal glands
C0001815|ICD9CM|PT|238.76|Myelofibrosis with myeloid metaplasia
C0001815|ICD9CM|AB|238.76|Myelofi w myelo metaplas
C0001819|ICD9CM|PT|300.22|Agoraphobia without mention of panic attacks
C0001819|ICD9CM|AB|300.22|Agoraphobia w/o panic
C0001860|ICD9CM|AB|136.0|Ainhum
C0001860|ICD9CM|PT|136.0|Ainhum
C0001906|ICD9CM|AB|050.1|Alastrim
C0001906|ICD9CM|PT|050.1|Alastrim
C0001940|ICD9CM|PT|291.1|Alcohol-induced persisting amnestic disorder
C0001940|ICD9CM|AB|291.1|Alcohol amnestic disordr
C0001950|ICD9CM|PT|291.4|Idiosyncratic alcohol intoxication
C0001950|ICD9CM|AB|291.4|Pathologic alcohol intox
C0001957|ICD9CM|PT|291.0|Alcohol withdrawal delirium
C0001957|ICD9CM|AB|291.0|Delirium tremens
C0001973|ICD9CM|HT|303|Alcohol dependence syndrome
C0002018|ICD9CM|AB|315.01|Alexia
C0002018|ICD9CM|PT|315.01|Alexia
C0002019|ICD9CM|AB|784.61|Alexia and dyslexia
C0002019|ICD9CM|PT|784.61|Alexia and dyslexia
C0002063|ICD9CM|AB|276.3|Alkalosis
C0002063|ICD9CM|PT|276.3|Alkalosis
C0002170|ICD9CM|HT|704.0|Alopecia
C0002170|ICD9CM|AB|704.00|Alopecia NOS
C0002170|ICD9CM|PT|704.00|Alopecia, unspecified
C0002171|ICD9CM|AB|704.01|Alopecia areata
C0002171|ICD9CM|PT|704.01|Alopecia areata
C0002181|ICD9CM|AB|091.82|Syphilitic alopecia
C0002181|ICD9CM|PT|091.82|Syphilitic alopecia
C0002312|ICD9CM|PT|282.43|Alpha thalassemia
C0002312|ICD9CM|AB|282.43|Alpha thalassemia
C0002390|ICD9CM|HT|495|Extrinsic allergic alveolitis
C0002390|ICD9CM|PT|495.9|Unspecified allergic alveolitis and pneumonitis
C0002390|ICD9CM|AB|495.9|Allerg alveol/pneum NOS
C0002393|ICD9CM|AB|24.5|Alveoloplasty
C0002393|ICD9CM|PT|24.5|Alveoloplasty
C0002395|ICD9CM|AB|331.0|Alzheimer's disease
C0002395|ICD9CM|PT|331.0|Alzheimer's disease
C0002418|ICD9CM|AB|368.00|Amblyopia NOS
C0002418|ICD9CM|PT|368.00|Amblyopia, unspecified
C0002438|ICD9CM|HT|006|Amebiasis
C0002438|ICD9CM|AB|006.9|Amebiasis NOS
C0002438|ICD9CM|PT|006.9|Amebiasis, unspecified
C0002453|ICD9CM|AB|626.0|Absence of menstruation
C0002453|ICD9CM|PT|626.0|Absence of menstruation
C0002514|ICD9CM|HT|270|Disorders of amino-acid transport and metabolism
C0002514|ICD9CM|PT|270.9|Unspecified disorder of amino-acid metabolism
C0002514|ICD9CM|AB|270.9|Dis amino-acid metab NOS
C0002625|ICD9CM|PT|294.0|Amnestic disorder in conditions classified elsewhere
C0002625|ICD9CM|AB|294.0|Amnestic disord oth dis
C0002627|ICD9CM|AB|75.1|Diagnostic amniocentesis
C0002627|ICD9CM|PT|75.1|Diagnostic amniocentesis
C0002631|ICD9CM|HT|658.4|Infection of amniotic cavity
C0002631|ICD9CM|PT|658.40|Infection of amniotic cavity, unspecified as to episode of care or not applicable
C0002631|ICD9CM|AB|658.40|Amniotic infection-unsp
C0002632|ICD9CM|AB|75.31|Amnioscopy
C0002632|ICD9CM|PT|75.31|Amnioscopy
C0002688|ICD9CM|AB|84.91|Amputation NOS
C0002688|ICD9CM|PT|84.91|Amputation, not otherwise specified
C0002691|ICD9CM|AB|84.17|Above knee amputation
C0002691|ICD9CM|PT|84.17|Amputation above knee
C0002726|ICD9CM|HT|277.3|Amyloidosis
C0002726|ICD9CM|AB|277.30|Amyloidosis NOS
C0002726|ICD9CM|PT|277.30|Amyloidosis, unspecified
C0002736|ICD9CM|PT|335.20|Amyotrophic lateral sclerosis
C0002736|ICD9CM|AB|335.20|Amyotrophic sclerosis
C0002753|ICD9CM|PT|569.0|Anal and rectal polyp
C0002753|ICD9CM|AB|569.0|Anal & rectal polyp
C0002758|ICD9CM|AB|569.42|Anal or rectal pain
C0002758|ICD9CM|PT|569.42|Anal or rectal pain
C0002871|ICD9CM|AB|285.9|Anemia NOS
C0002871|ICD9CM|PT|285.9|Anemia, unspecified
C0002873|ICD9CM|HT|285.2|Anemia of chronic disease
C0002874|ICD9CM|AB|284.9|Aplastic anemia NOS
C0002874|ICD9CM|PT|284.9|Aplastic anemia, unspecified
C0002879|ICD9CM|HT|283|Acquired hemolytic anemias
C0002879|ICD9CM|PT|283.9|Acquired hemolytic anemia, unspecified
C0002879|ICD9CM|AB|283.9|Acq hemolytic anemia NOS
C0002880|ICD9CM|PT|283.0|Autoimmune hemolytic anemias
C0002880|ICD9CM|AB|283.0|Autoimmun hemolytic anem
C0002881|ICD9CM|HT|282|Hereditary hemolytic anemias
C0002881|ICD9CM|PT|282.9|Hereditary hemolytic anemia, unspecified
C0002881|ICD9CM|AB|282.9|Hered hemolytic anem NOS
C0002892|ICD9CM|AB|281.0|Pernicious anemia
C0002892|ICD9CM|PT|281.0|Pernicious anemia
C0002895|ICD9CM|HT|282.6|Sickle-cell disease
C0002895|ICD9CM|AB|282.60|Sickle cell disease NOS
C0002895|ICD9CM|PT|282.60|Sickle-cell disease, unspecified
C0002896|ICD9CM|AB|285.0|Sideroblastic anemia
C0002896|ICD9CM|PT|285.0|Sideroblastic anemia
C0002899|ICD9CM|PT|282.2|Anemias due to disorders of glutathione metabolism
C0002899|ICD9CM|AB|282.2|Glutathione dis anemia
C0002902|ICD9CM|AB|740.0|Anencephalus
C0002902|ICD9CM|PT|740.0|Anencephalus
C0002940|ICD9CM|AB|442.9|Aneurysm NOS
C0002940|ICD9CM|PT|442.9|Aneurysm of unspecified site
C0002945|ICD9CM|HT|442.8|Aneurysm of other specified artery
C0002946|ICD9CM|AB|442.89|Aneurysm NEC
C0002946|ICD9CM|PT|442.89|Aneurysm of other specified artery
C0002962|ICD9CM|HT|413|Angina pectoris
C0002963|ICD9CM|AB|413.1|Prinzmetal angina
C0002963|ICD9CM|PT|413.1|Prinzmetal angina
C0002965|ICD9CM|PT|411.1|Intermediate coronary syndrome
C0002965|ICD9CM|AB|411.1|Intermed coronary synd
C0002971|ICD9CM|AB|88.50|Angiocardiography NOS
C0002971|ICD9CM|PT|88.50|Angiocardiography, not otherwise specified
C0002983|ICD9CM|PT|363.43|Angioid streaks of choroid
C0002983|ICD9CM|AB|363.43|Angioid streaks, choroid
C0002998|ICD9CM|AB|39.30|Suture of vessel NOS
C0002998|ICD9CM|PT|39.30|Suture of unspecified blood vessel
C0003028|ICD9CM|AB|705.0|Anhidrosis
C0003028|ICD9CM|PT|705.0|Anhidrosis
C0003044|ICD9CM|AB|E906.5|Animal bite NOS
C0003044|ICD9CM|PT|E906.5|Bite by unspecified animal
C0003076|ICD9CM|AB|743.45|Aniridia
C0003076|ICD9CM|PT|743.45|Aniridia
C0003078|ICD9CM|AB|367.32|Aniseikonia
C0003078|ICD9CM|PT|367.32|Aniseikonia
C0003079|ICD9CM|AB|379.41|Anisocoria
C0003079|ICD9CM|PT|379.41|Anisocoria
C0003081|ICD9CM|AB|367.31|Anisometropia
C0003081|ICD9CM|PT|367.31|Anisometropia
C0003089|ICD9CM|HT|720|Ankylosing spondylitis and other inflammatory spondylopathies
C0003090|ICD9CM|HT|718.5|Ankylosis of joint
C0003090|ICD9CM|PT|718.50|Ankylosis of joint, site unspecified
C0003090|ICD9CM|AB|718.50|Ankylosis-unspec
C0003110|ICD9CM|HT|524.1|Anomalies of relationship of jaw to cranial base
C0003110|ICD9CM|PT|524.10|Anomalies of relationship of jaw to cranial base, unspecified anomaly
C0003110|ICD9CM|AB|524.10|Unspcf anm jaw cranl bse
C0003119|ICD9CM|HT|743.0|Anophthalmos
C0003119|ICD9CM|PT|743.00|Clinical anophthalmos, unspecified
C0003119|ICD9CM|AB|743.00|Clinic anophthalmos NOS
C0003123|ICD9CM|AB|783.0|Anorexia
C0003123|ICD9CM|PT|783.0|Anorexia
C0003125|ICD9CM|AB|307.1|Anorexia nervosa
C0003125|ICD9CM|PT|307.1|Anorexia nervosa
C0003132|ICD9CM|AB|348.1|Anoxic brain damage
C0003132|ICD9CM|PT|348.1|Anoxic brain damage
C0003165|ICD9CM|AB|500|Coal workers' pneumocon
C0003165|ICD9CM|PT|500|Coal workers' pneumoconiosis
C0003175|ICD9CM|HT|022|Anthrax
C0003175|ICD9CM|AB|022.9|Anthrax NOS
C0003175|ICD9CM|PT|022.9|Anthrax, unspecified
C0003177|ICD9CM|AB|022.0|Cutaneous anthrax
C0003177|ICD9CM|PT|022.0|Cutaneous anthrax
C0003431|ICD9CM|PT|301.7|Antisocial personality disorder
C0003431|ICD9CM|AB|301.7|Antisocial personality
C0003477|ICD9CM|PT|309.21|Separation anxiety disorder
C0003477|ICD9CM|AB|309.21|Separation anxiety
C0003492|ICD9CM|AB|747.10|Coarctation of aorta
C0003492|ICD9CM|HT|747.1|Coarctation of aorta
C0003492|ICD9CM|PT|747.10|Coarctation of aorta (preductal) (postductal)
C0003511|ICD9CM|AB|093.1|Syphilitic aortitis
C0003511|ICD9CM|PT|093.1|Syphilitic aortitis
C0003515|ICD9CM|PT|88.42|Aortography
C0003515|ICD9CM|AB|88.42|Contrast aortogram
C0003534|ICD9CM|AB|379.31|Aphakia
C0003534|ICD9CM|PT|379.31|Aphakia
C0003537|ICD9CM|AB|784.3|Aphasia
C0003537|ICD9CM|PT|784.3|Aphasia
C0003564|ICD9CM|AB|784.41|Aphonia
C0003564|ICD9CM|PT|784.41|Aphonia
C0003571|ICD9CM|AB|23.73|Apicoectomy
C0003571|ICD9CM|PT|23.73|Apicoectomy
C0003578|ICD9CM|AB|786.03|Apnea
C0003578|ICD9CM|PT|786.03|Apnea
C0003611|ICD9CM|HT|47.0|Appendectomy
C0003615|ICD9CM|HT|540-543.99|APPENDICITIS
C0003615|ICD9CM|AB|541|Appendicitis NOS
C0003615|ICD9CM|PT|541|Appendicitis, unqualified
C0003626|ICD9CM|PT|23.41|Application of crown
C0003626|ICD9CM|AB|23.41|Crown application
C0003627|ICD9CM|PT|93.57|Application of other wound dressing
C0003627|ICD9CM|AB|93.57|Dressing of wound NEC
C0003721|ICD9CM|HT|065|Arthropod-borne hemorrhagic fever
C0003721|ICD9CM|PT|065.9|Arthropod-borne hemorrhagic fever, unspecified
C0003721|ICD9CM|AB|065.9|Arthropod hem fever NOS
C0003723|ICD9CM|HT|060-066.99|ARTHROPOD-BORNE VIRAL DISEASES
C0003723|ICD9CM|PT|066.9|Arthropod-borne viral disease, unspecified
C0003723|ICD9CM|AB|066.9|Arthropod virus NOS
C0003811|ICD9CM|HT|427|Cardiac dysrhythmias
C0003811|ICD9CM|AB|427.9|Cardiac dysrhythmia NOS
C0003811|ICD9CM|PT|427.9|Cardiac dysrhythmia, unspecified
C0003844|ICD9CM|HT|88.4|Arteriography using contrast material
C0003860|ICD9CM|AB|447.6|Arteritis NOS
C0003860|ICD9CM|PT|447.6|Arteritis, unspecified
C0003862|ICD9CM|AB|719.40|Joint pain-unspec
C0003862|ICD9CM|HT|719.4|Pain in joint
C0003862|ICD9CM|PT|719.40|Pain in joint, site unspecified
C0003868|ICD9CM|HT|274.0|Gouty arthropathy
C0003868|ICD9CM|AB|274.00|Gouty arthropathy NOS
C0003868|ICD9CM|PT|274.00|Gouty arthropathy, unspecified
C0003869|ICD9CM|AB|711.90|Inf arthritis NOS-unspec
C0003869|ICD9CM|HT|711.0|Pyogenic arthritis
C0003869|ICD9CM|HT|711.9|Unspecified infective arthritis
C0003869|ICD9CM|PT|711.90|Unspecified infective arthritis, site unspecified
C0003872|ICD9CM|AB|696.0|Psoriatic arthropathy
C0003872|ICD9CM|PT|696.0|Psoriatic arthropathy
C0003873|ICD9CM|AB|714.0|Rheumatoid arthritis
C0003873|ICD9CM|PT|714.0|Rheumatoid arthritis
C0003881|ICD9CM|AB|81.20|Arthrodesis NOS
C0003881|ICD9CM|PT|81.20|Arthrodesis of unspecified joint
C0003883|ICD9CM|PT|81.29|Arthrodesis of other specified joints
C0003883|ICD9CM|AB|81.29|Arthrodesis NEC
C0003885|ICD9CM|AB|88.32|Contrast arthrogram
C0003885|ICD9CM|PT|88.32|Contrast arthrogram
C0003892|ICD9CM|PT|713.5|Arthropathy associated with neurological disorders
C0003892|ICD9CM|AB|713.5|Arthropathy w nerve dis
C0003904|ICD9CM|HT|80.2|Arthroscopy
C0003906|MTH|PN|NOCODE|Arthroscopy NEC in ICD9CM_2014
C0003906|ICD9CM|AB|80.29|Arthroscopy NEC
C0003906|ICD9CM|PT|80.29|Arthroscopy, other specified sites
C0003907|ICD9CM|PT|995.21|Arthus phenomenon
C0003907|ICD9CM|AB|995.21|Arthus phenomenon
C0003949|ICD9CM|AB|501|Asbestosis
C0003949|ICD9CM|PT|501|Asbestosis
C0003950|ICD9CM|AB|127.0|Ascariasis
C0003950|ICD9CM|PT|127.0|Ascariasis
C0003962|ICD9CM|HT|789.5|Ascites
C0003969|ICD9CM|AB|267|Ascorbic acid deficiency
C0003969|ICD9CM|PT|267|Ascorbic acid deficiency
C0003977|ICD9CM|PT|733.42|Aseptic necrosis of head and neck of femur
C0003977|ICD9CM|AB|733.42|Aseptic necrosis femur
C0004030|ICD9CM|AB|117.3|Aspergillosis
C0004030|ICD9CM|PT|117.3|Aspergillosis
C0004031|ICD9CM|PT|518.6|Allergic bronchopulmonary aspergillosis
C0004031|ICD9CM|AB|518.6|Alrgc brncpul asprglosis
C0004044|ICD9CM|AB|799.01|Asphyxia
C0004044|ICD9CM|PT|799.01|Asphyxia
C0004045|ICD9CM|PT|768.9|Unspecified severity of birth asphyxia in liveborn infant
C0004045|ICD9CM|AB|768.9|Birth asphyxia NOS
C0004050|ICD9CM|PT|69.51|Aspiration curettage of uterus for termination of pregnancy
C0004050|ICD9CM|AB|69.51|Aspirat curet-preg termi
C0004063|ICD9CM|AB|E968.9|Assault NOS
C0004063|ICD9CM|PT|E968.9|Assault by unspecified means
C0004096|ICD9CM|HT|493|Asthma
C0004096|ICD9CM|HT|493.9|Asthma, unspecified
C0004106|ICD9CM|HT|367.2|Astigmatism
C0004106|ICD9CM|AB|367.20|Astigmatism NOS
C0004106|ICD9CM|PT|367.20|Astigmatism, unspecified
C0004144|ICD9CM|AB|518.0|Pulmonary collapse
C0004144|ICD9CM|PT|518.0|Pulmonary collapse
C0004153|ICD9CM|HT|440|Atherosclerosis
C0004155|ICD9CM|PT|440.8|Atherosclerosis of other specified arteries
C0004155|ICD9CM|AB|440.8|Atherosclerosis NEC
C0004187|ICD9CM|HT|691|Atopic dermatitis and related conditions
C0004238|ICD9CM|AB|427.31|Atrial fibrillation
C0004238|ICD9CM|PT|427.31|Atrial fibrillation
C0004239|ICD9CM|AB|427.32|Atrial flutter
C0004239|ICD9CM|PT|427.32|Atrial flutter
C0004245|ICD9CM|PT|426.10|Atrioventricular block, unspecified
C0004245|ICD9CM|AB|426.10|Atriovent block NOS
C0004269|ICD9CM|HT|314.0|Attention deficit disorder of childhood
C0004286|ICD9CM|AB|95.41|Audiometry
C0004286|ICD9CM|PT|95.41|Audiometry
C0004352|ICD9CM|HT|299.0|Autistic disorder
C0004398|ICD9CM|AB|89.8|Autopsy
C0004398|ICD9CM|PT|89.8|Autopsy
C0004402|ICD9CM|HT|758.3|Autosomal deletion syndromes
C0004444|ICD9CM|PT|301.82|Avoidant personality disorder
C0004444|ICD9CM|AB|301.82|Avoidant personality dis
C0004445|ICD9CM|AB|871.3|Avulsion of eye
C0004445|ICD9CM|PT|871.3|Avulsion of eye
C0004509|ICD9CM|AB|606.0|Azoospermia
C0004509|ICD9CM|PT|606.0|Azoospermia
C0004576|ICD9CM|AB|088.82|Babesiosis
C0004576|ICD9CM|PT|088.82|Babesiosis
C0004604|ICD9CM|AB|724.5|Backache NOS
C0004604|ICD9CM|PT|724.5|Backache, unspecified
C0004606|ICD9CM|PT|362.03|Nonproliferative diabetic retinopathy NOS
C0004606|ICD9CM|PT|362.01|Background diabetic retinopathy
C0004606|ICD9CM|AB|362.01|Diabetic retinopathy NOS
C0004606|ICD9CM|AB|362.03|Nonprolf db retnoph NOS
C0004608|ICD9CM|PT|362.10|Background retinopathy, unspecified
C0004608|ICD9CM|AB|362.10|Backgrnd retinopathy NOS
C0004610|ICD9CM|AB|790.7|Bacteremia
C0004610|ICD9CM|PT|790.7|Bacteremia
C0004622|ICD9CM|PT|041.9|Bacterial infection, unspecified, in conditions classified elsewhere and of unspecified site
C0004622|ICD9CM|AB|041.9|Bacterial infection NOS
C0004622|ICD9CM|HT|041|Bacterial infection in conditions classified elsewhere and of unspecified site
C0004626|ICD9CM|AB|482.9|Bacterial pneumonia NOS
C0004626|ICD9CM|PT|482.9|Bacterial pneumonia, unspecified
C0004681|ICD9CM|AB|495.1|Bagassosis
C0004681|ICD9CM|PT|495.1|Bagassosis
C0004691|ICD9CM|AB|607.1|Balanoposthitis
C0004691|ICD9CM|PT|607.1|Balanoposthitis
C0004692|ICD9CM|AB|007.0|Balantidiasis
C0004692|ICD9CM|PT|007.0|Balantidiasis
C0004763|ICD9CM|AB|530.85|Barrett's esophagus
C0004763|ICD9CM|PT|530.85|Barrett's esophagus
C0004766|ICD9CM|PT|616.3|Abscess of Bartholin's gland
C0004766|ICD9CM|AB|616.3|Bartholin's glnd abscess
C0004767|ICD9CM|AB|616.2|Bartholin's gland cyst
C0004767|ICD9CM|PT|616.2|Cyst of Bartholin's gland
C0004771|ICD9CM|AB|088.0|Bartonellosis
C0004771|ICD9CM|PT|088.0|Bartonellosis
C0004775|ICD9CM|AB|255.13|Bartter's syndrome
C0004775|ICD9CM|PT|255.13|Bartter's syndrome
C0004795|ICD9CM|AB|E007.3|Baseball
C0004795|ICD9CM|PT|E007.3|Activities involving baseball
C0004812|ICD9CM|AB|435.0|Basilar artery syndrome
C0004812|ICD9CM|PT|435.0|Basilar artery syndrome
C0004818|ICD9CM|AB|E007.6|Basketball
C0004818|ICD9CM|PT|E007.6|Activities involving basketball
C0004933|ICD9CM|AB|94.33|Behavior therapy
C0004933|ICD9CM|PT|94.33|Behavior therapy
C0004943|ICD9CM|AB|136.1|Behcet's syndrome
C0004943|ICD9CM|PT|136.1|Behcet's syndrome
C0004991|ICD9CM|PT|211.3|Benign neoplasm of colon
C0004991|ICD9CM|AB|211.3|Benign neoplasm lg bowel
C0004992|ICD9CM|PT|225.1|Benign neoplasm of cranial nerves
C0004992|ICD9CM|AB|225.1|Benign neo cranial nerve
C0004994|ICD9CM|PT|213.1|Benign neoplasm of lower jaw bone
C0004994|ICD9CM|AB|213.1|Ben neo lower jaw bone
C0004997|ICD9CM|PT|220|Benign neoplasm of ovary
C0004997|ICD9CM|AB|220|Benign neoplasm ovary
C0004998|ICD9CM|HT|216|Benign neoplasm of skin
C0004998|ICD9CM|AB|216.9|Benign neoplasm skin NOS
C0004998|ICD9CM|PT|216.9|Benign neoplasm of skin, site unspecified
C0005122|ICD9CM|AB|265.0|Beriberi
C0005122|ICD9CM|PT|265.0|Beriberi
C0005283|ICD9CM|PT|282.44|Beta thalassemia
C0005283|ICD9CM|AB|282.44|Beta thalassemia
C0005411|ICD9CM|AB|751.61|Biliary atresia
C0005411|ICD9CM|PT|751.61|Biliary atresia
C0005417|ICD9CM|AB|576.4|Fistula of bile duct
C0005417|ICD9CM|PT|576.4|Fistula of bile duct
C0005424|ICD9CM|PT|576.9|Unspecified disorder of biliary tract
C0005424|ICD9CM|AB|576.9|Dis of biliary tract NOS
C0005461|ICD9CM|PT|368.30|Binocular vision disorder, unspecified
C0005461|ICD9CM|AB|368.30|Binocular vision dis NOS
C0005586|ICD9CM|AB|296.80|Bipolar disorder NOS
C0005586|ICD9CM|PT|296.80|Bipolar disorder, unspecified
C0005592|ICD9CM|AB|495.2|Bird-fanciers' lung
C0005592|ICD9CM|PT|495.2|Bird-fanciers' lung
C0005604|ICD9CM|HT|767|Birth trauma
C0005604|ICD9CM|AB|767.9|Birth trauma NOS
C0005604|ICD9CM|PT|767.9|Birth trauma, unspecified
C0005656|ICD9CM|PT|E906.3|Bite of other animal except arthropod
C0005656|ICD9CM|AB|E906.3|Animal bite NEC
C0005660|ICD9CM|PT|E928.3|Human bite
C0005660|ICD9CM|AB|E928.3|Human bite - accidental
C0005681|ICD9CM|AB|084.8|Blackwater fever
C0005681|ICD9CM|PT|084.8|Blackwater fever
C0005684|ICD9CM|HT|188|Malignant neoplasm of bladder
C0005684|ICD9CM|PT|188.9|Malignant neoplasm of bladder, part unspecified
C0005684|ICD9CM|AB|188.9|Malig neo bladder NOS
C0005686|ICD9CM|PT|596.9|Unspecified disorder of bladder
C0005686|ICD9CM|AB|596.9|Bladder disorder NOS
C0005689|ICD9CM|AB|753.5|Bladder exstrophy
C0005689|ICD9CM|PT|753.5|Exstrophy of urinary bladder
C0005694|ICD9CM|AB|596.0|Bladder neck obstruction
C0005694|ICD9CM|PT|596.0|Bladder neck obstruction
C0005697|ICD9CM|AB|596.54|Neurogenic bladder NOS
C0005697|ICD9CM|PT|596.54|Neurogenic bladder NOS
C0005700|ICD9CM|PT|993.4|Effects of air pressure caused by explosion
C0005700|ICD9CM|AB|993.4|Eff air press by explos
C0005716|ICD9CM|AB|116.0|Blastomycosis
C0005716|ICD9CM|PT|116.0|Blastomycosis
C0005716|ICD9CM|HT|116|Blastomycotic infection
C0005741|ICD9CM|HT|373.0|Blepharitis
C0005741|ICD9CM|AB|373.00|Blepharitis NOS
C0005741|ICD9CM|AB|373.9|Inflammation eyelid NOS
C0005741|ICD9CM|PT|373.9|Unspecified inflammation of eyelid
C0005741|ICD9CM|PT|373.00|Blepharitis, unspecified
C0005742|ICD9CM|AB|374.34|Blepharochalasis
C0005742|ICD9CM|PT|374.34|Blepharochalasis
C0005743|ICD9CM|HT|372.2|Blepharoconjunctivitis
C0005743|ICD9CM|PT|372.20|Blepharoconjunctivitis, unspecified
C0005743|ICD9CM|AB|372.20|Blepharoconjunctivit NOS
C0005744|ICD9CM|AB|374.46|Blepharophimosis
C0005744|ICD9CM|PT|374.46|Blepharophimosis
C0005745|ICD9CM|HT|374.3|Ptosis of eyelid
C0005745|ICD9CM|AB|374.30|Ptosis of eyelid NOS
C0005745|ICD9CM|PT|374.30|Ptosis of eyelid, unspecified
C0005746|ICD9CM|AB|08.52|Blepharorrhaphy
C0005746|ICD9CM|PT|08.52|Blepharorrhaphy
C0005747|ICD9CM|AB|333.81|Blepharospasm
C0005747|ICD9CM|PT|333.81|Blepharospasm
C0005750|ICD9CM|AB|579.2|Blind loop syndrome
C0005750|ICD9CM|PT|579.2|Blind loop syndrome
C0005761|ICD9CM|PT|919.2|Blister of other, multiple, and unspecified sites, without mention of infection
C0005761|ICD9CM|AB|919.2|Blister NEC
C0005779|ICD9CM|HT|286|Coagulation defects
C0005843|ICD9CM|AB|75.2|Intrauterine transfusion
C0005843|ICD9CM|PT|75.2|Intrauterine transfusion
C0005933|ICD9CM|HT|77.4|Biopsy of bone
C0005933|ICD9CM|AB|77.40|Bone biopsy NOS
C0005933|ICD9CM|PT|77.40|Biopsy of bone, unspecified site
C0005937|ICD9CM|HT|733.2|Cyst of bone
C0005937|ICD9CM|AB|733.20|Cyst of bone NOS
C0005937|ICD9CM|AB|733.21|Solitary bone cyst
C0005937|ICD9CM|PT|733.21|Solitary bone cyst
C0005937|ICD9CM|PT|733.20|Cyst of bone (localized), unspecified
C0005949|ICD9CM|HT|78.3|Limb lengthening procedures
C0005949|ICD9CM|PT|78.30|Limb lengthening procedures, unspecified site
C0005949|ICD9CM|AB|78.30|Limb lengthen proc NOS
C0005954|ICD9CM|AB|41.31|Bone marrow biopsy
C0005954|ICD9CM|PT|41.31|Biopsy of bone marrow
C0005961|ICD9CM|PT|41.00|Bone marrow transplant, not otherwise specified
C0005961|ICD9CM|AB|41.00|Bone marrow trnsplnt NOS
C0005976|ICD9CM|HT|78.0|Bone graft
C0005976|ICD9CM|AB|78.00|Bone graft NOS
C0005976|ICD9CM|PT|78.00|Bone graft, unspecified site
C0006012|ICD9CM|PT|301.83|Borderline personality disorder
C0006012|ICD9CM|AB|301.83|Borderline personality
C0006060|ICD9CM|AB|082.1|Boutonneuse fever
C0006060|ICD9CM|PT|082.1|Boutonneuse fever
C0006080|ICD9CM|AB|E008.0|Boxing
C0006080|ICD9CM|PT|E008.0|Activities involving boxing
C0006091|ICD9CM|AB|353.0|Brachial plexus lesions
C0006091|ICD9CM|PT|353.0|Brachial plexus lesions
C0006107|ICD9CM|HT|850|Concussion
C0006107|ICD9CM|AB|850.9|Concussion NOS
C0006107|ICD9CM|PT|850.9|Concussion, unspecified
C0006110|ICD9CM|AB|348.82|Brain death
C0006110|ICD9CM|PT|348.82|Brain death
C0006111|ICD9CM|PT|348.9|Unspecified condition of brain
C0006111|ICD9CM|AB|348.9|Brain condition NOS
C0006112|ICD9CM|AB|348.31|Metabolic encephalopathy
C0006112|ICD9CM|PT|348.31|Metabolic encephalopathy
C0006114|ICD9CM|AB|348.5|Cerebral edema
C0006114|ICD9CM|PT|348.5|Cerebral edema
C0006118|ICD9CM|AB|239.6|Brain neoplasm NOS
C0006118|ICD9CM|PT|239.6|Neoplasm of unspecified nature of brain
C0006123|ICD9CM|PT|362.32|Retinal arterial branch occlusion
C0006123|ICD9CM|AB|362.32|Arterial branch occlus
C0006131|ICD9CM|AB|744.42|Branchial cleft cyst
C0006131|ICD9CM|PT|744.42|Branchial cleft cyst
C0006145|ICD9CM|HT|610-612.99|DISORDERS OF BREAST
C0006145|ICD9CM|AB|611.9|Breast disorder NOS
C0006145|ICD9CM|PT|611.9|Unspecified breast disorder
C0006155|ICD9CM|PT|93.18|Breathing exercise
C0006155|ICD9CM|AB|93.18|Pt breathing exercise
C0006158|ICD9CM|HT|652.2|Breech presentation without mention of version
C0006181|ICD9CM|AB|081.1|Brill's disease
C0006181|ICD9CM|PT|081.1|Brill's disease
C0006267|ICD9CM|HT|494|Bronchiectasis
C0006277|ICD9CM|AB|490|Bronchitis NOS
C0006277|ICD9CM|PT|490|Bronchitis, not specified as acute or chronic
C0006285|ICD9CM|PT|485|Bronchopneumonia, organism unspecified
C0006285|ICD9CM|AB|485|Bronchopneumonia org NOS
C0006309|ICD9CM|HT|023|Brucellosis
C0006309|ICD9CM|AB|023.9|Brucellosis NOS
C0006309|ICD9CM|PT|023.9|Brucellosis, unspecified
C0006384|ICD9CM|AB|426.50|Bundle branch block NOS
C0006384|ICD9CM|PT|426.50|Bundle branch block, unspecified
C0006386|ICD9CM|AB|727.1|Bunion
C0006386|ICD9CM|PT|727.1|Bunion
C0006413|ICD9CM|HT|200.2|Burkitt's tumor or lymphoma
C0006420|ICD9CM|HT|947|Burn of internal organs
C0006420|ICD9CM|AB|947.9|Burn internal organ NOS
C0006420|ICD9CM|PT|947.9|Burn of internal organs, unspecified site
C0006421|ICD9CM|PT|941.02|Burn of unspecified degree of eye (with other parts of face, head, and neck)
C0006421|ICD9CM|AB|941.02|Burn NOS eye
C0006434|ICD9CM|HT|940-949.99|BURNS
C0006434|ICD9CM|AB|949.0|Burn NOS
C0006434|ICD9CM|PT|949.0|Burn of unspecified site, unspecified degree
C0006625|ICD9CM|AB|799.4|Cachexia
C0006625|ICD9CM|PT|799.4|Cachexia
C0006690|ICD9CM|PT|727.82|Calcium deposits in tendon and bursa
C0006690|ICD9CM|AB|727.82|Calcium deposit tendon
C0006705|ICD9CM|HT|275.4|Disorders of calcium metabolism
C0006705|ICD9CM|PT|275.40|Unspecified disorder of calcium metabolism
C0006705|ICD9CM|AB|275.40|Dis calcium metablsm NOS
C0006739|ICD9CM|HT|574.5|Calculus of bile duct without mention of cholecystitis
C0006741|ICD9CM|HT|574.2|Calculus of gallbladder without mention of cholecystitis
C0006742|ICD9CM|PT|574.20|Calculus of gallbladder without mention of cholecystitis, without mention of obstruction
C0006742|ICD9CM|AB|574.20|Cholelithiasis NOS
C0006759|ICD9CM|AB|E009.1|Calisthenics
C0006759|ICD9CM|PT|E009.1|Activity involving calisthenics
C0006826|ICD9CM|HT|199|Malignant neoplasm without specification of site
C0006840|ICD9CM|HT|112|Candidiasis
C0006840|ICD9CM|PT|112.9|Candidiasis of unspecified site
C0006840|ICD9CM|AB|112.9|Candidiasis site NOS
C0006842|ICD9CM|PT|112.3|Candidiasis of skin and nails
C0006842|ICD9CM|AB|112.3|Cutaneous candidiasis
C0006849|ICD9CM|PT|112.0|Candidiasis of mouth
C0006849|ICD9CM|AB|112.0|Thrush
C0006868|ICD9CM|HT|305.2|Cannabis abuse
C0006870|ICD9CM|HT|304.3|Cannabis dependence
C0006897|ICD9CM|AB|127.5|Capillariasis
C0006897|ICD9CM|PT|127.5|Capillariasis
C0007079|ICD9CM|PT|680.9|Carbuncle and furuncle of unspecified site
C0007079|ICD9CM|AB|680.9|Carbuncle NOS
C0007099|ICD9CM|HT|230-234.99|CARCINOMA IN SITU
C0007099|ICD9CM|PT|234.9|Carcinoma in situ, site unspecified
C0007099|ICD9CM|AB|234.9|Ca in situ NOS
C0007100|ICD9CM|PT|234.8|Carcinoma in situ of other specified sites
C0007100|ICD9CM|AB|234.8|Ca in situ NEC
C0007102|ICD9CM|HT|153|Malignant neoplasm of colon
C0007102|ICD9CM|PT|153.9|Malignant neoplasm of colon, unspecified site
C0007102|ICD9CM|AB|153.9|Malignant neo colon NOS
C0007107|ICD9CM|HT|161|Malignant neoplasm of larynx
C0007107|ICD9CM|PT|161.9|Malignant neoplasm of larynx, unspecified
C0007107|ICD9CM|AB|161.9|Malignant neo larynx NOS
C0007115|ICD9CM|PT|193|Malignant neoplasm of thyroid gland
C0007115|ICD9CM|AB|193|Malign neopl thyroid
C0007177|ICD9CM|PT|423.3|Cardiac tamponade
C0007177|ICD9CM|AB|423.3|Cardiac tamponade
C0007192|ICD9CM|AB|425.5|Alcoholic cardiomyopathy
C0007192|ICD9CM|PT|425.5|Alcoholic cardiomyopathy
C0007194|ICD9CM|HT|425.1|Hypertrophic cardiomyopathy
C0007203|ICD9CM|PT|99.60|Cardiopulmonary resuscitation, not otherwise specified
C0007203|ICD9CM|AB|99.60|Cardiopulm resuscita NOS
C0007222|ICD9CM|AB|429.2|Ascvd
C0007222|ICD9CM|PT|429.2|Cardiovascular disease, unspecified
C0007233|ICD9CM|PT|V57.0|Care involving breathing exercises
C0007233|ICD9CM|AB|V57.0|Breathing exercises
C0007234|ICD9CM|HT|V57.2|Care involving occupational therapy and vocational rehabilitation
C0007235|MTH|PN|NOCODE|Physical therapy NEC in ICD9CM_2014
C0007235|ICD9CM|PT|V57.1|Care involving other physical therapy
C0007235|ICD9CM|AB|V57.1|Physical therapy NEC
C0007237|ICD9CM|PT|V57.9|Care involving unspecified rehabilitation procedure
C0007237|ICD9CM|HT|V57|Care involving use of rehabilitation procedures
C0007237|ICD9CM|AB|V57.9|Rehabilitation proc NOS
C0007286|ICD9CM|AB|354.0|Carpal tunnel syndrome
C0007286|ICD9CM|PT|354.0|Carpal tunnel syndrome
C0007294|ICD9CM|AB|V18.9|Fam hx genet dis carrier
C0007294|ICD9CM|PT|V18.9|Family history of genetic disease carrier
C0007347|ICD9CM|HT|62.4|Bilateral orchiectomy
C0007361|ICD9CM|AB|078.3|Cat-scratch disease
C0007361|ICD9CM|PT|078.3|Cat-scratch disease
C0007431|ICD9CM|AB|38.91|Arterial catheterization
C0007431|ICD9CM|PT|38.91|Arterial catheterization
C0007459|ICD9CM|PT|344.61|Cauda equina syndrome with neurogenic bladder
C0007459|ICD9CM|AB|344.61|Neurogenic bladder
C0007570|ICD9CM|AB|579.0|Celiac disease
C0007570|ICD9CM|PT|579.0|Celiac disease
C0007643|ICD9CM|PT|528.3|Cellulitis and abscess of oral soft tissues
C0007643|ICD9CM|AB|528.3|Cellulitis/abscess mouth
C0007644|ICD9CM|PT|681.9|Cellulitis and abscess of unspecified digit
C0007644|ICD9CM|AB|681.9|Cellulitis of digit NOS
C0007645|ICD9CM|AB|682.9|Cellulitis NOS
C0007645|ICD9CM|PT|682.9|Cellulitis and abscess of unspecified sites
C0007686|ICD9CM|PT|371.03|Central opacity of cornea
C0007686|ICD9CM|AB|371.03|Central opacity, cornea
C0007688|ICD9CM|PT|362.31|Central retinal artery occlusion
C0007688|ICD9CM|AB|362.31|Cent retina artery occlu
C0007767|ICD9CM|PT|88.41|Arteriography of cerebral arteries
C0007767|ICD9CM|AB|88.41|Contr cerebr arteriogram
C0007773|ICD9CM|AB|437.4|Cerebral arteritis
C0007773|ICD9CM|PT|437.4|Cerebral arteritis
C0007775|ICD9CM|AB|437.0|Cerebral atherosclerosis
C0007775|ICD9CM|PT|437.0|Cerebral atherosclerosis
C0007780|ICD9CM|HT|434.1|Cerebral embolism
C0007788|ICD9CM|AB|330.1|Cerebral lipidoses
C0007788|ICD9CM|PT|330.1|Cerebral lipidoses
C0007795|ICD9CM|AB|341.1|Schilder's disease
C0007795|ICD9CM|PT|341.1|Schilder's disease
C0007814|ICD9CM|PT|388.61|Cerebrospinal fluid otorrhea
C0007814|ICD9CM|AB|388.61|Cerebrosp fluid otorrhea
C0007815|ICD9CM|PT|349.81|Cerebrospinal fluid rhinorrhea
C0007815|ICD9CM|AB|349.81|Cerebrospinal rhinorrhea
C0007820|ICD9CM|PT|437.9|Unspecified cerebrovascular disease
C0007820|ICD9CM|HT|430-438.99|CEREBROVASCULAR DISEASE
C0007820|ICD9CM|AB|437.9|Cerebrovasc disease NOS
C0007832|ICD9CM|HT|364.2|Certain types of iridocyclitis
C0007847|ICD9CM|HT|180|Malignant neoplasm of cervix uteri
C0007847|ICD9CM|PT|180.9|Malignant neoplasm of cervix uteri, unspecified site
C0007847|ICD9CM|AB|180.9|Mal neo cervix uteri NOS
C0007859|ICD9CM|AB|723.1|Cervicalgia
C0007859|ICD9CM|PT|723.1|Cervicalgia
C0007861|ICD9CM|AB|616.0|Cervicitis
C0007861|ICD9CM|PT|616.0|Cervicitis and endocervicitis
C0007868|ICD9CM|AB|622.10|Dysplasia of cervix NOS
C0007868|ICD9CM|HT|622.1|Dysplasia of cervix (uteri)
C0007868|ICD9CM|PT|622.10|Dysplasia of cervix, unspecified
C0007871|ICD9CM|AB|622.5|Incompetence of cervix
C0007871|ICD9CM|PT|622.5|Incompetence of cervix
C0007876|ICD9CM|HT|74.9|Cesarean section of unspecified type
C0007876|ICD9CM|HT|74|Cesarean section and removal of fetus
C0007878|ICD9CM|PT|74.4|Cesarean section of other specified type
C0007878|ICD9CM|AB|74.4|Cesarean section NEC
C0007894|ICD9CM|AB|123.9|Cestode infection NOS
C0007894|ICD9CM|PT|123.9|Cestode infection, unspecified
C0007930|ICD9CM|PT|086.0|Chagas' disease with heart involvement
C0007930|ICD9CM|AB|086.0|Chagas disease of heart
C0007932|ICD9CM|PT|086.2|Chagas' disease without mention of organ involvement
C0007932|ICD9CM|AB|086.2|Chagas disease NOS
C0007933|ICD9CM|AB|373.2|Chalazion
C0007933|ICD9CM|PT|373.2|Chalazion
C0007947|ICD9CM|AB|099.0|Chancroid
C0007947|ICD9CM|PT|099.0|Chancroid
C0007953|ICD9CM|AB|94.03|Character analysis
C0007953|ICD9CM|PT|94.03|Character analysis
C0007959|ICD9CM|PT|356.1|Peroneal muscular atrophy
C0007959|ICD9CM|AB|356.1|Peroneal muscle atrophy
C0008031|ICD9CM|HT|786.5|Chest pain
C0008031|ICD9CM|AB|786.50|Chest pain NOS
C0008031|ICD9CM|PT|786.50|Chest pain, unspecified
C0008039|ICD9CM|PT|786.04|Cheyne-Stokes respiration
C0008039|ICD9CM|AB|786.04|Cheyne-stokes respiratn
C0008049|ICD9CM|HT|052|Chickenpox
C0008058|ICD9CM|AB|991.5|Chilblains
C0008058|ICD9CM|PT|991.5|Chilblains
C0008060|ICD9CM|AB|995.50|Child abuse NOS
C0008060|ICD9CM|HT|995.5|Child maltreatment syndrome
C0008060|ICD9CM|PT|995.50|Child abuse, unspecified
C0008062|ICD9CM|AB|995.53|Child sexual abuse
C0008062|ICD9CM|PT|995.53|Child sexual abuse
C0008297|ICD9CM|AB|748.0|Choanal atresia
C0008297|ICD9CM|PT|748.0|Choanal atresia
C0008310|ICD9CM|PT|51.10|Endoscopic retrograde cholangiopancreatography [ERCP]
C0008310|ICD9CM|AB|51.10|Endosc retro cholangiopa
C0008311|ICD9CM|AB|576.1|Cholangitis
C0008311|ICD9CM|PT|576.1|Cholangitis
C0008320|ICD9CM|AB|51.22|Cholecystectomy
C0008320|ICD9CM|HT|51.2|Cholecystectomy
C0008320|ICD9CM|PT|51.22|Cholecystectomy
C0008325|ICD9CM|AB|575.10|Cholecystitis NOS
C0008325|ICD9CM|PT|575.10|Cholecystitis, unspecified
C0008338|ICD9CM|PT|51.91|Repair of laceration of gallbladder
C0008338|ICD9CM|AB|51.91|Repair gb laceration
C0008350|ICD9CM|HT|574|Cholelithiasis
C0008354|ICD9CM|HT|001|Cholera
C0008354|ICD9CM|AB|001.9|Cholera NOS
C0008354|ICD9CM|PT|001.0|Cholera due to vibrio cholerae
C0008354|ICD9CM|PT|001.9|Cholera, unspecified
C0008354|ICD9CM|AB|001.0|Cholera d/t vib cholerae
C0008370|ICD9CM|AB|576.2|Obstruction of bile duct
C0008370|ICD9CM|PT|576.2|Obstruction of bile duct
C0008373|ICD9CM|AB|385.30|Cholesteatoma NOS
C0008373|ICD9CM|PT|385.30|Cholesteatoma, unspecified
C0008374|ICD9CM|HT|385.3|Cholesteatoma of middle ear and mastoid
C0008374|ICD9CM|PT|385.33|Cholesteatoma of middle ear and mastoid
C0008374|ICD9CM|AB|385.33|Cholestma mid ear/mstoid
C0008449|ICD9CM|AB|756.4|Chondrodystrophy
C0008449|ICD9CM|PT|756.4|Chondrodystrophy
C0008475|ICD9CM|AB|717.7|Chondromalacia patellae
C0008475|ICD9CM|PT|717.7|Chondromalacia of patella
C0008511|ICD9CM|HT|363|Chorioretinal inflammations, scars, and other disorders of choroid
C0008512|ICD9CM|HT|363.3|Chorioretinal scars
C0008512|ICD9CM|AB|363.30|Chorioretinal scar NOS
C0008512|ICD9CM|PT|363.30|Chorioretinal scar, unspecified
C0008513|ICD9CM|AB|363.20|Chorioretinitis NOS
C0008513|ICD9CM|PT|363.20|Chorioretinitis, unspecified
C0008521|ICD9CM|PT|363.9|Unspecified disorder of choroid
C0008521|ICD9CM|AB|363.9|Choroidal disorder NOS
C0008522|ICD9CM|PT|363.61|Choroidal hemorrhage, unspecified
C0008522|ICD9CM|AB|363.61|Choroidal hemorrhage NOS
C0008525|ICD9CM|AB|363.55|Choroideremia
C0008525|ICD9CM|PT|363.55|Choroideremia
C0008533|ICD9CM|PT|286.1|Congenital factor IX disorder
C0008533|ICD9CM|AB|286.1|Cong factor IX disorder
C0008582|ICD9CM|AB|117.2|Chromoblastomycosis
C0008582|ICD9CM|PT|117.2|Chromoblastomycosis
C0008626|ICD9CM|PT|758.9|Conditions due to anomaly of unspecified chromosome
C0008626|ICD9CM|HT|758|Chromosomal anomalies
C0008626|ICD9CM|AB|758.9|Chromosome anomaly NOS
C0008677|ICD9CM|HT|491|Chronic bronchitis
C0008677|ICD9CM|AB|491.9|Chronic bronchitis NOS
C0008677|ICD9CM|PT|491.9|Unspecified chronic bronchitis
C0008681|ICD9CM|PT|473.2|Chronic ethmoidal sinusitis
C0008681|ICD9CM|AB|473.2|Chr ethmoidal sinusitis
C0008682|ICD9CM|PT|301.51|Chronic factitious illness with physical symptoms
C0008682|ICD9CM|AB|301.51|Chr factitious illness
C0008683|ICD9CM|PT|473.1|Chronic frontal sinusitis
C0008683|ICD9CM|AB|473.1|Chr frontal sinusitis
C0008684|ICD9CM|HT|523.1|Chronic gingivitis
C0008685|ICD9CM|PT|582.2|Chronic glomerulonephritis with lesion of membranoproliferative glomerulonephritis
C0008685|ICD9CM|AB|582.2|Chr membranoprolif nephr
C0008686|ICD9CM|PT|582.1|Chronic glomerulonephritis with lesion of membranous glomerulonephritis
C0008686|ICD9CM|AB|582.1|Chr membranous nephritis
C0008698|ICD9CM|PT|473.0|Chronic maxillary sinusitis
C0008698|ICD9CM|AB|473.0|Chr maxillary sinusitis
C0008701|ICD9CM|PT|307.22|Chronic motor or vocal tic disorder
C0008701|ICD9CM|AB|307.22|Chr motor/vocal tic dis
C0008707|ICD9CM|HT|730.1|Chronic osteomyelitis
C0008707|ICD9CM|PT|730.10|Chronic osteomyelitis, site unspecified
C0008707|ICD9CM|AB|730.10|Chr osteomyelitis-unsp
C0008711|ICD9CM|AB|472.0|Chronic rhinitis
C0008711|ICD9CM|PT|472.0|Chronic rhinitis
C0008712|ICD9CM|PT|473.3|Chronic sphenoidal sinusitis
C0008712|ICD9CM|AB|473.3|Chr sphenoidal sinusitis
C0008819|ICD9CM|AB|64.0|Circumcision
C0008819|ICD9CM|PT|64.0|Circumcision
C0008827|ICD9CM|PT|571.5|Cirrhosis of liver without mention of alcohol
C0008827|ICD9CM|AB|571.5|Cirrhosis of liver NOS
C0008924|ICD9CM|HT|749.1|Cleft lip
C0008924|ICD9CM|AB|749.10|Cleft lip NOS
C0008924|ICD9CM|PT|749.10|Cleft lip, unspecified
C0008925|ICD9CM|HT|749.0|Cleft palate
C0008925|ICD9CM|AB|749.00|Cleft palate NOS
C0008925|ICD9CM|PT|749.00|Cleft palate, unspecified
C0009021|ICD9CM|AB|121.1|Clonorchiasis
C0009021|ICD9CM|PT|121.1|Clonorchiasis
C0009039|ICD9CM|PT|99.63|Closed chest cardiac massage
C0009039|ICD9CM|AB|99.63|Closed chest card massag
C0009041|ICD9CM|HT|835.0|Closed dislocation of hip
C0009043|ICD9CM|PT|839.8|Closed dislocation, multiple and ill-defined sites
C0009043|ICD9CM|AB|839.8|Dislocation NEC-closed
C0009044|ICD9CM|HT|814.0|Closed fractures of carpal bones
C0009044|ICD9CM|PT|814.00|Closed fracture of carpal bone, unspecified
C0009044|ICD9CM|AB|814.00|Fx carpal bone NOS-close
C0009045|ICD9CM|PT|802.4|Closed fracture of malar and maxillary bones
C0009045|ICD9CM|AB|802.4|Fx malar/maxillary-close
C0009048|ICD9CM|PT|805.8|Closed fracture of unspecified vertebral column without mention of spinal cord injury
C0009048|ICD9CM|AB|805.8|Vertebral fx NOS-closed
C0009080|ICD9CM|AB|781.5|Clubbing of fingers
C0009080|ICD9CM|PT|781.5|Clubbing of fingers
C0009081|ICD9CM|AB|754.51|Talipes equinovarus
C0009081|ICD9CM|PT|754.51|Talipes equinovarus
C0009088|ICD9CM|PT|339.02|Chronic cluster headache
C0009088|ICD9CM|AB|339.02|Chronic cluster headache
C0009088|ICD9CM|PT|339.00|Cluster headache syndrome, unspecified
C0009088|ICD9CM|AB|339.00|Cluster headache syn NOS
C0009171|ICD9CM|HT|305.6|Cocaine abuse
C0009171|ICD9CM|PT|305.60|Cocaine abuse, unspecified
C0009171|ICD9CM|AB|305.60|Cocaine abuse-unspec
C0009186|ICD9CM|HT|114|Coccidioidomycosis
C0009186|ICD9CM|AB|114.9|Coccidioidomycosis NOS
C0009186|ICD9CM|PT|114.9|Coccidioidomycosis, unspecified
C0009324|ICD9CM|HT|556|Ulcerative colitis
C0009324|ICD9CM|PT|556.9|Ulcerative colitis, unspecified
C0009324|ICD9CM|AB|556.9|Ulceratve colitis unspcf
C0009354|ICD9CM|PT|813.41|Closed Colles' fracture
C0009354|ICD9CM|AB|813.41|Colles' fracture-closed
C0009378|ICD9CM|AB|45.23|Colonoscopy
C0009378|ICD9CM|PT|45.23|Colonoscopy
C0009410|ICD9CM|HT|46.1|Colostomy
C0009410|ICD9CM|AB|46.10|Colostomy NOS
C0009410|ICD9CM|PT|46.10|Colostomy, not otherwise specified
C0009421|ICD9CM|AB|780.01|Coma
C0009421|ICD9CM|PT|780.01|Coma
C0009443|ICD9CM|AB|460|Acute nasopharyngitis
C0009443|ICD9CM|PT|460|Acute nasopharyngitis [common cold]
C0009447|ICD9CM|PT|279.06|Common variable immunodeficiency
C0009447|ICD9CM|AB|279.06|Common variabl immunodef
C0009451|ICD9CM|PT|331.3|Communicating hydrocephalus
C0009451|ICD9CM|AB|331.3|Communicat hydrocephalus
C0009492|ICD9CM|AB|958.90|Compartment syndrome NOS
C0009492|ICD9CM|PT|958.90|Compartment syndrome, unspecified
C0009557|ICD9CM|AB|25.3|Complete glossectomy
C0009557|ICD9CM|PT|25.3|Complete glossectomy
C0009568|ICD9CM|HT|996.8|Complications of transplanted organ
C0009592|ICD9CM|AB|348.4|Compression of brain
C0009592|ICD9CM|PT|348.4|Compression of brain
C0009595|ICD9CM|PT|301.4|Obsessive-compulsive personality disorder
C0009595|ICD9CM|AB|301.4|Obsessive-compulsive dis
C0009663|ICD9CM|AB|078.11|Condyloma acuminatum
C0009663|ICD9CM|PT|078.11|Condyloma acuminatum
C0009677|ICD9CM|AB|750.15|Cong macroglossia
C0009677|ICD9CM|PT|750.15|Macroglossia
C0009680|ICD9CM|HT|756.7|Anomalies of abdominal wall, congenital
C0009680|ICD9CM|PT|756.70|Anomaly of abdominal wall, unspecified
C0009680|ICD9CM|AB|756.70|Congn anoml abd wall NOS
C0009681|ICD9CM|HT|747.3|Anomalies of pulmonary artery, congenital
C0009691|ICD9CM|AB|743.30|Congenital cataract NOS
C0009691|ICD9CM|PT|743.30|Congenital cataract, unspecified
C0009699|ICD9CM|PT|286.3|Congenital deficiency of other clotting factors
C0009699|ICD9CM|AB|286.3|Cong def clot factor NEC
C0009702|ICD9CM|PT|754.30|Congenital dislocation of hip, unilateral
C0009702|ICD9CM|AB|754.30|Cong hip disloc, unilat
C0009726|ICD9CM|PT|757.33|Congenital pigmentary anomalies of skin
C0009726|ICD9CM|AB|757.33|Cong skin pigment anomal
C0009733|ICD9CM|PT|750.3|Tracheoesophageal fistula, esophageal atresia and stenosis
C0009733|ICD9CM|AB|750.3|Cong esoph fistula/atres
C0009759|ICD9CM|PT|372.9|Unspecified disorder of conjunctiva
C0009759|ICD9CM|HT|372|Disorders of conjunctiva
C0009759|ICD9CM|AB|372.9|Conjunctiva disorder NOS
C0009760|ICD9CM|AB|372.72|Conjunctival hemorrhage
C0009760|ICD9CM|PT|372.72|Conjunctival hemorrhage
C0009763|ICD9CM|AB|372.30|Conjunctivitis NOS
C0009763|ICD9CM|PT|372.30|Conjunctivitis, unspecified
C0009765|ICD9CM|PT|077.4|Epidemic hemorrhagic conjunctivitis
C0009765|ICD9CM|AB|077.4|Epidem hem conjunctivit
C0009770|ICD9CM|AB|077.0|Inclusion conjunctivitis
C0009770|ICD9CM|PT|077.0|Inclusion conjunctivitis
C0009773|ICD9CM|AB|372.13|Vernal conjunctivitis
C0009773|ICD9CM|PT|372.13|Vernal conjunctivitis
C0009806|ICD9CM|HT|564.0|Constipation
C0009806|ICD9CM|AB|564.00|Constipation NOS
C0009806|ICD9CM|PT|564.00|Constipation, unspecified
C0009818|ICD9CM|AB|89.09|Consultation NOS
C0009818|ICD9CM|PT|89.09|Consultation, not otherwise specified
C0009833|ICD9CM|HT|692|Contact dermatitis and other eczema
C0009834|ICD9CM|HT|692.8|Contact dermatitis and other eczema due to other specified agents
C0009834|ICD9CM|PT|692.89|Contact dermatitis and other eczema due to other specified agents
C0009834|ICD9CM|AB|692.89|Dermatitis NEC
C0009918|ICD9CM|HT|718.4|Contracture of joint
C0009918|ICD9CM|PT|718.40|Contracture of joint, site unspecified
C0009918|ICD9CM|AB|718.40|Jt contracture-unspec
C0009926|ICD9CM|AB|87.66|Contrast pancreatogram
C0009926|ICD9CM|PT|87.66|Contrast pancreatogram
C0009938|ICD9CM|AB|924.9|Contusion NOS
C0009938|ICD9CM|PT|924.9|Contusion of unspecified site
C0009941|ICD9CM|PT|V66.5|Convalescence following other treatment
C0009941|ICD9CM|AB|V66.5|Convalescence NEC
C0009946|ICD9CM|AB|300.11|Conversion disorder
C0009946|ICD9CM|PT|300.11|Conversion disorder
C0009952|ICD9CM|AB|780.31|Febrile convulsions NOS
C0009952|ICD9CM|PT|780.31|Febrile convulsions (simple), unspecified
C0009995|ICD9CM|AB|746.82|Cor triatriatum
C0009995|ICD9CM|PT|746.82|Cor triatriatum
C0010009|ICD9CM|HT|03.2|Chordotomy
C0010034|ICD9CM|PT|371.9|Unspecified corneal disorder
C0010034|ICD9CM|AB|371.9|Corneal disorder NOS
C0010035|ICD9CM|HT|371.5|Hereditary corneal dystrophies
C0010035|ICD9CM|AB|371.50|Corneal dystrophy NOS
C0010035|ICD9CM|PT|371.50|Hereditary corneal dystrophy, unspecified
C0010037|ICD9CM|HT|371.2|Corneal edema
C0010037|ICD9CM|AB|371.20|Corneal edema NOS
C0010037|ICD9CM|PT|371.20|Corneal edema, unspecified
C0010038|ICD9CM|AB|371.00|Corneal opacity NOS
C0010038|ICD9CM|PT|371.00|Corneal opacity, unspecified
C0010042|ICD9CM|HT|11.6|Corneal transplant
C0010042|ICD9CM|AB|11.60|Corneal transplant NOS
C0010042|ICD9CM|PT|11.60|Corneal transplant, not otherwise specified
C0010043|ICD9CM|HT|370.0|Corneal ulcer
C0010043|ICD9CM|AB|370.00|Corneal ulcer NOS
C0010043|ICD9CM|PT|370.00|Corneal ulcer, unspecified
C0010051|ICD9CM|PT|414.11|Aneurysm of coronary vessels
C0010051|ICD9CM|AB|414.11|Aneurysm coronary vessel
C0010054|ICD9CM|HT|414.0|Coronary atherosclerosis
C0010055|ICD9CM|AB|36.10|Aortocoronary bypass NOS
C0010055|ICD9CM|HT|36.1|Bypass anastomosis for heart revascularization
C0010055|ICD9CM|PT|36.10|Aortocoronary bypass for heart revascularization, not otherwise specified
C0010200|ICD9CM|AB|786.2|Cough
C0010200|ICD9CM|PT|786.2|Cough
C0010232|ICD9CM|PT|051.01|Cowpox
C0010232|ICD9CM|AB|051.01|Cowpox
C0010244|ICD9CM|PT|079.2|Coxsackie virus infection in conditions classified elsewhere and of unspecified site
C0010244|ICD9CM|AB|079.2|Coxsackie virus inf NOS
C0010261|ICD9CM|PT|521.81|Cracked tooth
C0010261|ICD9CM|AB|521.81|Cracked tooth
C0010263|ICD9CM|PT|729.82|Cramp of limb
C0010263|ICD9CM|AB|729.82|Cramp in limb
C0010266|ICD9CM|PT|352.9|Unspecified disorder of cranial nerves
C0010266|ICD9CM|AB|352.9|Cranial nerve dis NOS
C0010308|ICD9CM|PT|243|Congenital hypothyroidism
C0010308|ICD9CM|AB|243|Congenital hypothyroidsm
C0010314|ICD9CM|AB|758.31|Cri-du-chat syndrome
C0010314|ICD9CM|PT|758.31|Cri-du-chat syndrome
C0010332|ICD9CM|AB|94.35|Crisis intervention
C0010332|ICD9CM|PT|94.35|Crisis intervention
C0010380|ICD9CM|AB|464.4|Croup
C0010380|ICD9CM|PT|464.4|Croup
C0010414|ICD9CM|AB|117.5|Cryptococcosis
C0010414|ICD9CM|PT|117.5|Cryptococcosis
C0010417|ICD9CM|AB|752.51|Undescended testis
C0010417|ICD9CM|PT|752.51|Undescended testis
C0010418|ICD9CM|AB|007.4|Cryptosporidiosis
C0010418|ICD9CM|PT|007.4|Cryptosporidiosis
C0010443|ICD9CM|AB|70.22|Culdoscopy
C0010443|ICD9CM|PT|70.22|Culdoscopy
C0010481|ICD9CM|AB|255.0|Cushing's syndrome
C0010481|ICD9CM|PT|255.0|Cushing's syndrome
C0010487|ICD9CM|PT|031.1|Cutaneous diseases due to other mycobacteria
C0010487|ICD9CM|AB|031.1|Cutaneous mycobacteria
C0010520|ICD9CM|AB|782.5|Cyanosis
C0010520|ICD9CM|PT|782.5|Cyanosis
C0010598|ICD9CM|AB|301.13|Cyclothymic disorder
C0010598|ICD9CM|PT|301.13|Cyclothymic disorder
C0010598|ICD9CM|HT|301.1|Affective personality disorder
C0010598|ICD9CM|PT|301.10|Affective personality disorder, unspecified
C0010598|ICD9CM|AB|301.10|Affectiv personality NOS
C0010623|ICD9CM|PT|577.2|Cyst and pseudocyst of pancreas
C0010623|ICD9CM|AB|577.2|Pancreat cyst/pseudocyst
C0010674|ICD9CM|HT|277.0|Cystic fibrosis
C0010676|ICD9CM|PT|277.00|Cystic fibrosis without mention of meconium ileus
C0010676|ICD9CM|AB|277.00|Cystic fibros w/o ileus
C0010678|ICD9CM|AB|123.1|Cysticercosis
C0010678|ICD9CM|PT|123.1|Cysticercosis
C0010692|ICD9CM|HT|595|Cystitis
C0010692|ICD9CM|AB|595.9|Cystitis NOS
C0010692|ICD9CM|PT|595.9|Cystitis, unspecified
C0010700|ICD9CM|PT|57.81|Suture of laceration of bladder
C0010700|ICD9CM|AB|57.81|Suture bladder lacerat
C0010705|ICD9CM|AB|57.21|Vesicostomy
C0010705|ICD9CM|HT|57.2|Vesicostomy
C0010705|ICD9CM|PT|57.21|Vesicostomy
C0010823|ICD9CM|AB|078.5|Cytomegaloviral disease
C0010823|ICD9CM|PT|078.5|Cytomegaloviral disease
C0010930|ICD9CM|AB|375.30|Dacryocystitis NOS
C0010930|ICD9CM|PT|375.30|Dacryocystitis, unspecified
C0010931|ICD9CM|AB|09.81|Dacryocystorhinostomy
C0010931|ICD9CM|PT|09.81|Dacryocystorhinostomy [DCR]
C0010932|ICD9CM|PT|09.53|Incision of lacrimal sac
C0010932|ICD9CM|AB|09.53|Lacrimal sac incision
C0010963|ICD9CM|AB|E005.0|Dancing
C0010963|ICD9CM|PT|E005.0|Activities involving dancing
C0011057|ICD9CM|AB|388.2|Sudden hearing loss NOS
C0011057|ICD9CM|PT|388.2|Sudden hearing loss, unspecified
C0011119|ICD9CM|AB|993.3|Caisson disease
C0011119|ICD9CM|PT|993.3|Caisson disease
C0011124|ICD9CM|AB|799.81|Decreased libido
C0011124|ICD9CM|PT|799.81|Decreased libido
C0011127|ICD9CM|HT|707.0|Pressure ulcer
C0011127|ICD9CM|AB|707.00|Pressure ulcer, site NOS
C0011127|ICD9CM|PT|707.00|Pressure ulcer, unspecified site
C0011157|ICD9CM|PT|269.1|Deficiency of other vitamins
C0011157|ICD9CM|AB|269.1|Vitamin Deficiency NEC
C0011168|ICD9CM|HT|787.2|Dysphagia
C0011168|ICD9CM|AB|787.20|Dysphagia NOS
C0011168|ICD9CM|PT|787.20|Dysphagia, unspecified
C0011175|ICD9CM|AB|276.51|Dehydration
C0011175|ICD9CM|PT|276.51|Dehydration
C0011251|ICD9CM|AB|297.1|Delusional disorder
C0011251|ICD9CM|PT|297.1|Delusional disorder
C0011265|ICD9CM|HT|290.1|Presenile dementia
C0011269|ICD9CM|HT|290.4|Vascular dementia
C0011302|ICD9CM|PT|341.9|Demyelinating disease of central nervous system, unspecified
C0011302|ICD9CM|AB|341.9|Cns demyelination NOS
C0011311|ICD9CM|AB|061|Dengue
C0011311|ICD9CM|PT|061|Dengue
C0011334|ICD9CM|HT|521.0|Dental caries
C0011334|ICD9CM|AB|521.00|Dental caries NOS
C0011334|ICD9CM|PT|521.00|Dental caries, unspecified
C0011346|ICD9CM|AB|523.6|Accretions on teeth
C0011346|ICD9CM|PT|523.6|Accretions on teeth
C0011407|ICD9CM|AB|522.1|Necrosis of tooth pulp
C0011407|ICD9CM|PT|522.1|Necrosis of the pulp
C0011417|ICD9CM|PT|96.54|Dental scaling, polishing, and debridement
C0011417|ICD9CM|AB|96.54|Dental scaling & debride
C0011548|ICD9CM|PT|301.6|Dependent personality disorder
C0011548|ICD9CM|AB|301.6|Dependent personality
C0011593|ICD9CM|AB|86.25|Dermabrasion
C0011593|ICD9CM|PT|86.25|Dermabrasion
C0011604|ICD9CM|PT|693.0|Dermatitis due to drugs and medicines taken internally
C0011604|ICD9CM|AB|693.0|Drug dermatitis NOS
C0011608|ICD9CM|AB|694.0|Dermatitis herpetiformis
C0011608|ICD9CM|PT|694.0|Dermatitis herpetiformis
C0011630|ICD9CM|AB|111.9|Dermatomycosis NOS
C0011630|ICD9CM|HT|111|Dermatomycosis, other and unspecified
C0011630|ICD9CM|PT|111.9|Dermatomycosis, unspecified
C0011633|ICD9CM|AB|710.3|Dermatomyositis
C0011633|ICD9CM|PT|710.3|Dermatomyositis
C0011636|ICD9CM|HT|110|Dermatophytosis
C0011636|ICD9CM|PT|110.9|Dermatophytosis of unspecified site
C0011636|ICD9CM|AB|110.9|Dermatophytosis site NOS
C0011638|ICD9CM|PT|110.3|Dermatophytosis of groin and perianal area
C0011638|ICD9CM|AB|110.3|Dermatophytosis of groin
C0011640|ICD9CM|PT|110.0|Dermatophytosis of scalp and beard
C0011640|ICD9CM|AB|110.0|Dermatophyt scalp/beard
C0011757|ICD9CM|PT|315.4|Developmental coordination disorder
C0011757|ICD9CM|AB|315.4|Devel coordination dis
C0011848|ICD9CM|AB|253.5|Diabetes insipidus
C0011848|ICD9CM|PT|253.5|Diabetes insipidus
C0011849|ICD9CM|HT|250|Diabetes mellitus
C0011870|ICD9CM|HT|250.3|Diabetes with other coma
C0011871|ICD9CM|HT|250.7|Diabetes with peripheral circulatory disorders
C0011876|ICD9CM|AB|366.41|Diabetic cataract
C0011876|ICD9CM|PT|366.41|Diabetic cataract
C0011880|ICD9CM|HT|250.1|Diabetes with ketoacidosis
C0011881|ICD9CM|HT|250.4|Diabetes with renal manifestations
C0011882|ICD9CM|HT|250.6|Diabetes with neurological manifestations
C0011884|ICD9CM|HT|362.0|Diabetic retinopathy
C0011923|ICD9CM|AB|88.90|Diagnostic imaging NOS
C0011923|ICD9CM|PT|88.90|Diagnostic imaging, not elsewhere classified
C0011931|ICD9CM|PT|88.71|Diagnostic ultrasound of head and neck
C0011931|ICD9CM|AB|88.71|Dx ultrasound-head/neck
C0011974|ICD9CM|AB|691.0|Diaper or napkin rash
C0011974|ICD9CM|PT|691.0|Diaper or napkin rash
C0011991|ICD9CM|AB|787.91|Diarrhea
C0011991|ICD9CM|PT|787.91|Diarrhea
C0011999|ICD9CM|AB|742.51|Diastematomyelia
C0011999|ICD9CM|PT|742.51|Diastematomyelia
C0012002|ICD9CM|AB|93.34|Diathermy
C0012002|ICD9CM|PT|93.34|Diathermy
C0012236|ICD9CM|AB|279.11|Digeorge's syndrome
C0012236|ICD9CM|PT|279.11|Digeorge's syndrome
C0012242|ICD9CM|HT|520-579.99|DISEASES OF THE DIGESTIVE SYSTEM
C0012243|ICD9CM|PT|239.0|Neoplasm of unspecified nature of digestive system
C0012243|ICD9CM|AB|239.0|Digestive neoplasm NOS
C0012246|ICD9CM|PT|619.1|Digestive-genital tract fistula, female
C0012246|ICD9CM|AB|619.1|Digest-genit fistul, fem
C0012358|ICD9CM|HT|69.0|Dilation and curettage of uterus
C0012517|ICD9CM|AB|125.4|Dipetalonemiasis
C0012517|ICD9CM|PT|125.4|Dipetalonemiasis
C0012546|ICD9CM|HT|032|Diphtheria
C0012546|ICD9CM|AB|032.9|Diphtheria NOS
C0012546|ICD9CM|PT|032.9|Diphtheria, unspecified
C0012553|ICD9CM|PT|032.2|Anterior nasal diphtheria
C0012553|ICD9CM|AB|032.2|Ant nasal diphtheria
C0012554|ICD9CM|AB|032.81|Conjunctival diphtheria
C0012554|ICD9CM|PT|032.81|Conjunctival diphtheria
C0012555|ICD9CM|AB|032.85|Cutaneous diphtheria
C0012555|ICD9CM|PT|032.85|Cutaneous diphtheria
C0012556|ICD9CM|AB|032.0|Faucial diphtheria
C0012556|ICD9CM|PT|032.0|Faucial diphtheria
C0012557|ICD9CM|AB|032.3|Laryngeal diphtheria
C0012557|ICD9CM|PT|032.3|Laryngeal diphtheria
C0012558|ICD9CM|PT|032.1|Nasopharyngeal diphtheria
C0012558|ICD9CM|AB|032.1|Nasopharynx diphtheria
C0012561|ICD9CM|PT|123.4|Diphyllobothriasis, intestinal
C0012561|ICD9CM|AB|123.4|Diphyllobothrias intest
C0012569|ICD9CM|AB|368.2|Diplopia
C0012569|ICD9CM|PT|368.2|Diplopia
C0012691|ICD9CM|HT|830-839.99|DISLOCATION
C0012711|ICD9CM|PT|277.4|Disorders of bilirubin excretion
C0012711|ICD9CM|AB|277.4|Dis bilirubin excretion
C0012714|ICD9CM|PT|275.1|Disorders of copper metabolism
C0012714|ICD9CM|AB|275.1|Dis copper metabolism
C0012715|ICD9CM|HT|275.0|Disorders of iron metabolism
C0012716|ICD9CM|PT|275.2|Disorders of magnesium metabolism
C0012716|ICD9CM|AB|275.2|Dis magnesium metabolism
C0012736|ICD9CM|HT|441.0|Dissecting aneurysm of aorta
C0012736|ICD9CM|HT|441|Aortic aneurysm and dissection
C0012739|ICD9CM|AB|286.6|Defibrination syndrome
C0012739|ICD9CM|PT|286.6|Defibrination syndrome
C0012746|ICD9CM|AB|300.15|Dissociative react NOS
C0012746|ICD9CM|PT|300.15|Dissociative disorder or reaction, unspecified
C0012765|ICD9CM|PT|527.7|Disturbance of salivary secretion
C0012765|ICD9CM|AB|527.7|Salivary secretion dis
C0012766|ICD9CM|PT|782.0|Disturbance of skin sensation
C0012766|ICD9CM|AB|782.0|Skin sensation disturb
C0012767|ICD9CM|PT|520.6|Disturbances in tooth eruption
C0012767|ICD9CM|AB|520.6|Tooth eruption disturb
C0012811|ICD9CM|HT|562.1|Diverticula of colon
C0012827|ICD9CM|PT|04.03|Division or crushing of other cranial and peripheral nerves
C0012827|ICD9CM|AB|04.03|Periph nerve div NEC
C0013019|ICD9CM|PT|V59.9|Donors of unspecified organ or tissue
C0013019|ICD9CM|AB|V59.9|Org or tissue donor NOS
C0013069|ICD9CM|PT|745.11|Double outlet right ventricle
C0013069|ICD9CM|AB|745.11|Double outlet rt ventric
C0013080|ICD9CM|AB|758.0|Down's syndrome
C0013080|ICD9CM|PT|758.0|Down's syndrome
C0013100|ICD9CM|AB|125.7|Dracontiasis
C0013100|ICD9CM|PT|125.7|Dracontiasis
C0013143|ICD9CM|PT|994.1|Drowning and nonfatal submersion
C0013143|ICD9CM|AB|994.1|Drowning/nonfatal submer
C0013221|ICD9CM|PT|977.9|Poisoning by unspecified drug or medicinal substance
C0013221|ICD9CM|AB|977.9|Poison-medicinal agt NOS
C0013240|ICD9CM|AB|526.5|Alveolitis of jaw
C0013240|ICD9CM|PT|526.5|Alveolitis of jaw
C0013261|ICD9CM|AB|378.71|Duane's syndrome
C0013261|ICD9CM|PT|378.71|Duane's syndrome
C0013274|ICD9CM|AB|747.0|Patent ductus arteriosus
C0013274|ICD9CM|PT|747.0|Patent ductus arteriosus
C0013295|ICD9CM|HT|532|Duodenal ulcer
C0013298|ICD9CM|HT|535.6|Duodenitis
C0013312|ICD9CM|PT|728.6|Contracture of palmar fascia
C0013312|ICD9CM|AB|728.6|Contracted palmar fascia
C0013338|ICD9CM|AB|253.3|Pituitary dwarfism
C0013338|ICD9CM|PT|253.3|Pituitary dwarfism
C0013362|ICD9CM|PT|784.51|Dysarthria
C0013362|ICD9CM|AB|784.51|Dysarthria
C0013362|ICD9CM|AB|438.13|Late eff CV-dysarthria
C0013362|ICD9CM|PT|438.13|Late effects of cerebrovascular disease, dysarthria
C0013369|ICD9CM|PT|009.2|Infectious diarrhea
C0013369|ICD9CM|AB|009.2|Infectious diarrhea NOS
C0013371|ICD9CM|HT|004|Shigellosis
C0013371|ICD9CM|AB|004.9|Shigellosis NOS
C0013371|ICD9CM|PT|004.9|Shigellosis, unspecified
C0013373|ICD9CM|PT|780.56|Dysfunctions associated with sleep stages or arousal from sleep
C0013373|ICD9CM|AB|780.56|Sleep stage dysfunctions
C0013390|ICD9CM|AB|625.3|Dysmenorrhea
C0013390|ICD9CM|PT|625.3|Dysmenorrhea
C0013394|ICD9CM|AB|625.0|Dyspareunia
C0013394|ICD9CM|PT|625.0|Dyspareunia
C0013396|ICD9CM|PT|536.8|Dyspepsia and other specified disorders of function of stomach
C0013396|ICD9CM|AB|536.8|Stomach function dis NEC
C0013404|ICD9CM|AB|786.05|Shortness of breath
C0013404|ICD9CM|PT|786.05|Shortness of breath
C0013415|ICD9CM|AB|300.4|Dysthymic disorder
C0013415|ICD9CM|PT|300.4|Dysthymic disorder
C0013418|ICD9CM|HT|661.9|Unspecified abnormality of labor
C0013423|ICD9CM|PT|333.6|Genetic torsion dystonia
C0013423|ICD9CM|AB|333.6|Genetic torsion dystonia
C0013426|ICD9CM|HT|624.0|Dystrophy of vulva
C0013428|ICD9CM|AB|788.1|Dysuria
C0013428|ICD9CM|PT|788.1|Dysuria
C0013447|ICD9CM|PT|388.9|Unspecified disorder of ear
C0013447|ICD9CM|AB|388.9|Disorder of ear NOS
C0013456|ICD9CM|HT|388.7|Otalgia
C0013456|ICD9CM|AB|388.70|Otalgia NOS
C0013456|ICD9CM|PT|388.70|Otalgia, unspecified
C0013473|ICD9CM|AB|307.50|Eating disorder NOS
C0013473|ICD9CM|PT|307.50|Eating disorder, unspecified
C0013481|ICD9CM|AB|746.2|Ebstein's anomaly
C0013481|ICD9CM|PT|746.2|Ebstein's anomaly
C0013502|ICD9CM|HT|122|Echinococcosis
C0013504|ICD9CM|PT|122.8|Echinococcosis, unspecified, of liver
C0013504|ICD9CM|AB|122.8|Echinococcosis NOS liver
C0013515|ICD9CM|PT|079.1|Echo virus infection in conditions classified elsewhere and of unspecified site
C0013515|ICD9CM|AB|079.1|Echo virus infect NOS
C0013516|ICD9CM|PT|88.72|Diagnostic ultrasound of heart
C0013516|ICD9CM|AB|88.72|Dx ultrasound-heart
C0013570|ICD9CM|AB|051.2|Contagious pustular derm
C0013570|ICD9CM|PT|051.2|Contagious pustular dermatitis
C0013575|ICD9CM|PT|757.31|Congenital ectodermal dysplasia
C0013575|ICD9CM|AB|757.31|Cong ectodermal dysplas
C0013581|ICD9CM|AB|743.37|Congenital ectopic lens
C0013581|ICD9CM|PT|743.37|Congenital ectopic lens
C0013592|ICD9CM|HT|374.1|Ectropion
C0013592|ICD9CM|AB|374.10|Ectropion NOS
C0013592|ICD9CM|PT|374.10|Ectropion, unspecified
C0013604|ICD9CM|AB|782.3|Edema
C0013604|ICD9CM|PT|782.3|Edema
C0013654|ICD9CM|PT|V62.3|Educational circumstances
C0013654|ICD9CM|AB|V62.3|Educational circumstance
C0013679|ICD9CM|HT|990-995.99|OTHER AND UNSPECIFIED EFFECTS OF EXTERNAL CAUSES
C0013679|ICD9CM|HT|994|Effects of other external causes
C0013680|ICD9CM|AB|994.3|Effects of thirst
C0013680|ICD9CM|PT|994.3|Effects of thirst
C0013720|ICD9CM|PT|756.83|Ehlers-Danlos syndrome
C0013720|ICD9CM|AB|756.83|Ehlers-danlos syndrome
C0013778|ICD9CM|HT|99.6|Conversion of cardiac rhythm
C0013798|ICD9CM|AB|89.52|Electrocardiogram
C0013798|ICD9CM|PT|89.52|Electrocardiogram
C0013805|ICD9CM|AB|20.31|Electrocochleography
C0013805|ICD9CM|PT|20.31|Electrocochleography
C0013819|ICD9CM|AB|89.14|Electroencephalogram
C0013819|ICD9CM|PT|89.14|Electroencephalogram
C0013839|ICD9CM|AB|93.08|Electromyography
C0013839|ICD9CM|PT|93.08|Electromyography
C0013853|ICD9CM|PT|95.24|Electronystagmogram [ENG]
C0013853|ICD9CM|AB|95.24|Electronystagmogram
C0013854|ICD9CM|PT|95.22|Electro-oculogram [EOG]
C0013854|ICD9CM|AB|95.22|Electro-oculogram
C0013867|ICD9CM|PT|95.21|Electroretinogram [ERG]
C0013867|ICD9CM|AB|95.21|Electroretinogram
C0013902|ICD9CM|PT|282.1|Hereditary elliptocytosis
C0013902|ICD9CM|AB|282.1|Heredit elliptocytosis
C0013903|ICD9CM|AB|756.55|Chondroectoderm dysplas
C0013903|ICD9CM|PT|756.55|Chondroectodermal dysplasia
C0013923|ICD9CM|HT|444.0|Embolism and thrombosis of abdominal aorta
C0013924|ICD9CM|PT|444.9|Embolism and thrombosis of unspecified artery
C0013924|ICD9CM|AB|444.9|Arterial embolism NOS
C0013927|ICD9CM|HT|673.1|Amniotic fluid embolism
C0013927|ICD9CM|PT|673.10|Amniotic fluid embolism, unspecified as to episode of care or not applicable
C0013927|ICD9CM|AB|673.10|Amniotic embolism-unspec
C0013946|ICD9CM|PT|752.11|Embryonic cyst of fallopian tubes and broad ligaments
C0013946|ICD9CM|AB|752.11|Embryonic cyst of adnexa
C0014009|ICD9CM|HT|510|Empyema
C0014053|ICD9CM|AB|062.5|California encephalitis
C0014053|ICD9CM|PT|062.5|California virus encephalitis
C0014054|ICD9CM|PT|063.2|Central european encephalitis
C0014054|ICD9CM|AB|063.2|Cent Europe encephalitis
C0014057|ICD9CM|AB|062.0|Japanese encephalitis
C0014057|ICD9CM|PT|062.0|Japanese encephalitis
C0014058|ICD9CM|HT|323|Encephalitis, myelitis, and encephalomyelitis
C0014060|ICD9CM|PT|062.3|St. Louis encephalitis
C0014060|ICD9CM|AB|062.3|St Louis encephalitis
C0014061|ICD9CM|HT|063|Tick-borne viral encephalitis
C0014061|ICD9CM|PT|063.9|Tick-borne viral encephalitis, unspecified
C0014061|ICD9CM|AB|063.9|Tick-borne enceph NOS
C0014078|ICD9CM|AB|066.2|Venezuelan equine fever
C0014078|ICD9CM|PT|066.2|Venezuelan equine fever
C0014089|ICD9CM|AB|307.7|Encopresis
C0014089|ICD9CM|PT|307.7|Encopresis
C0014098|ICD9CM|HT|38.1|Endarterectomy
C0014116|ICD9CM|HT|745.6|Endocardial cushion defects
C0014116|ICD9CM|PT|745.60|Endocardial cushion defect, unspecified type
C0014116|ICD9CM|AB|745.60|Endocard cushion def NOS
C0014117|ICD9CM|PT|425.3|Endocardial fibroelastosis
C0014117|ICD9CM|AB|425.3|Endocard fibroelastosis
C0014130|ICD9CM|AB|259.9|Endocrine disorder NOS
C0014130|ICD9CM|PT|259.9|Unspecified endocrine disorder
C0014169|ICD9CM|AB|20.71|Endolymphatic shunt
C0014169|ICD9CM|PT|20.71|Endolymphatic shunt
C0014173|ICD9CM|HT|621.3|Endometrial hyperplasia
C0014173|ICD9CM|PT|621.30|Endometrial hyperplasia, unspecified
C0014173|ICD9CM|AB|621.30|Endometrial hyperpla NOS
C0014175|ICD9CM|HT|617|Endometriosis
C0014175|ICD9CM|AB|617.9|Endometriosis NOS
C0014175|ICD9CM|PT|617.9|Endometriosis, site unspecified
C0014177|ICD9CM|PT|617.2|Endometriosis of fallopian tube
C0014177|ICD9CM|AB|617.2|Tubal endometriosis
C0014178|ICD9CM|PT|617.8|Endometriosis of other specified sites
C0014178|ICD9CM|AB|617.8|Endometriosis NEC
C0014238|ICD9CM|PT|360.13|Parasitic endophthalmitis NOS
C0014238|ICD9CM|AB|360.13|Parasitic endophthal NOS
C0014306|ICD9CM|HT|376.5|Enophthalmos
C0014306|ICD9CM|AB|376.50|Enophthalmos NOS
C0014306|ICD9CM|PT|376.50|Enophthalmos, unspecified as to cause
C0014329|ICD9CM|PT|96.6|Enteral infusion of concentrated nutritional substances
C0014329|ICD9CM|AB|96.6|Entral infus nutrit sub
C0014370|ICD9CM|PT|46.01|Exteriorization of small intestine
C0014370|ICD9CM|AB|46.01|Sm bowel exteriorization
C0014390|ICD9CM|AB|374.00|Entropion NOS
C0014390|ICD9CM|PT|374.00|Entropion, unspecified
C0014394|ICD9CM|AB|307.6|Enuresis
C0014394|ICD9CM|PT|307.6|Enuresis
C0014457|ICD9CM|AB|288.3|Eosinophilia
C0014457|ICD9CM|PT|288.3|Eosinophilia
C0014493|ICD9CM|PT|077.1|Epidemic keratoconjunctivitis
C0014493|ICD9CM|AB|077.1|Epidem keratoconjunctiv
C0014498|ICD9CM|PT|078.82|Epidemic vomiting syndrome
C0014498|ICD9CM|AB|078.82|Epidemic vomiting synd
C0014511|ICD9CM|AB|706.2|Sebaceous cyst
C0014511|ICD9CM|PT|706.2|Sebaceous cyst
C0014518|ICD9CM|PT|695.15|Toxic epidermal necrolysis
C0014518|ICD9CM|AB|695.15|Toxic epidrml necrolysis
C0014544|ICD9CM|HT|345.9|Epilepsy, unspecified
C0014586|ICD9CM|AB|73.6|Episiotomy
C0014586|ICD9CM|PT|73.6|Episiotomy
C0014591|ICD9CM|AB|784.7|Epistaxis
C0014591|ICD9CM|PT|784.7|Epistaxis
C0014719|ICD9CM|PT|622.0|Erosion and ectropion of cervix
C0014719|ICD9CM|AB|622.0|Erosion/ectropion cervix
C0014733|ICD9CM|AB|035|Erysipelas
C0014733|ICD9CM|PT|035|Erysipelas
C0014736|ICD9CM|AB|027.1|Erysipelothrix infection
C0014736|ICD9CM|PT|027.1|Erysipelothrix infection
C0014742|ICD9CM|HT|695.1|Erythema multiforme
C0014742|ICD9CM|AB|695.10|Erythema multiforme NOS
C0014742|ICD9CM|PT|695.10|Erythema multiforme, unspecified
C0014743|ICD9CM|AB|695.2|Erythema nodosum
C0014743|ICD9CM|PT|695.2|Erythema nodosum
C0014744|ICD9CM|HT|017.1|Erythema nodosum with hypersensitivity reaction in tuberculosis
C0014744|ICD9CM|AB|017.10|Erythema nodos tb-unspec
C0014744|ICD9CM|PT|017.10|Erythema nodosum with hypersensitivity reaction in tuberculosis, unspecified
C0014747|ICD9CM|HT|690|Erythematosquamous dermatosis
C0014761|ICD9CM|HT|773|Hemolytic disease of fetus or newborn, due to isoimmunization
C0014761|ICD9CM|PT|773.2|Hemolytic disease of fetus or newborn due to other and unspecified isoimmunization
C0014761|ICD9CM|AB|773.2|NB hemolyt dis-isoim NEC
C0014804|ICD9CM|AB|443.82|Erythromelalgia
C0014804|ICD9CM|PT|443.82|Erythromelalgia
C0014835|ICD9CM|HT|041.4|Escherichia coli [E. coli] infection in conditions classified elsewhere and of unspecified site
C0014836|ICD9CM|PT|041.49|Other and unspecified Escherichia coli [E. coli]
C0014836|ICD9CM|AB|041.49|E.coli infection NEC/NOS
C0014848|ICD9CM|PT|530.0|Achalasia and cardiospasm
C0014848|ICD9CM|AB|530.0|Achalasia & cardiospasm
C0014852|ICD9CM|AB|530.9|Esophageal disorder NOS
C0014852|ICD9CM|HT|530|Diseases of esophagus
C0014852|ICD9CM|PT|530.9|Unspecified disorder of esophagus
C0014858|ICD9CM|AB|530.5|Dyskinesia of esophagus
C0014858|ICD9CM|PT|530.5|Dyskinesia of esophagus
C0014860|ICD9CM|AB|530.4|Perforation of esophagus
C0014860|ICD9CM|PT|530.4|Perforation of esophagus
C0014864|ICD9CM|PT|93.73|Esophageal speech training
C0014864|ICD9CM|AB|93.73|Esophag speech training
C0014868|ICD9CM|HT|530.1|Esophagitis
C0014868|ICD9CM|AB|530.10|Esophagitis, unspecified
C0014868|ICD9CM|PT|530.10|Esophagitis, unspecified
C0014869|ICD9CM|AB|530.11|Reflux esophagitis
C0014869|ICD9CM|PT|530.11|Reflux esophagitis
C0014875|ICD9CM|HT|42.1|Esophagostomy
C0014875|ICD9CM|AB|42.10|Esophagostomy NOS
C0014875|ICD9CM|PT|42.10|Esophagostomy, not otherwise specified
C0014877|ICD9CM|HT|378.0|Esotropia
C0014877|ICD9CM|AB|378.00|Esotropia NOS
C0014877|ICD9CM|PT|378.00|Esotropia, unspecified
C0015190|ICD9CM|AB|790.94|Euthyroid sick syndrome
C0015190|ICD9CM|PT|790.94|Euthyroid sick syndrome
C0015222|ICD9CM|HT|V72.1|Examination of ears and hearing
C0015230|ICD9CM|PT|782.1|Rash and other nonspecific skin eruption
C0015230|ICD9CM|AB|782.1|Nonspecif skin erupt NEC
C0015231|ICD9CM|HT|058.1|Roseola infantum
C0015231|ICD9CM|AB|058.10|Roseola infantum NOS
C0015231|ICD9CM|PT|058.10|Roseola infantum, unspecified
C0015233|ICD9CM|PT|E901.0|Accident due to excessive cold due to weather conditions
C0015233|ICD9CM|AB|E901.0|Excessive cold: weather
C0015236|ICD9CM|AB|99.01|Exchange transfusion
C0015236|ICD9CM|PT|99.01|Exchange transfusion
C0015263|ICD9CM|PT|493.81|Exercise induced bronchospasm
C0015263|ICD9CM|AB|493.81|Exercse ind bronchospasm
C0015269|ICD9CM|AB|302.4|Exhibitionism
C0015269|ICD9CM|PT|302.4|Exhibitionism
C0015300|ICD9CM|AB|376.30|Exophthalmos NOS
C0015300|ICD9CM|PT|376.30|Exophthalmos, unspecified
C0015310|ICD9CM|HT|378.1|Exotropia
C0015310|ICD9CM|AB|378.10|Exotropia NOS
C0015310|ICD9CM|PT|378.10|Exotropia, unspecified
C0015332|ICD9CM|PT|E926.8|Exposure to other specified radiation
C0015332|ICD9CM|AB|E926.8|Radiation exposure NEC
C0015333|ICD9CM|HT|E926|Exposure to radiation
C0015333|ICD9CM|AB|E926.9|Radiation exposure NOS
C0015333|ICD9CM|PT|E926.9|Exposure to unspecified radiation
C0015335|ICD9CM|PT|E926.2|Exposure to visible and ultraviolet light sources
C0015335|ICD9CM|AB|E926.2|Vis/ultraviol lght expos
C0015355|ICD9CM|PT|39.61|Extracorporeal circulation auxiliary to open heart surgery
C0015355|ICD9CM|AB|39.61|Extracorporeal circulat
C0015357|ICD9CM|PT|39.65|Extracorporeal membrane oxygenation [ECMO]
C0015357|ICD9CM|AB|39.65|Extracorporeal memb oxy
C0015359|ICD9CM|HT|98.5|Extracorporeal shockwave lithotripsy [ESWL]
C0015359|ICD9CM|PT|59.95|Ultrasonic fragmentation of urinary stones
C0015359|ICD9CM|AB|59.95|Ultrason fragment-stone
C0015393|ICD9CM|HT|743|Congenital anomalies of eye
C0015393|ICD9CM|PT|743.9|Unspecified anomaly of eye
C0015393|ICD9CM|AB|743.9|Eye anomaly NOS
C0015397|ICD9CM|AB|379.90|Eye disorder NOS
C0015397|ICD9CM|HT|360|Disorders of the globe
C0015397|ICD9CM|AB|360.9|Disorder of globe NOS
C0015397|ICD9CM|PT|360.9|Unspecified disorder of globe
C0015397|ICD9CM|PT|379.90|Disorder of eye, unspecified
C0015400|ICD9CM|HT|16.4|Enucleation of eyeball
C0015401|ICD9CM|PT|360.60|Foreign body, intraocular, unspecified
C0015401|ICD9CM|AB|360.60|Intraocular FB NOS
C0015409|ICD9CM|PT|871.7|Unspecified ocular penetration
C0015409|ICD9CM|AB|871.7|Ocular penetration NOS
C0015423|ICD9CM|PT|374.9|Unspecified disorder of eyelid
C0015423|ICD9CM|AB|374.9|Disorder of eyelid NOS
C0015464|ICD9CM|HT|351|Facial nerve disorders
C0015464|ICD9CM|PT|351.9|Facial nerve disorder, unspecified
C0015464|ICD9CM|AB|351.9|Facial nerve dis NOS
C0015481|ICD9CM|PT|300.16|Factitious disorder with predominantly psychological signs and symptoms
C0015481|ICD9CM|AB|300.16|Factitious dis w symptom
C0015523|ICD9CM|PT|286.2|Congenital factor XI deficiency
C0015523|ICD9CM|AB|286.2|Cong factor xi disorder
C0015544|ICD9CM|PT|783.41|Failure to thrive
C0015544|ICD9CM|AB|783.41|Failure to thrive-child
C0015584|ICD9CM|AB|V19.7|Consanguinity
C0015584|ICD9CM|PT|V19.7|Family history of consanguinity
C0015618|ICD9CM|AB|94.42|Family therapy
C0015618|ICD9CM|PT|94.42|Family therapy
C0015632|ICD9CM|PT|063.0|Russian spring-summer [taiga] encephalitis
C0015632|ICD9CM|AB|063.0|Russia spr-summer enceph
C0015634|ICD9CM|AB|495.0|Farmers' lung
C0015634|ICD9CM|PT|495.0|Farmers' lung
C0015645|ICD9CM|AB|729.4|Fasciitis NOS
C0015645|ICD9CM|PT|729.4|Fasciitis, unspecified
C0015652|ICD9CM|AB|121.3|Fascioliasis
C0015652|ICD9CM|PT|121.3|Fascioliasis
C0015656|ICD9CM|AB|121.4|Fasciolopsiasis
C0015656|ICD9CM|PT|121.4|Fasciolopsiasis
C0015674|ICD9CM|AB|780.71|Chronic fatigue syndrome
C0015674|ICD9CM|PT|780.71|Chronic fatigue syndrome
C0015696|ICD9CM|AB|571.0|Alcoholic fatty liver
C0015696|ICD9CM|PT|571.0|Alcoholic fatty liver
C0015732|ICD9CM|HT|787.6|Incontinence of feces
C0015734|ICD9CM|PT|560.32|Fecal impaction
C0015734|ICD9CM|AB|560.32|Fecal impaction
C0015773|ICD9CM|AB|714.1|Felty's syndrome
C0015773|ICD9CM|PT|714.1|Felty's syndrome
C0015806|ICD9CM|HT|820|Fracture of neck of femur
C0015825|ICD9CM|HT|20.6|Fenestration of inner ear
C0015931|ICD9CM|HT|656.3|Fetal distress affecting management of mother
C0015934|ICD9CM|HT|764.9|Fetal growth retardation, unspecified
C0015934|ICD9CM|PT|764.90|Fetal growth retardation, unspecified, unspecified [weight]
C0015934|ICD9CM|AB|764.90|Fet growth retard wtNOS
C0015944|ICD9CM|HT|658.1|Premature rupture of membranes
C0015957|ICD9CM|AB|302.81|Fetishism
C0015957|ICD9CM|PT|302.81|Fetishism
C0015959|ICD9CM|PT|656.00|Fetal-maternal hemorrhage, unspecified as to episode of care or not applicable
C0015959|ICD9CM|AB|656.00|Fetal-maternal hem-unsp
C0015967|ICD9CM|AB|780.60|Fever NOS
C0015967|ICD9CM|PT|780.60|Fever, unspecified
C0016034|ICD9CM|PT|610.1|Diffuse cystic mastopathy
C0016034|ICD9CM|AB|610.1|Diffus cystic mastopathy
C0016037|ICD9CM|PT|728.11|Progressive myositis ossificans
C0016037|ICD9CM|AB|728.11|Prog myositis ossificans
C0016065|ICD9CM|PT|756.54|Polyostotic fibrous dysplasia of bone
C0016065|ICD9CM|AB|756.54|Polyostotic fibros dyspl
C0016085|ICD9CM|AB|125.9|Filariasis NOS
C0016085|ICD9CM|PT|125.9|Unspecified filariasis
C0016089|ICD9CM|PT|125.5|Mansonella ozzardi infection
C0016089|ICD9CM|AB|125.5|Mansonella ozzardi infec
C0016124|ICD9CM|PT|959.5|Finger injury
C0016124|ICD9CM|AB|959.5|Finger injury NOS
C0016142|ICD9CM|AB|312.33|Pyromania
C0016142|ICD9CM|PT|312.33|Pyromania
C0016167|ICD9CM|AB|565.0|Anal fissure
C0016167|ICD9CM|PT|565.0|Anal fissure
C0016171|ICD9CM|PT|569.81|Fistula of intestine, excluding rectum and anus
C0016171|ICD9CM|AB|569.81|Intestinal fistula
C0016196|ICD9CM|AB|807.4|Flail chest
C0016196|ICD9CM|PT|807.4|Flail chest
C0016205|ICD9CM|PT|787.3|Flatulence, eructation, and gas pain
C0016205|ICD9CM|AB|787.3|Flatul/eructat/gas pain
C0016234|ICD9CM|AB|45.24|Flexible sigmoidoscopy
C0016234|ICD9CM|PT|45.24|Flexible sigmoidoscopy
C0016382|ICD9CM|AB|782.62|Flushing
C0016382|ICD9CM|PT|782.62|Flushing
C0016429|ICD9CM|AB|620.0|Follicular cyst of ovary
C0016429|ICD9CM|PT|620.0|Follicular cyst of ovary
C0016479|ICD9CM|AB|005.9|Food poisoning NOS
C0016479|ICD9CM|PT|005.9|Food poisoning, unspecified
C0016514|ICD9CM|PT|078.4|Foot and mouth disease
C0016514|ICD9CM|AB|078.4|Foot & mouth disease
C0016545|ICD9CM|PT|728.82|Foreign body granuloma of muscle
C0016545|ICD9CM|AB|728.82|FB granuloma of muscle
C0016546|ICD9CM|PT|938|Foreign body in digestive system, unspecified
C0016546|ICD9CM|AB|938|Foreign body GI NOS
C0016574|ICD9CM|PT|56.61|Formation of other cutaneous ureterostomy
C0016574|ICD9CM|AB|56.61|Form cutan ureterostomy
C0016632|ICD9CM|AB|705.82|Fox-fordyce disease
C0016632|ICD9CM|PT|705.82|Fox-Fordyce disease
C0016644|ICD9CM|HT|814|Fracture of carpal bone(s)
C0016652|ICD9CM|PT|813.81|Closed fracture of unspecified part of radius (alone)
C0016652|ICD9CM|AB|813.81|Fx radius NOS-closed
C0016653|ICD9CM|PT|813.82|Closed fracture of unspecified part of ulna (alone)
C0016653|ICD9CM|AB|813.82|Fracture ulna NOS-closed
C0016658|ICD9CM|HT|800-829.99|FRACTURES
C0016658|ICD9CM|HT|829|Fracture of unspecified bones
C0016658|ICD9CM|AB|E887|Fracture, cause NOS
C0016658|ICD9CM|PT|E887|Fracture, cause unspecified
C0016659|ICD9CM|AB|829.0|Fracture NOS-closed
C0016659|ICD9CM|PT|829.0|Fracture of unspecified bone, closed
C0016662|ICD9CM|AB|829.1|Fracture NOS-open
C0016662|ICD9CM|PT|829.1|Fracture of unspecified bone, open
C0016663|ICD9CM|HT|733.1|Pathologic fracture
C0016663|ICD9CM|PT|733.10|Pathologic fracture, unspecified site
C0016663|ICD9CM|AB|733.10|Path fx unspecified site
C0016663|ICD9CM|AB|V13.51|Hx pathological fracture
C0016663|ICD9CM|PT|V13.51|Personal history of pathologic fracture
C0016665|ICD9CM|AB|733.82|Nonunion of fracture
C0016665|ICD9CM|PT|733.82|Nonunion of fracture
C0016667|ICD9CM|PT|759.83|Fragile X syndrome
C0016667|ICD9CM|AB|759.83|Fragile x syndrome
C0016708|ICD9CM|HT|788.4|Frequency of urination and polyuria
C0016719|ICD9CM|AB|334.0|Friedreich's ataxia
C0016719|ICD9CM|PT|334.0|Friedreich's ataxia
C0016737|ICD9CM|PT|991.3|Frostbite of other and unspecified sites
C0016737|ICD9CM|AB|991.3|Frostbite NEC/NOS
C0016751|ICD9CM|PT|271.2|Hereditary fructose intolerance
C0016751|ICD9CM|AB|271.2|Hered fructose intoleran
C0016782|ICD9CM|PT|364.21|Fuchs' heterochromic cyclitis
C0016782|ICD9CM|AB|364.21|Fuch hetrochrom cyclitis
C0016807|ICD9CM|PT|564.9|Unspecified functional disorder of intestine
C0016807|ICD9CM|AB|564.9|Funct dis intestine NOS
C0016808|ICD9CM|PT|288.1|Functional disorders of polymorphonuclear neutrophils
C0016808|ICD9CM|AB|288.1|Function dis neutrophils
C0016809|ICD9CM|PT|429.4|Functional disturbances following cardiac surgery
C0016809|ICD9CM|AB|429.4|Hrt dis postcardiac surg
C0016842|ICD9CM|AB|754.81|Pectus excavatum
C0016842|ICD9CM|PT|754.81|Pectus excavatum
C0016952|ICD9CM|AB|271.1|Galactosemia
C0016952|ICD9CM|PT|271.1|Galactosemia
C0016977|ICD9CM|PT|575.9|Unspecified disorder of gallbladder
C0016977|ICD9CM|AB|575.9|Dis of gallbladder NOS
C0017086|ICD9CM|AB|785.4|Gangrene
C0017086|ICD9CM|PT|785.4|Gangrene
C0017105|ICD9CM|AB|040.0|Gas gangrene
C0017105|ICD9CM|PT|040.0|Gas gangrene
C0017131|ICD9CM|AB|96.32|Gastric freezing
C0017131|ICD9CM|PT|96.32|Gastric freezing
C0017131|ICD9CM|AB|96.31|Gastric cooling
C0017131|ICD9CM|PT|96.31|Gastric cooling
C0017134|ICD9CM|AB|96.33|Gastric lavage
C0017134|ICD9CM|PT|96.33|Gastric lavage
C0017154|ICD9CM|HT|535.1|Atrophic gastritis
C0017155|ICD9CM|HT|535.2|Gastric mucosal hypertrophy
C0017166|ICD9CM|HT|44.3|Gastroenterostomy without gastrectomy
C0017168|ICD9CM|AB|530.81|Esophageal reflux
C0017168|ICD9CM|PT|530.81|Esophageal reflux
C0017181|ICD9CM|HT|578|Gastrointestinal hemorrhage
C0017181|ICD9CM|AB|578.9|Gastrointest hemorr NOS
C0017181|ICD9CM|PT|578.9|Hemorrhage of gastrointestinal tract, unspecified
C0017183|ICD9CM|PT|306.4|Gastrointestinal malfunction arising from mental factors
C0017183|ICD9CM|AB|306.4|Psychogenic GI disease
C0017196|ICD9CM|HT|43.1|Gastrostomy
C0017327|ICD9CM|AB|440.9|Atherosclerosis NOS
C0017327|ICD9CM|PT|440.9|Generalized and unspecified atherosclerosis
C0017332|ICD9CM|HT|345.0|Generalized nonconvulsive epilepsy
C0017377|ICD9CM|PT|288.2|Genetic anomalies of leukocytes
C0017377|ICD9CM|AB|288.2|Genetic anomaly leukocyt
C0017394|MTH|PN|NOCODE|Encounter for Genetic screening NEC in ICD9CM
C0017394|ICD9CM|HT|V82.7|Genetic screening
C0017394|ICD9CM|PT|V82.79|Other genetic screening
C0017394|ICD9CM|AB|V82.79|Genetic screening NEC
C0017407|ICD9CM|AB|351.1|Geniculate ganglionitis
C0017407|ICD9CM|PT|351.1|Geniculate ganglionitis
C0017409|ICD9CM|AB|053.11|Geniculate herpes zoster
C0017409|ICD9CM|PT|053.11|Geniculate herpes zoster
C0017411|ICD9CM|PT|629.9|Unspecified disorder of female genital organs
C0017411|ICD9CM|AB|629.9|Female genital dis NOS
C0017412|ICD9CM|PT|608.9|Unspecified disorder of male genital organs
C0017412|ICD9CM|HT|600-608.99|DISEASES OF MALE GENITAL ORGANS
C0017412|ICD9CM|AB|608.9|Male genital dis NOS
C0017418|ICD9CM|AB|091.0|Primary genital syphilis
C0017418|ICD9CM|PT|091.0|Genital syphilis (primary)
C0017495|ICD9CM|PT|046.71|Gerstmann-Sträussler-Scheinker syndrome
C0017495|ICD9CM|AB|046.71|Gerstmn-Straus-Schnk syn
C0017536|ICD9CM|AB|007.1|Giardiasis
C0017536|ICD9CM|PT|007.1|Giardiasis
C0017572|ICD9CM|HT|523.2|Gingival recession
C0017572|ICD9CM|AB|523.20|Gingival recession NOS
C0017572|ICD9CM|PT|523.20|Gingival recession, unspecified
C0017576|ICD9CM|AB|24.2|Gingivoplasty
C0017576|ICD9CM|PT|24.2|Gingivoplasty
C0017589|ICD9CM|AB|024|Glanders
C0017589|ICD9CM|PT|024|Glanders
C0017601|ICD9CM|HT|365|Glaucoma
C0017601|ICD9CM|AB|365.9|Glaucoma NOS
C0017601|ICD9CM|PT|365.9|Unspecified glaucoma
C0017606|ICD9CM|HT|365.2|Primary angle-closure glaucoma
C0017606|ICD9CM|PT|365.20|Primary angle-closure glaucoma, unspecified
C0017606|ICD9CM|AB|365.20|Prim angl-clos glauc NOS
C0017612|ICD9CM|HT|365.1|Open-angle glaucoma
C0017612|ICD9CM|AB|365.10|Open-angle glaucoma NOS
C0017612|ICD9CM|PT|365.13|Pigmentary open-angle glaucoma
C0017612|ICD9CM|AB|365.13|Pigmentary glaucoma
C0017612|ICD9CM|PT|365.10|Open-angle glaucoma, unspecified
C0017672|ICD9CM|AB|529.6|Glossodynia
C0017672|ICD9CM|PT|529.6|Glossodynia
C0017675|ICD9CM|AB|529.0|Glossitis
C0017675|ICD9CM|PT|529.0|Glossitis
C0017677|ICD9CM|AB|529.1|Geographic tongue
C0017677|ICD9CM|PT|529.1|Geographic tongue
C0017919|ICD9CM|AB|271.0|Glycogenosis
C0017919|ICD9CM|PT|271.0|Glycogenosis
C0017979|ICD9CM|AB|791.5|Glycosuria
C0017979|ICD9CM|PT|791.5|Glycosuria
C0017980|ICD9CM|AB|271.4|Renal glycosuria
C0017980|ICD9CM|PT|271.4|Renal glycosuria
C0018013|ICD9CM|AB|128.1|Gnathostomiasis
C0018013|ICD9CM|PT|128.1|Gnathostomiasis
C0018021|ICD9CM|AB|240.9|Goiter NOS
C0018021|ICD9CM|PT|240.9|Goiter, unspecified
C0018022|ICD9CM|AB|240.0|Simple goiter
C0018022|ICD9CM|PT|240.0|Goiter, specified as simple
C0018041|ICD9CM|AB|E006.2|Golf
C0018041|ICD9CM|PT|E006.2|Activities involving golf
C0018051|ICD9CM|AB|758.6|Gonadal dysgenesis
C0018051|ICD9CM|PT|758.6|Gonadal dysgenesis
C0018074|ICD9CM|PT|098.0|Gonococcal infection (acute) of lower genitourinary tract
C0018074|ICD9CM|AB|098.0|Acute gc infect lower gu
C0018075|ICD9CM|AB|098.81|Gonococcal keratosis
C0018075|ICD9CM|PT|098.81|Gonococcal keratosis (blennorrhagica)
C0018077|ICD9CM|AB|098.86|Gonococcal peritonitis
C0018077|ICD9CM|PT|098.86|Gonococcal peritonitis
C0018081|ICD9CM|HT|098|Gonococcal infections
C0018099|ICD9CM|HT|274|Gout
C0018099|ICD9CM|AB|274.9|Gout NOS
C0018099|ICD9CM|PT|274.9|Gout, unspecified
C0018133|ICD9CM|HT|279.5|Graft-versus-host disease
C0018133|ICD9CM|AB|279.50|Graft-versus-host NOS
C0018133|ICD9CM|PT|279.50|Graft-versus-host disease, unspecified
C0018179|ICD9CM|PT|371.53|Granular corneal dystrophy
C0018179|ICD9CM|AB|371.53|Granular cornea dystrphy
C0018190|ICD9CM|AB|099.2|Granuloma inguinale
C0018190|ICD9CM|PT|099.2|Granuloma inguinale
C0018197|ICD9CM|AB|446.3|Lethal midline granuloma
C0018197|ICD9CM|PT|446.3|Lethal midline granuloma
C0018409|ICD9CM|AB|E005.2|Gymnastics
C0018409|ICD9CM|PT|E005.2|Activities involving gymnastics
C0018524|ICD9CM|AB|780.1|Hallucinations
C0018524|ICD9CM|PT|780.1|Hallucinations
C0018526|ICD9CM|HT|305.3|Hallucinogen abuse
C0018528|ICD9CM|HT|304.5|Hallucinogen dependence
C0018528|ICD9CM|PT|304.50|Hallucinogen dependence, unspecified
C0018528|ICD9CM|AB|304.50|Hallucinogen dep-unspec
C0018572|ICD9CM|PT|074.3|Hand, foot, and mouth disease
C0018572|ICD9CM|AB|074.3|Hand, foot & mouth dis
C0018621|ICD9CM|PT|477.0|Allergic rhinitis due to pollen
C0018621|ICD9CM|AB|477.0|Rhinitis due to pollen
C0018674|ICD9CM|AB|959.01|Head injury NOS
C0018674|ICD9CM|PT|959.01|Head injury, unspecified
C0018681|ICD9CM|AB|784.0|Headache
C0018681|ICD9CM|PT|784.0|Headache
C0018776|ICD9CM|AB|389.14|Central hearing loss
C0018776|ICD9CM|PT|389.14|Central hearing loss
C0018777|ICD9CM|HT|389.0|Conductive hearing loss
C0018777|ICD9CM|PT|389.00|Conductive hearing loss, unspecified
C0018777|ICD9CM|AB|389.00|Conduct hearing loss NOS
C0018781|ICD9CM|PT|388.12|Noise-induced hearing loss
C0018781|ICD9CM|AB|388.12|Hearing loss d/t noise
C0018784|ICD9CM|HT|389.1|Sensorineural hearing loss
C0018784|ICD9CM|PT|389.10|Sensorineural hearing loss, unspecified
C0018784|ICD9CM|AB|389.10|Sensorneur hear loss NOS
C0018786|ICD9CM|AB|95.47|Hearing examination NOS
C0018786|ICD9CM|PT|95.42|Clinical test of hearing
C0018786|ICD9CM|AB|95.42|Clinical hearing test
C0018786|ICD9CM|PT|95.47|Hearing examination, not otherwise specified
C0018790|ICD9CM|AB|427.5|Cardiac arrest
C0018790|ICD9CM|PT|427.5|Cardiac arrest
C0018791|ICD9CM|AB|39.63|Cardioplegia
C0018791|ICD9CM|PT|39.63|Cardioplegia
C0018798|ICD9CM|PT|746.9|Unspecified congenital anomaly of heart
C0018798|ICD9CM|AB|746.9|Cong heart anomaly NOS
C0018799|ICD9CM|AB|429.9|Heart disease NOS
C0018799|ICD9CM|PT|429.9|Heart disease, unspecified
C0018800|ICD9CM|AB|429.3|Cardiomegaly
C0018800|ICD9CM|PT|429.3|Cardiomegaly
C0018801|ICD9CM|HT|428|Heart failure
C0018801|ICD9CM|AB|428.9|Heart failure NOS
C0018801|ICD9CM|PT|428.9|Heart failure, unspecified
C0018802|ICD9CM|AB|428.0|CHF NOS
C0018802|ICD9CM|PT|428.0|Congestive heart failure, unspecified
C0018812|ICD9CM|PT|V42.1|Heart replaced by transplant
C0018812|ICD9CM|AB|V42.1|Heart transplant status
C0018818|ICD9CM|PT|745.4|Ventricular septal defect
C0018818|ICD9CM|AB|745.4|Ventricular sept defect
C0018823|ICD9CM|AB|37.51|Heart transplantation
C0018823|ICD9CM|PT|37.51|Heart transplantation
C0018833|ICD9CM|PT|33.6|Combined heart-lung transplantation
C0018833|ICD9CM|AB|33.6|Comb heart/lung transpla
C0018834|ICD9CM|AB|787.1|Heartburn
C0018834|ICD9CM|PT|787.1|Heartburn
C0018839|ICD9CM|AB|992.5|Heat exhaustion NOS
C0018839|ICD9CM|PT|992.5|Heat exhaustion, unspecified
C0018844|ICD9CM|PT|992.0|Heat stroke and sunstroke
C0018844|ICD9CM|AB|992.0|Heat stroke & sunstroke
C0018889|ICD9CM|HT|120-129.99|HELMINTHIASES
C0018889|ICD9CM|AB|128.9|Helminthiasis NOS
C0018889|ICD9CM|PT|128.9|Helminth infection, unspecified
C0018916|ICD9CM|AB|228.00|Hemangioma NOS
C0018916|ICD9CM|PT|228.00|Hemangioma of unspecified site
C0018916|ICD9CM|HT|228.0|Hemangioma, any site
C0018918|ICD9CM|PT|228.09|Hemangioma of other sites
C0018918|ICD9CM|AB|228.09|Hemangioma NEC
C0018924|ICD9CM|HT|719.1|Hemarthrosis
C0018924|ICD9CM|AB|719.10|Hemarthrosis-unspec
C0018924|ICD9CM|PT|719.10|Hemarthrosis, site unspecified
C0018926|ICD9CM|AB|578.0|Hematemesis
C0018926|ICD9CM|PT|578.0|Hematemesis
C0018939|ICD9CM|AB|289.9|Blood disease NOS
C0018939|ICD9CM|PT|289.9|Unspecified diseases of blood and blood-forming organs
C0018939|ICD9CM|HT|280-289.99|DISEASES OF THE BLOOD AND BLOOD-FORMING ORGANS
C0018946|ICD9CM|AB|432.1|Subdural hemorrhage
C0018946|ICD9CM|PT|432.1|Subdural hemorrhage
C0018948|ICD9CM|AB|621.4|Hematometra
C0018948|ICD9CM|PT|621.4|Hematometra
C0018965|ICD9CM|HT|599.7|Hematuria
C0018965|ICD9CM|AB|599.70|Hematuria NOS
C0018965|ICD9CM|PT|599.70|Hematuria, unspecified
C0018990|ICD9CM|PT|84.19|Abdominopelvic amputation
C0018990|ICD9CM|AB|84.19|Hindquarter amputation
C0018991|ICD9CM|HT|342.9|Hemiplegia, unspecified
C0019004|ICD9CM|AB|39.95|Hemodialysis
C0019004|ICD9CM|PT|39.95|Hemodialysis
C0019034|ICD9CM|PT|282.63|Sickle-cell/Hb-C disease without crisis
C0019034|ICD9CM|AB|282.63|Hb-SS/hb-C dis w/o crsis
C0019048|ICD9CM|AB|791.2|Hemoglobinuria
C0019048|ICD9CM|PT|791.2|Hemoglobinuria
C0019049|ICD9CM|PT|283.2|Hemoglobinuria due to hemolysis from external causes
C0019049|ICD9CM|AB|283.2|Hemolytic hemoglobinuria
C0019061|ICD9CM|PT|283.11|Hemolytic-uremic syndrome
C0019061|ICD9CM|AB|283.11|Hemolytic uremic synd
C0019064|ICD9CM|AB|423.0|Hemopericardium
C0019064|ICD9CM|PT|423.0|Hemopericardium
C0019066|ICD9CM|PT|568.81|Hemoperitoneum (nontraumatic)
C0019066|ICD9CM|AB|568.81|Hemoperitoneum
C0019069|ICD9CM|PT|286.0|Congenital factor VIII disorder
C0019069|ICD9CM|AB|286.0|Cong factor viii diord
C0019073|ICD9CM|PT|041.5|Hemophilus influenzae [H. influenzae] infection in conditions classified elsewhere and of unspecified site
C0019073|ICD9CM|AB|041.5|H. influenzae infect NOS
C0019079|ICD9CM|HT|786.3|Hemoptysis
C0019079|ICD9CM|AB|786.30|Hemoptysis NOS
C0019079|ICD9CM|PT|786.30|Hemoptysis, unspecified
C0019080|ICD9CM|AB|459.0|Hemorrhage NOS
C0019080|ICD9CM|PT|459.0|Hemorrhage, unspecified
C0019081|ICD9CM|PT|569.3|Hemorrhage of rectum and anus
C0019081|ICD9CM|AB|569.3|Rectal & anal hemorrhage
C0019087|ICD9CM|PT|287.9|Unspecified hemorrhagic conditions
C0019087|ICD9CM|AB|287.9|Hemorrhagic cond NOS
C0019088|ICD9CM|PT|776.0|Hemorrhagic disease of newborn
C0019088|ICD9CM|AB|776.0|NB hemorrhagic disease
C0019099|ICD9CM|PT|065.0|Crimean hemorrhagic fever [CHF Congo virus]
C0019099|ICD9CM|AB|065.0|Crimean hemorrhagic fev
C0019101|ICD9CM|PT|078.6|Hemorrhagic nephrosonephritis
C0019101|ICD9CM|AB|078.6|Hem nephrosonephritis
C0019103|ICD9CM|AB|065.1|Omsk hemorrhagic fever
C0019103|ICD9CM|PT|065.1|Omsk hemorrhagic fever
C0019108|ICD9CM|AB|49.46|Hemorrhoidectomy
C0019108|ICD9CM|PT|49.46|Excision of hemorrhoids
C0019112|ICD9CM|HT|455|Hemorrhoids
C0019151|ICD9CM|PT|572.2|Hepatic encephalopathy
C0019151|ICD9CM|AB|572.2|Hepatic encephalopathy
C0019158|ICD9CM|AB|573.3|Hepatitis NOS
C0019158|ICD9CM|PT|573.3|Hepatitis, unspecified
C0019189|ICD9CM|HT|571.4|Chronic hepatitis
C0019189|ICD9CM|AB|571.40|Chronic hepatitis NOS
C0019189|ICD9CM|PT|571.40|Chronic hepatitis, unspecified
C0019196|ICD9CM|HT|070.7|Unspecified viral hepatitis C
C0019209|ICD9CM|AB|789.1|Hepatomegaly
C0019209|ICD9CM|PT|789.1|Hepatomegaly
C0019212|ICD9CM|AB|572.4|Hepatorenal syndrome
C0019212|ICD9CM|PT|572.4|Hepatorenal syndrome
C0019275|ICD9CM|PT|553.9|Hernia of unspecified site without mention of obstruction or gangrene
C0019275|ICD9CM|AB|553.9|Hernia NOS
C0019275|ICD9CM|AB|553.8|Hernia NEC
C0019275|ICD9CM|PT|553.8|Hernia of other specified sites without mention of obstruction or gangrene
C0019294|ICD9CM|HT|550|Inguinal hernia
C0019328|ICD9CM|HT|53|Repair of hernia
C0019333|ICD9CM|HT|53.4|Repair of umbilical hernia
C0019338|ICD9CM|AB|074.0|Herpangina
C0019338|ICD9CM|PT|074.0|Herpangina
C0019342|ICD9CM|HT|054.1|Genital herpes
C0019342|ICD9CM|AB|054.10|Genital herpes NOS
C0019342|ICD9CM|PT|054.10|Genital herpes, unspecified
C0019348|ICD9CM|HT|054|Herpes simplex
C0019359|ICD9CM|AB|054.71|Visceral herpes simplex
C0019359|ICD9CM|PT|054.71|Visceral herpes simplex
C0019360|ICD9CM|HT|053|Herpes zoster
C0019362|ICD9CM|PT|053.20|Herpes zoster dermatitis of eyelid
C0019362|ICD9CM|AB|053.20|Herpes zoster of eyelid
C0019364|ICD9CM|HT|053.2|Herpes zoster with ophthalmic complications
C0019366|ICD9CM|PT|053.9|Herpes zoster without mention of complication
C0019366|ICD9CM|AB|053.9|Herpes zoster NOS
C0019385|ICD9CM|PT|054.3|Herpetic meningoencephalitis
C0019385|ICD9CM|AB|054.3|Herpetic encephalitis
C0019386|ICD9CM|AB|054.11|Herpetic vulvovaginitis
C0019386|ICD9CM|PT|054.11|Herpetic vulvovaginitis
C0019521|ICD9CM|AB|786.8|Hiccough
C0019521|ICD9CM|PT|786.8|Hiccough
C0019554|ICD9CM|HT|835|Dislocation of hip
C0019555|ICD9CM|HT|754.3|Congenital dislocation of hip
C0019570|ICD9CM|PT|751.3|Hirschsprung's disease and other congenital functional disorders of colon
C0019570|ICD9CM|AB|751.3|Hirschsprung's disease
C0019572|ICD9CM|AB|704.1|Hirsutism
C0019572|ICD9CM|PT|704.1|Hirsutism
C0019575|ICD9CM|AB|134.2|Hirudiniasis
C0019575|ICD9CM|PT|134.2|Hirudiniasis
C0019623|ICD9CM|HT|202.3|Malignant histiocytosis
C0019655|ICD9CM|HT|115|Histoplasmosis
C0019655|ICD9CM|HT|115.9|Histoplasmosis, unspecified
C0019657|ICD9CM|PT|115.99|Histoplasmosis, unspecified, other
C0019657|ICD9CM|AB|115.99|Histoplasmosis NEC
C0019681|ICD9CM|HT|301.5|Histrionic personality disorder
C0019681|ICD9CM|AB|301.50|Histrionic person NOS
C0019681|ICD9CM|PT|301.50|Histrionic personality disorder, unspecified
C0019693|ICD9CM|HT|042-042.99|HUMAN IMMUNODEFICIENCY VIRUS [HIV] INFECTION
C0019693|ICD9CM|PT|042|Human immunodeficiency virus [HIV] disease
C0019693|ICD9CM|AB|042|Human immuno virus dis
C0019829|ICD9CM|HT|201|Hodgkin's disease
C0019829|ICD9CM|HT|201.1|Hodgkin's granuloma
C0019829|ICD9CM|HT|201.0|Hodgkin's paragranuloma
C0019829|ICD9CM|HT|201.9|Hodgkin's disease, unspecified type
C0019918|ICD9CM|HT|373.1|Hordeolum and other deep inflammation of eyelid
C0019919|ICD9CM|AB|373.11|Hordeolum externum
C0019919|ICD9CM|PT|373.11|Hordeolum externum
C0020162|ICD9CM|HT|812|Fracture of humerus
C0020179|ICD9CM|AB|333.4|Huntington's chorea
C0020179|ICD9CM|PT|333.4|Huntington's chorea
C0020217|ICD9CM|AB|630|Hydatidiform mole
C0020217|ICD9CM|PT|630|Hydatidiform mole
C0020224|ICD9CM|HT|657.0|Polyhydramnios
C0020224|ICD9CM|HT|657|Polyhydramnios
C0020256|ICD9CM|AB|742.3|Congenital hydrocephalus
C0020256|ICD9CM|PT|742.3|Congenital hydrocephalus
C0020295|ICD9CM|AB|591|Hydronephrosis
C0020295|ICD9CM|PT|591|Hydronephrosis
C0020413|ICD9CM|AB|123.6|Hymenolepiasis
C0020413|ICD9CM|PT|123.6|Hymenolepiasis
C0020428|ICD9CM|HT|255.1|Hyperaldosteronism
C0020428|ICD9CM|AB|255.10|Hyperaldosteronism NOS
C0020428|ICD9CM|PT|255.10|Hyperaldosteronism, unspecified
C0020431|ICD9CM|AB|93.95|Hyperbaric oxygenation
C0020431|ICD9CM|PT|93.95|Hyperbaric oxygenation
C0020437|ICD9CM|AB|275.42|Hypercalcemia
C0020437|ICD9CM|PT|275.42|Hypercalcemia
C0020441|ICD9CM|AB|521.5|Hypercementosis
C0020441|ICD9CM|PT|521.5|Hypercementosis
C0020450|ICD9CM|HT|643|Excessive vomiting in pregnancy
C0020451|ICD9CM|HT|643.0|Mild hyperemesis gravidarum
C0020461|ICD9CM|AB|276.7|Hyperpotassemia
C0020461|ICD9CM|PT|276.7|Hyperpotassemia
C0020480|ICD9CM|AB|272.1|Pure hyperglyceridemia
C0020480|ICD9CM|PT|272.1|Pure hyperglyceridemia
C0020490|ICD9CM|AB|367.0|Hypermetropia
C0020490|ICD9CM|PT|367.0|Hypermetropia
C0020496|ICD9CM|AB|733.3|Hyperostosis of skull
C0020496|ICD9CM|PT|733.3|Hyperostosis of skull
C0020498|ICD9CM|PT|721.6|Ankylosing vertebral hyperostosis
C0020498|ICD9CM|AB|721.6|Ankyl vert hyperostosis
C0020502|ICD9CM|HT|252.0|Hyperparathyroidism
C0020502|ICD9CM|AB|252.00|Hyperparathyroidism NOS
C0020502|ICD9CM|PT|252.00|Hyperparathyroidism, unspecified
C0020505|ICD9CM|AB|783.6|Polyphagia
C0020505|ICD9CM|PT|783.6|Polyphagia
C0020532|ICD9CM|AB|289.4|Hypersplenism
C0020532|ICD9CM|PT|289.4|Hypersplenism
C0020534|ICD9CM|AB|376.41|Hypertelorism of orbit
C0020534|ICD9CM|PT|376.41|Hypertelorism of orbit
C0020538|ICD9CM|HT|401-405.99|HYPERTENSIVE DISEASE
C0020538|ICD9CM|PT|997.91|Complications affecting other specified body systems, not elsewhere classified, hypertension
C0020538|ICD9CM|AB|997.91|Surg comp - hypertension
C0020541|ICD9CM|AB|572.3|Portal hypertension
C0020541|ICD9CM|PT|572.3|Portal hypertension
C0020561|ICD9CM|PT|622.6|Hypertrophic elongation of cervix
C0020561|ICD9CM|AB|622.6|Hypertrophic elong cervx
C0020565|ICD9CM|AB|611.1|Hypertrophy of breast
C0020565|ICD9CM|PT|611.1|Hypertrophy of breast
C0020569|ICD9CM|PT|527.1|Hypertrophy of salivary gland
C0020569|ICD9CM|AB|527.1|Salivary glnd hyprtrophy
C0020575|ICD9CM|AB|378.31|Hypertropia
C0020575|ICD9CM|PT|378.31|Hypertropia
C0020578|ICD9CM|AB|786.01|Hyperventilation
C0020578|ICD9CM|PT|786.01|Hyperventilation
C0020579|ICD9CM|PT|278.2|Hypervitaminosis A
C0020579|ICD9CM|AB|278.2|Hypervitaminosis a
C0020582|ICD9CM|PT|364.41|Hyphema of iris and ciliary body
C0020582|ICD9CM|AB|364.41|Hyphema
C0020587|ICD9CM|AB|94.32|Hypnotherapy
C0020587|ICD9CM|PT|94.32|Hypnotherapy
C0020594|ICD9CM|PT|302.71|Hypoactive sexual desire disorder
C0020594|ICD9CM|AB|302.71|Hypoactive sex desire
C0020598|ICD9CM|AB|275.41|Hypocalcemia
C0020598|ICD9CM|PT|275.41|Hypocalcemia
C0020604|ICD9CM|AB|300.7|Hypochondriasis
C0020604|ICD9CM|PT|300.7|Hypochondriasis
C0020615|ICD9CM|AB|251.2|Hypoglycemia NOS
C0020615|ICD9CM|PT|251.2|Hypoglycemia, unspecified
C0020617|ICD9CM|AB|251.0|Hypoglycemic coma
C0020617|ICD9CM|PT|251.0|Hypoglycemic coma
C0020621|ICD9CM|AB|276.8|Hypopotassemia
C0020621|ICD9CM|PT|276.8|Hypopotassemia
C0020623|ICD9CM|AB|272.5|Lipoprotein deficiencies
C0020623|ICD9CM|PT|272.5|Lipoprotein deficiencies
C0020626|ICD9CM|AB|252.1|Hypoparathyroidism
C0020626|ICD9CM|PT|252.1|Hypoparathyroidism
C0020632|ICD9CM|HT|07.6|Hypophysectomy
C0020632|ICD9CM|PT|07.69|Total excision of pituitary gland, unspecified approach
C0020632|ICD9CM|AB|07.69|Total exc pituitary NOS
C0020641|ICD9CM|AB|364.05|Hypopyon
C0020641|ICD9CM|PT|364.05|Hypopyon
C0020645|ICD9CM|PT|276.1|Hyposmolality and/or hyponatremia
C0020645|ICD9CM|AB|276.1|Hyposmolality
C0020649|ICD9CM|HT|458|Hypotension
C0020649|ICD9CM|AB|458.9|Hypotension NOS
C0020649|ICD9CM|PT|458.9|Hypotension, unspecified
C0020651|ICD9CM|AB|458.0|Orthostatic hypotension
C0020651|ICD9CM|PT|458.0|Orthostatic hypotension
C0020673|ICD9CM|PT|99.81|Hypothermia (central) (local)
C0020673|ICD9CM|AB|99.81|Hypothermia
C0020676|ICD9CM|AB|244.9|Hypothyroidism NOS
C0020676|ICD9CM|PT|244.9|Unspecified acquired hypothyroidism
C0020700|ICD9CM|HT|68.5|Vaginal hysterectomy
C0020701|ICD9CM|AB|300.10|Hysteria NOS
C0020701|ICD9CM|PT|300.10|Hysteria, unspecified
C0020703|ICD9CM|AB|300.13|Dissociative fugue
C0020703|ICD9CM|PT|300.13|Dissociative fugue
C0020708|ICD9CM|PT|69.41|Suture of laceration of uterus
C0020708|ICD9CM|AB|69.41|Suture uterine lacerat
C0020710|ICD9CM|AB|68.12|Hysteroscopy
C0020710|ICD9CM|PT|68.12|Hysteroscopy
C0020711|ICD9CM|AB|68.0|Hysterotomy
C0020711|ICD9CM|PT|68.0|Hysterotomy
C0020748|ICD9CM|AB|E003.1|Ice hockey
C0020748|ICD9CM|PT|E003.1|Activities involving ice hockey
C0020749|ICD9CM|AB|E003.0|Ice Skating
C0020749|ICD9CM|PT|E003.0|Activities involving ice skating
C0020758|ICD9CM|AB|757.1|Ichthyosis congenita
C0020758|ICD9CM|PT|757.1|Ichthyosis congenita
C0020795|ICD9CM|AB|313.82|Identity disorder
C0020795|ICD9CM|PT|313.82|Identity disorder of childhood or adolescence
C0020807|ICD9CM|PT|516.1|Idiopathic pulmonary hemosiderosis
C0020807|ICD9CM|AB|516.1|Idio pulm hemosiderosis
C0020883|ICD9CM|HT|46.2|Ileostomy
C0020883|ICD9CM|AB|46.20|Ileostomy NOS
C0020883|ICD9CM|PT|46.20|Ileostomy, not otherwise specified
C0020941|ICD9CM|AB|991.4|Immersion foot
C0020941|ICD9CM|PT|991.4|Immersion foot
C0021051|ICD9CM|PT|279.3|Unspecified immunity deficiency
C0021051|ICD9CM|AB|279.3|Immunity deficiency NOS
C0021092|ICD9CM|AB|380.4|Impacted cerumen
C0021092|ICD9CM|PT|380.4|Impacted cerumen
C0021099|ICD9CM|AB|684|Impetigo
C0021099|ICD9CM|PT|684|Impetigo
C0021109|ICD9CM|PT|20.96|Implantation or replacement of cochlear prosthetic device, not otherwise specified
C0021109|ICD9CM|AB|20.96|Implt cochlear prost NOS
C0021122|ICD9CM|PT|312.30|Impulse control disorder, unspecified
C0021122|ICD9CM|AB|312.30|Impulse control dis NOS
C0021138|ICD9CM|PT|V60.2|Inadequate material resources
C0021138|ICD9CM|AB|V60.2|Economic problem
C0021192|ICD9CM|AB|030.2|Indeterminate leprosy
C0021192|ICD9CM|PT|030.2|Indeterminate leprosy [group I]
C0021193|ICD9CM|PT|752.7|Indeterminate sex and pseudohermaphroditism
C0021193|ICD9CM|AB|752.7|Indeterminate sex
C0021293|ICD9CM|AB|766.21|Post-term infant
C0021293|ICD9CM|PT|766.21|Post-term infant
C0021313|ICD9CM|HT|590|Infections of kidney
C0021313|ICD9CM|AB|590.9|Infection of kidney NOS
C0021313|ICD9CM|PT|590.9|Infection of kidney, unspecified
C0021345|ICD9CM|AB|075|Infectious mononucleosis
C0021345|ICD9CM|PT|075|Infectious mononucleosis
C0021355|ICD9CM|HT|380.1|Infective otitis externa
C0021355|ICD9CM|PT|380.10|Infective otitis externa, unspecified
C0021355|ICD9CM|AB|380.10|Infec otitis externa NOS
C0021360|ICD9CM|PT|606.8|Infertility due to extratesticular causes
C0021360|ICD9CM|AB|606.8|Male infertility NEC
C0021361|ICD9CM|HT|628|Infertility, female
C0021361|ICD9CM|AB|628.9|Female infertility NOS
C0021361|ICD9CM|PT|628.9|Infertility, female, of unspecified origin
C0021362|ICD9CM|PT|628.8|Infertility, female, of other specified origin
C0021362|ICD9CM|AB|628.8|Female infertility NEC
C0021364|ICD9CM|HT|606|Infertility, male
C0021364|ICD9CM|AB|606.9|Male infertility NOS
C0021364|ICD9CM|PT|606.9|Male infertility, unspecified
C0021396|ICD9CM|PT|720.81|Inflammatory spondylopathies in diseases classified elsewhere
C0021396|ICD9CM|AB|720.81|Spondylopathy in oth dis
C0021400|ICD9CM|HT|487|Influenza
C0021414|ICD9CM|PT|487.1|Influenza with other respiratory manifestations
C0021414|ICD9CM|AB|487.1|Flu w resp manifest NEC
C0021447|ICD9CM|HT|550.9|Inguinal hernia, without mention of obstruction or gangrene
C0021482|ICD9CM|PT|39.92|Injection of sclerosing agent into vein
C0021482|ICD9CM|AB|39.92|Vein inject-scleros agnt
C0021498|ICD9CM|PT|03.92|Injection of other agent into spinal canal
C0021498|ICD9CM|AB|03.92|Spinal canal inject NEC
C0021505|ICD9CM|PT|862.0|Injury to diaphragm, without mention of open wound into cavity
C0021505|ICD9CM|AB|862.0|Diaphragm injury-closed
C0021567|ICD9CM|PT|919.4|Insect bite, nonvenomous, of other, multiple, and unspecified sites, without mention of infection
C0021567|ICD9CM|AB|919.4|Insect bite NEC
C0021587|ICD9CM|AB|69.92|Artificial insemination
C0021587|ICD9CM|PT|69.92|Artificial insemination
C0021607|ICD9CM|PT|327.00|Organic insomnia, unspecified
C0021607|ICD9CM|AB|327.00|Organic insomnia NOS
C0021614|ICD9CM|AB|798.1|Instantaneous death
C0021614|ICD9CM|PT|798.1|Instantaneous death
C0021705|ICD9CM|PT|94.01|Administration of intelligence test
C0021705|ICD9CM|AB|94.01|Intelligence test admin
C0021776|ICD9CM|PT|312.34|Intermittent explosive disorder
C0021776|ICD9CM|AB|312.34|Intermitt explosive dis
C0021777|ICD9CM|AB|93.91|Ippb
C0021777|ICD9CM|PT|93.91|Intermittent positive pressure breathing [IPPB]
C0021779|ICD9CM|PT|869.0|Internal injury to unspecified or ill-defined organs without mention of open wound into cavity
C0021779|ICD9CM|AB|869.0|Internal inj NOS-closed
C0021781|ICD9CM|PT|36.15|Single internal mammary-coronary artery bypass
C0021781|ICD9CM|AB|36.15|1 int mam-cor art bypass
C0021816|ICD9CM|PT|80.52|Intervertebral chemonucleolysis
C0021816|ICD9CM|AB|80.52|Chemonucleolysis iv disc
C0021830|ICD9CM|PT|271.3|Intestinal disaccharidase deficiencies and disaccharide malabsorption
C0021830|ICD9CM|AB|271.3|Disaccharidase def/malab
C0021831|ICD9CM|PT|569.9|Unspecified disorder of intestine
C0021831|ICD9CM|AB|569.9|Intestinal disorder NOS
C0021832|ICD9CM|PT|129|Intestinal parasitism, unspecified
C0021832|ICD9CM|AB|129|Intestin parasitism NOS
C0021843|ICD9CM|PT|560.9|Unspecified intestinal obstruction
C0021843|ICD9CM|AB|560.9|Intestinal obstruct NOS
C0021844|ICD9CM|HT|560|Intestinal obstruction without mention of hernia
C0021845|ICD9CM|AB|569.83|Perforation of intestine
C0021845|ICD9CM|PT|569.83|Perforation of intestine
C0021859|ICD9CM|PT|39.1|Intra-abdominal venous shunt
C0021859|ICD9CM|AB|39.1|Intra-abd venous shunt
C0021874|ICD9CM|AB|324.0|Intracranial abscess
C0021874|ICD9CM|PT|324.0|Intracranial abscess
C0021878|ICD9CM|HT|854.0|Intracranial injury of other and unspecified nature without mention of open intracranial wound
C0021879|ICD9CM|PT|854.00|Intracranial injury of other and unspecified nature without mention of open intracranial wound, unspecified state of consciousness
C0021879|ICD9CM|AB|854.00|Brain injury NEC
C0021932|ICD9CM|PT|96.04|Insertion of endotracheal tube
C0021932|ICD9CM|AB|96.04|Insert endotracheal tube
C0021933|ICD9CM|AB|560.0|Intussusception
C0021933|ICD9CM|PT|560.0|Intussusception
C0022024|ICD9CM|AB|99.27|Iontophoresis
C0022024|ICD9CM|PT|99.27|Iontophoresis
C0022073|ICD9CM|AB|364.3|Iridocyclitis NOS
C0022073|ICD9CM|PT|364.3|Unspecified iridocyclitis
C0022102|ICD9CM|AB|96.51|Irrigation of eye
C0022102|ICD9CM|PT|96.51|Irrigation of eye
C0022104|ICD9CM|AB|564.1|Irritable bowel syndrome
C0022104|ICD9CM|PT|564.1|Irritable bowel syndrome
C0022107|ICD9CM|AB|799.22|Irritability
C0022107|ICD9CM|PT|799.22|Irritability
C0022336|ICD9CM|HT|046.1|Jakob-Creutzfeldt disease
C0022362|ICD9CM|HT|526|Diseases of the jaws
C0022362|ICD9CM|AB|526.9|Jaw disease NOS
C0022362|ICD9CM|PT|526.9|Unspecified disease of the jaws
C0022408|ICD9CM|AB|719.90|Joint dis NOS-unspec jt
C0022408|ICD9CM|HT|716.9|Arthropathy, unspecified
C0022408|ICD9CM|HT|719.9|Unspecified disorder of joint
C0022408|ICD9CM|PT|716.90|Arthropathy, unspecified, site unspecified
C0022408|ICD9CM|PT|719.90|Unspecified disorder of joint, site unspecified
C0022408|ICD9CM|AB|716.90|Arthropathy NOS-unspec
C0022411|ICD9CM|HT|718.1|Loose body in joint
C0022411|ICD9CM|AB|718.10|Loose body-unspec
C0022411|ICD9CM|PT|718.10|Loose body in joint, site unspecified
C0022548|ICD9CM|AB|701.4|Keloid scar
C0022548|ICD9CM|PT|701.4|Keloid scar
C0022568|ICD9CM|HT|370|Keratitis
C0022568|ICD9CM|AB|370.9|Keratitis NOS
C0022568|ICD9CM|PT|370.9|Unspecified keratitis
C0022570|ICD9CM|AB|054.42|Dendritic keratitis
C0022570|ICD9CM|PT|054.42|Dendritic keratitis
C0022573|ICD9CM|AB|370.40|Keratoconjunctivitis NOS
C0022573|ICD9CM|PT|370.40|Keratoconjunctivitis, unspecified
C0022578|ICD9CM|HT|371.6|Keratoconus
C0022578|ICD9CM|AB|371.60|Keratoconus NOS
C0022578|ICD9CM|PT|371.60|Keratoconus, unspecified
C0022581|ICD9CM|AB|701.1|Keratoderma, acquired
C0022581|ICD9CM|PT|701.1|Keratoderma, acquired
C0022602|ICD9CM|AB|702.0|Actinic keratosis
C0022602|ICD9CM|PT|702.0|Actinic keratosis
C0022603|ICD9CM|HT|702.1|Seborrheic keratosis
C0022607|ICD9CM|AB|11.75|Radial keratotomy
C0022607|ICD9CM|PT|11.75|Radial keratotomy
C0022650|ICD9CM|AB|592.0|Calculus of kidney
C0022650|ICD9CM|PT|592.0|Calculus of kidney
C0022660|ICD9CM|HT|584|Acute kidney failure
C0022660|ICD9CM|AB|584.9|Acute kidney failure NOS
C0022660|ICD9CM|PT|584.9|Acute kidney failure, unspecified
C0022661|ICD9CM|AB|585.6|End stage renal disease
C0022661|ICD9CM|PT|585.6|End stage renal disease
C0022671|ICD9CM|HT|55.6|Transplant of kidney
C0022680|ICD9CM|AB|753.12|Polycystic kidney NOS
C0022680|ICD9CM|PT|753.12|Polycystic kidney, unspecified type
C0022681|ICD9CM|AB|753.17|Medullary sponge kidney
C0022681|ICD9CM|PT|753.17|Medullary sponge kidney
C0022734|ICD9CM|AB|312.32|Kleptomania
C0022734|ICD9CM|PT|312.32|Kleptomania
C0022735|ICD9CM|AB|758.7|Klinefelter's syndrome
C0022735|ICD9CM|PT|758.7|Klinefelter's syndrome
C0022738|ICD9CM|PT|756.16|Klippel-Feil syndrome
C0022738|ICD9CM|AB|756.16|Klippel-feil syndrome
C0022782|ICD9CM|AB|607.0|Leukoplakia of penis
C0022782|ICD9CM|PT|607.0|Leukoplakia of penis
C0022802|ICD9CM|AB|046.0|Kuru
C0022802|ICD9CM|PT|046.0|Kuru
C0022806|ICD9CM|AB|260|Kwashiorkor
C0022806|ICD9CM|PT|260|Kwashiorkor
C0022810|ICD9CM|AB|065.2|Kyasanur forest disease
C0022810|ICD9CM|PT|065.2|Kyasanur forest disease
C0022820|ICD9CM|HT|737.3|Kyphoscoliosis and scoliosis
C0022822|ICD9CM|HT|737.1|Kyphosis (acquired)
C0022823|ICD9CM|PT|737.10|Kyphosis (acquired) (postural)
C0022823|ICD9CM|AB|737.10|Kyphosis NOS
C0022893|ICD9CM|HT|386.3|Labyrinthitis
C0022893|ICD9CM|AB|386.30|Labyrinthitis NOS
C0022893|ICD9CM|PT|386.30|Labyrinthitis, unspecified
C0022904|ICD9CM|HT|375|Disorders of lacrimal system
C0022904|ICD9CM|PT|375.9|Unspecified disorder of lacrimal system
C0022904|ICD9CM|AB|375.9|Lacrimal syst dis NOS
C0022927|ICD9CM|HT|676.9|Unspecified disorder of lactation
C0022927|ICD9CM|PT|676.90|Unspecified disorder of lactation, unspecified as to episode of care or not applicable
C0022927|ICD9CM|AB|676.90|Lactation dis NOS-unspec
C0022972|ICD9CM|HT|358.3|Lambert-Eaton syndrome
C0023035|ICD9CM|HT|54.6|Suture of abdominal wall and peritoneum
C0023038|ICD9CM|HT|54.1|Laparotomy
C0023051|ICD9CM|PT|478.70|Unspecified disease of larynx
C0023051|ICD9CM|AB|478.70|Disease of larynx NOS
C0023052|ICD9CM|AB|478.6|Edema of larynx
C0023052|ICD9CM|PT|478.6|Edema of larynx
C0023065|ICD9CM|HT|30|Excision of larynx
C0023066|ICD9CM|AB|478.75|Laryngeal spasm
C0023066|ICD9CM|PT|478.75|Laryngeal spasm
C0023071|ICD9CM|PT|31.61|Suture of laceration of larynx
C0023071|ICD9CM|AB|31.61|Suture of laryngeal lac
C0023073|ICD9CM|PT|31.42|Laryngoscopy and other tracheoscopy
C0023073|ICD9CM|AB|31.42|Larygnoscopy/tracheoscop
C0023075|ICD9CM|AB|478.74|Stenosis of larynx
C0023075|ICD9CM|PT|478.74|Stenosis of larynx
C0023105|ICD9CM|HT|295.5|Latent schizophrenia
C0023105|ICD9CM|PT|295.50|Latent schizophrenia, unspecified
C0023105|ICD9CM|AB|295.50|Latent schizophren-unsp
C0023176|ICD9CM|PT|984.9|Toxic effect of unspecified lead compound
C0023176|ICD9CM|HT|984|Toxic effect of lead and its compounds (including fumes)
C0023176|ICD9CM|AB|984.9|Tox eff lead compnd NOS
C0023212|ICD9CM|AB|428.1|Left heart failure
C0023212|ICD9CM|PT|428.1|Left heart failure
C0023241|ICD9CM|AB|482.84|Legionnaires' disease
C0023241|ICD9CM|PT|482.84|Pneumonia due to Legionnaires' disease
C0023281|ICD9CM|HT|085|Leishmaniasis
C0023281|ICD9CM|AB|085.9|Leishmaniasis NOS
C0023281|ICD9CM|PT|085.9|Leishmaniasis, unspecified
C0023285|ICD9CM|PT|085.2|Cutaneous leishmaniasis, Asian desert
C0023285|ICD9CM|AB|085.2|Cutan leishmanias asian
C0023290|ICD9CM|AB|085.0|Visceral leishmaniasis
C0023290|ICD9CM|PT|085.0|Visceral [kala-azar] leishmaniasis
C0023311|ICD9CM|HT|13.7|Insertion of prosthetic lens [pseudophakos]
C0023311|ICD9CM|PT|13.70|Insertion of pseudophakos, not otherwise specified
C0023311|ICD9CM|AB|13.70|Insert pseudophakos NOS
C0023316|ICD9CM|AB|379.32|Subluxation of lens
C0023316|ICD9CM|PT|379.32|Subluxation of lens
C0023343|ICD9CM|HT|030|Leprosy
C0023343|ICD9CM|AB|030.9|Leprosy NOS
C0023343|ICD9CM|PT|030.9|Leprosy, unspecified
C0023346|ICD9CM|AB|030.3|Borderline leprosy
C0023346|ICD9CM|PT|030.3|Borderline leprosy [group B]
C0023348|ICD9CM|AB|030.0|Lepromatous leprosy
C0023348|ICD9CM|PT|030.0|Lepromatous leprosy [type L]
C0023351|ICD9CM|AB|030.1|Tuberculoid leprosy
C0023351|ICD9CM|PT|030.1|Tuberculoid leprosy [type T]
C0023364|ICD9CM|HT|100|Leptospirosis
C0023364|ICD9CM|AB|100.9|Leptospirosis NOS
C0023364|ICD9CM|PT|100.9|Leptospirosis, unspecified
C0023370|ICD9CM|PT|444.01|Saddle embolus of abdominal aorta
C0023370|ICD9CM|AB|444.01|Saddle embolus abd aorta
C0023381|ICD9CM|HT|202.5|Letterer-Siwe disease
C0023416|ICD9CM|PT|99.72|Therapeutic leukopheresis
C0023416|ICD9CM|AB|99.72|Therapeutc leukopheresis
C0023418|ICD9CM|HT|208|Leukemia of unspecified cell type
C0023418|ICD9CM|HT|208.9|Unspecified leukemia
C0023434|ICD9CM|HT|204.1|Lymphoid leukemia, chronic
C0023443|ICD9CM|HT|202.4|Leukemic reticuloendotheliosis
C0023448|ICD9CM|HT|204|Lymphoid leukemia
C0023448|ICD9CM|HT|204.9|Unspecified lymphoid leukemia
C0023449|ICD9CM|HT|204.0|Lymphoid leukemia, acute
C0023462|ICD9CM|HT|207.2|Megakaryocytic leukemia
C0023465|ICD9CM|HT|206.0|Monocytic leukemia, acute
C0023466|ICD9CM|HT|206.1|Monocytic leukemia, chronic
C0023467|ICD9CM|HT|205.0|Myeloid leukemia, acute
C0023470|ICD9CM|HT|205|Myeloid leukemia
C0023470|ICD9CM|HT|205.9|Unspecified myeloid leukemia
C0023473|ICD9CM|HT|205.1|Myeloid leukemia, chronic
C0023484|ICD9CM|HT|203.1|Plasma cell leukemia
C0023501|ICD9CM|PT|288.62|Leukemoid reaction
C0023501|ICD9CM|AB|288.62|Leukemoid reaction
C0023510|ICD9CM|HT|288|Diseases of white blood cells
C0023510|ICD9CM|PT|288.9|Unspecified disease of white blood cells
C0023510|ICD9CM|AB|288.9|Wbc disease NOS
C0023518|ICD9CM|AB|288.60|Leukocytosis NOS
C0023518|ICD9CM|PT|288.60|Leukocytosis, unspecified
C0023520|ICD9CM|AB|330.0|Leukodystrophy
C0023520|ICD9CM|PT|330.0|Leukodystrophy
C0023524|ICD9CM|PT|046.3|Progressive multifocal leukoencephalopathy
C0023524|ICD9CM|AB|046.3|Prog multifoc leukoencep
C0023529|ICD9CM|PT|779.7|Periventricular leukomalacia
C0023529|ICD9CM|AB|779.7|Perivent leukomalacia
C0023530|ICD9CM|AB|288.50|Leukocytopenia NOS
C0023530|ICD9CM|PT|288.50|Leukocytopenia, unspecified
C0023534|ICD9CM|PT|623.5|Leukorrhea, not specified as infective
C0023534|ICD9CM|AB|623.5|Noninfect vag leukorrhea
C0023643|ICD9CM|PT|697.9|Lichen, unspecified
C0023643|ICD9CM|HT|697|Lichen
C0023643|ICD9CM|AB|697.9|Lichen NOS
C0023646|ICD9CM|AB|697.0|Lichen planus
C0023646|ICD9CM|PT|697.0|Lichen planus
C0023654|ICD9CM|PT|698.3|Lichenification and lichen simplex chronicus
C0023654|ICD9CM|AB|698.3|Lichenification
C0023702|ICD9CM|AB|994.0|Effects of lightning
C0023702|ICD9CM|PT|994.0|Effects of lightning
C0023760|ICD9CM|AB|528.5|Diseases of lips
C0023760|ICD9CM|PT|528.5|Diseases of lips
C0023787|ICD9CM|AB|272.6|Lipodystrophy
C0023787|ICD9CM|PT|272.6|Lipodystrophy
C0023788|ICD9CM|AB|040.2|Whipple's disease
C0023788|ICD9CM|PT|040.2|Whipple's disease
C0023794|ICD9CM|AB|272.7|Lipidoses
C0023794|ICD9CM|PT|272.7|Lipidoses
C0023798|ICD9CM|HT|214|Lipoma
C0023798|ICD9CM|AB|214.9|Lipoma NOS
C0023798|ICD9CM|PT|214.9|Lipoma, unspecified site
C0023800|ICD9CM|PT|214.8|Lipoma of other specified sites
C0023800|ICD9CM|AB|214.8|Lipoma NEC
C0023817|ICD9CM|AB|272.3|Hyperchylomicronemia
C0023817|ICD9CM|PT|272.3|Hyperchylomicronemia
C0023860|ICD9CM|AB|027.0|Listeriosis
C0023860|ICD9CM|PT|027.0|Listeriosis
C0023885|ICD9CM|AB|572.0|Abscess of liver
C0023885|ICD9CM|PT|572.0|Abscess of liver
C0023886|ICD9CM|AB|006.3|Amebic liver abscess
C0023886|ICD9CM|PT|006.3|Amebic liver abscess
C0023891|ICD9CM|PT|571.2|Alcoholic cirrhosis of liver
C0023891|ICD9CM|AB|571.2|Alcohol cirrhosis liver
C0023892|ICD9CM|AB|571.6|Biliary cirrhosis
C0023892|ICD9CM|PT|571.6|Biliary cirrhosis
C0023895|ICD9CM|PT|573.9|Unspecified disorder of liver
C0023895|ICD9CM|AB|573.9|Liver disorder NOS
C0023908|ICD9CM|PT|V42.7|Liver replaced by transplant
C0023908|ICD9CM|AB|V42.7|Liver transplant status
C0023911|ICD9CM|HT|50.5|Liver transplant
C0023944|ICD9CM|AB|344.81|Locked-in state
C0023944|ICD9CM|PT|344.81|Locked-in state
C0023968|ICD9CM|AB|125.2|Loiasis
C0023968|ICD9CM|PT|125.2|Loiasis
C0023976|ICD9CM|AB|426.82|Long QT syndrome
C0023976|ICD9CM|PT|426.82|Long QT syndrome
C0023985|ICD9CM|AB|46.22|Continent ileostomy
C0023985|ICD9CM|PT|46.22|Continent ileostomy
C0023988|ICD9CM|PT|718.18|Loose body in joint, other specified sites
C0023988|ICD9CM|AB|718.18|Loose body-joint NEC
C0024004|ICD9CM|HT|737.2|Lordosis (acquired)
C0024005|ICD9CM|AB|737.20|Lordosis NOS
C0024005|ICD9CM|PT|737.20|Lordosis (acquired) (postural)
C0024025|ICD9CM|AB|063.1|Louping ill
C0024025|ICD9CM|PT|063.1|Louping ill
C0024031|ICD9CM|AB|724.2|Lumbago
C0024031|ICD9CM|PT|724.2|Lumbago
C0024054|ICD9CM|PT|426.81|Lown-Ganong-Levine syndrome
C0024054|ICD9CM|AB|426.81|Lown-ganong-levine synd
C0024103|ICD9CM|AB|611.72|Lump or mass in breast
C0024103|ICD9CM|PT|611.72|Lump or mass in breast
C0024110|ICD9CM|AB|513.0|Abscess of lung
C0024110|ICD9CM|PT|513.0|Abscess of lung
C0024128|ICD9CM|HT|33.5|Lung transplant
C0024128|ICD9CM|AB|33.50|Lung transplant NOS
C0024128|ICD9CM|PT|33.50|Lung transplantation, not otherwise specified
C0024141|ICD9CM|PT|710.0|Systemic lupus erythematosus
C0024141|ICD9CM|AB|710.0|Syst lupus erythematosus
C0024198|ICD9CM|PT|088.81|Lyme Disease
C0024198|ICD9CM|AB|088.81|Lyme disease
C0024207|ICD9CM|PT|289.3|Lymphadenitis, unspecified, except mesenteric
C0024207|ICD9CM|AB|289.3|Lymphadenitis NOS
C0024221|ICD9CM|AB|228.1|Lymphangioma, any site
C0024221|ICD9CM|PT|228.1|Lymphangioma, any site
C0024225|ICD9CM|AB|457.2|Lymphangitis
C0024225|ICD9CM|PT|457.2|Lymphangitis
C0024286|ICD9CM|AB|099.1|Lymphogranuloma venereum
C0024286|ICD9CM|PT|099.1|Lymphogranuloma venereum
C0024301|ICD9CM|HT|202.0|Nodular lymphoma
C0024302|ICD9CM|HT|200.0|Reticulosarcoma
C0024302|ICD9CM|HT|200.7|Large cell lymphoma
C0024312|ICD9CM|PT|288.51|Lymphocytopenia
C0024312|ICD9CM|AB|288.51|Lymphocytopenia
C0024419|ICD9CM|AB|273.3|Macroglobulinemia
C0024419|ICD9CM|PT|273.3|Macroglobulinemia
C0024433|ICD9CM|AB|744.83|Macrostomia
C0024433|ICD9CM|PT|744.83|Macrostomia
C0024439|ICD9CM|PT|371.55|Macular corneal dystrophy
C0024439|ICD9CM|AB|371.55|Macular cornea dystrophy
C0024486|ICD9CM|PT|88.97|Magnetic resonance imaging of other and unspecified sites
C0024486|ICD9CM|AB|88.97|Magnetic res image unsp
C0024508|ICD9CM|HT|524.0|Major anomalies of jaw size
C0024508|ICD9CM|PT|524.00|Major anomalies of jaw size, unspecified anomaly
C0024508|ICD9CM|AB|524.00|Unspcf anomaly jaw size
C0024517|ICD9CM|HT|296.2|Major depressive disorder, single episode
C0024517|ICD9CM|PT|296.20|Major depressive affective disorder, single episode, unspecified
C0024517|ICD9CM|AB|296.20|Depress psychosis-unspec
C0024523|ICD9CM|PT|579.9|Unspecified intestinal malabsorption
C0024523|ICD9CM|HT|579|Intestinal malabsorption
C0024523|ICD9CM|AB|579.9|Intest malabsorption NOS
C0024528|ICD9CM|HT|780.7|Malaise and fatigue
C0024530|ICD9CM|HT|084|Malaria
C0024530|ICD9CM|AB|084.6|Malaria NOS
C0024530|ICD9CM|PT|084.6|Malaria, unspecified
C0024535|ICD9CM|AB|084.0|Falciparum malaria
C0024535|ICD9CM|PT|084.0|Falciparum malaria [malignant tertian]
C0024536|ICD9CM|AB|084.2|Quartan malaria
C0024536|ICD9CM|PT|084.2|Quartan malaria
C0024537|ICD9CM|AB|084.1|Vivax malaria
C0024537|ICD9CM|PT|084.1|Vivax malaria [benign tertian]
C0024559|ICD9CM|AB|63.70|Male sterilization NOS
C0024559|ICD9CM|PT|63.70|Male sterilization procedure, not otherwise specified
C0024586|ICD9CM|AB|259.2|Carcinoid syndrome
C0024586|ICD9CM|PT|259.2|Carcinoid syndrome
C0024588|ICD9CM|PT|401.0|Malignant essential hypertension
C0024588|ICD9CM|AB|401.0|Malignant hypertension
C0024591|ICD9CM|AB|995.86|Malignant hyperthermia
C0024591|ICD9CM|PT|995.86|Malignant hyperthermia
C0024620|ICD9CM|PT|155.0|Malignant neoplasm of liver, primary
C0024620|ICD9CM|AB|155.0|Mal neo liver, primary
C0024621|ICD9CM|PT|174.0|Malignant neoplasm of nipple and areola of female breast
C0024621|ICD9CM|AB|174.0|Malig neo nipple
C0024622|ICD9CM|PT|190.5|Malignant neoplasm of retina
C0024622|ICD9CM|AB|190.5|Malign neopl retina
C0024623|ICD9CM|HT|151|Malignant neoplasm of stomach
C0024623|ICD9CM|PT|151.9|Malignant neoplasm of stomach, unspecified site
C0024623|ICD9CM|AB|151.9|Malig neopl stomach NOS
C0024624|ICD9CM|PT|162.3|Malignant neoplasm of upper lobe, bronchus or lung
C0024624|ICD9CM|AB|162.3|Mal neo upper lobe lung
C0024633|ICD9CM|AB|530.7|Mallory-weiss syndrome
C0024633|ICD9CM|PT|530.7|Gastroesophageal laceration-hemorrhage syndrome
C0024636|ICD9CM|AB|524.4|Malocclusion NOS
C0024636|ICD9CM|PT|524.4|Malocclusion, unspecified
C0024649|ICD9CM|PT|746.87|Malposition of heart and cardiac apex
C0024649|ICD9CM|AB|746.87|Malposition of heart
C0024713|ICD9CM|PT|296.40|Bipolar I disorder, most recent episode (or current) manic, unspecified
C0024713|ICD9CM|AB|296.40|Bipol I currnt manic NOS
C0024796|ICD9CM|AB|759.82|Marfan syndrome
C0024796|ICD9CM|PT|759.82|Marfan syndrome
C0024881|ICD9CM|HT|85.4|Mastectomy
C0024885|ICD9CM|AB|85.23|Subtotal mastectomy
C0024885|ICD9CM|PT|85.23|Subtotal mastectomy
C0024886|ICD9CM|PT|85.41|Unilateral simple mastectomy
C0024886|ICD9CM|AB|85.41|Unilat simple mastectomy
C0024902|ICD9CM|AB|611.71|Mastodynia
C0024902|ICD9CM|PT|611.71|Mastodynia
C0024904|ICD9CM|AB|383.9|Mastoiditis NOS
C0024904|ICD9CM|PT|383.9|Unspecified mastoiditis
C0025007|ICD9CM|HT|055|Measles
C0025037|ICD9CM|AB|751.0|Meckel's diverticulum
C0025037|ICD9CM|PT|751.0|Meckel's diverticulum
C0025064|ICD9CM|AB|519.2|Mediastinitis
C0025064|ICD9CM|PT|519.2|Mediastinitis
C0025065|ICD9CM|AB|34.22|Mediastinoscopy
C0025065|ICD9CM|PT|34.22|Mediastinoscopy
C0025229|ICD9CM|AB|025|Melioidosis
C0025229|ICD9CM|PT|025|Melioidosis
C0025267|ICD9CM|AB|258.01|Mult endo neoplas type I
C0025267|ICD9CM|PT|258.01|Multiple endocrine neoplasia [MEN] type I
C0025268|ICD9CM|AB|258.02|Mult endo neop type IIA
C0025268|ICD9CM|PT|258.02|Multiple endocrine neoplasia [MEN] type IIA
C0025269|ICD9CM|AB|258.03|Mult endo neop type IIB
C0025269|ICD9CM|PT|258.03|Multiple endocrine neoplasia [MEN] type IIB
C0025281|ICD9CM|HT|386.0|Meniere's disease
C0025281|ICD9CM|AB|386.00|Meniere's disease NOS
C0025281|ICD9CM|PT|386.00|Ménière's disease, unspecified
C0025287|ICD9CM|AB|781.6|Meningismus
C0025287|ICD9CM|PT|781.6|Meningismus
C0025289|ICD9CM|AB|322.9|Meningitis NOS
C0025289|ICD9CM|HT|322|Meningitis of unspecified cause
C0025289|ICD9CM|PT|322.9|Meningitis, unspecified
C0025292|ICD9CM|AB|320.0|Hemophilus meningitis
C0025292|ICD9CM|PT|320.0|Hemophilus meningitis
C0025294|ICD9CM|AB|036.0|Meningococcal meningitis
C0025294|ICD9CM|PT|036.0|Meningococcal meningitis
C0025295|ICD9CM|AB|320.1|Pneumococcal meningitis
C0025295|ICD9CM|PT|320.1|Pneumococcal meningitis
C0025297|ICD9CM|AB|047.9|Viral meningitis NOS
C0025297|ICD9CM|PT|047.9|Unspecified viral meningitis
C0025303|ICD9CM|HT|036|Meningococcal infection
C0025303|ICD9CM|PT|036.9|Meningococcal infection, unspecified
C0025303|ICD9CM|AB|036.9|Meningococcal infect NOS
C0025306|ICD9CM|AB|036.2|Meningococcemia
C0025306|ICD9CM|PT|036.2|Meningococcemia
C0025322|ICD9CM|AB|256.31|Premature menopause
C0025322|ICD9CM|PT|256.31|Premature menopause
C0025335|ICD9CM|PT|69.6|Menstrual extraction or regulation
C0025335|ICD9CM|AB|69.6|Menstrual extraction
C0025427|ICD9CM|PT|985.0|Toxic effect of mercury and its compounds
C0025427|ICD9CM|AB|985.0|Toxic effect mercury
C0025469|ICD9CM|AB|289.2|Mesenteric lymphadenitis
C0025469|ICD9CM|PT|289.2|Nonspecific mesenteric lymphadenitis
C0025517|ICD9CM|PT|277.9|Unspecified disorder of metabolism
C0025517|ICD9CM|AB|277.9|Metabolism disorder NOS
C0025530|ICD9CM|AB|121.5|Metagonimiasis
C0025530|ICD9CM|PT|121.5|Metagonimiasis
C0025637|ICD9CM|AB|289.7|Methemoglobinemia
C0025637|ICD9CM|PT|289.7|Methemoglobinemia
C0025874|ICD9CM|AB|626.6|Metrorrhagia
C0025874|ICD9CM|PT|626.6|Metrorrhagia
C0025958|ICD9CM|AB|742.1|Microcephalus
C0025958|ICD9CM|PT|742.1|Microcephalus
C0025988|ICD9CM|AB|750.16|Microglossia
C0025988|ICD9CM|PT|750.16|Microglossia
C0025990|ICD9CM|AB|524.04|Mandibular hypoplasia
C0025990|ICD9CM|PT|524.04|Major anomalies of jaw size, mandibular hypoplasia
C0026010|ICD9CM|HT|743.1|Microphthalmos
C0026010|ICD9CM|AB|743.10|Microphthalmos NOS
C0026010|ICD9CM|AB|743.11|Simple microphthalmos
C0026010|ICD9CM|PT|743.11|Simple microphthalmos
C0026010|ICD9CM|PT|743.10|Microphthalmos, unspecified
C0026034|ICD9CM|AB|744.84|Microstomia
C0026034|ICD9CM|PT|744.84|Microstomia
C0026106|ICD9CM|PT|317|Mild intellectual disabilities
C0026106|ICD9CM|AB|317|Mild intellect disabilty
C0026143|ICD9CM|AB|051.9|Paravaccinia NOS
C0026143|ICD9CM|AB|051.1|Pseudocowpox
C0026143|ICD9CM|PT|051.1|Pseudocowpox
C0026143|ICD9CM|PT|051.9|Paravaccinia, unspecified
C0026205|ICD9CM|PT|379.42|Miosis (persistent), not due to miotics
C0026205|ICD9CM|AB|379.42|Miosis not d/t miotics
C0026229|ICD9CM|HT|133|Acariasis
C0026229|ICD9CM|AB|133.9|Acariasis NOS
C0026229|ICD9CM|PT|133.9|Acariasis, unspecified
C0026265|ICD9CM|AB|424.0|Mitral valve disorder
C0026265|ICD9CM|PT|424.0|Mitral valve disorders
C0026351|ICD9CM|PT|318.0|Moderate intellectual disabilities
C0026351|ICD9CM|AB|318.0|Mod intellect disability
C0026393|ICD9CM|AB|078.0|Molluscum contagiosum
C0026393|ICD9CM|PT|078.0|Molluscum contagiosum
C0026471|ICD9CM|PT|273.1|Monoclonal paraproteinemia
C0026471|ICD9CM|AB|273.1|Monoclon paraproteinemia
C0026509|ICD9CM|PT|813.03|Closed Monteggia's fracture
C0026509|ICD9CM|AB|813.03|Monteggia's fx-closed
C0026603|ICD9CM|AB|994.6|Motion sickness
C0026603|ICD9CM|PT|994.6|Motion sickness
C0026614|ICD9CM|HT|E819|Motor vehicle traffic accident of unspecified nature
C0026618|ICD9CM|AB|520.3|Mottled teeth
C0026618|ICD9CM|PT|520.3|Mottled teeth
C0026654|ICD9CM|AB|437.5|Moyamoya disease
C0026654|ICD9CM|PT|437.5|Moyamoya disease
C0026686|ICD9CM|PT|527.6|Mucocele of salivary gland
C0026686|ICD9CM|AB|527.6|Salivary gland mucocele
C0026691|ICD9CM|PT|446.1|Acute febrile mucocutaneous lymph node syndrome [MCLS]
C0026691|ICD9CM|AB|446.1|Mucocutan lymph node syn
C0026703|ICD9CM|AB|277.5|Mucopolysaccharidosis
C0026703|ICD9CM|PT|277.5|Mucopolysaccharidosis
C0026725|ICD9CM|AB|622.7|Mucous polyp of cervix
C0026725|ICD9CM|PT|622.7|Mucous polyp of cervix
C0026758|ICD9CM|PT|759.7|Multiple congenital anomalies, so described
C0026758|ICD9CM|AB|759.7|Mult congen anomal NEC
C0026760|ICD9CM|PT|756.56|Multiple epiphyseal dysplasia
C0026760|ICD9CM|AB|756.56|Mult epiphyseal dysplas
C0026764|ICD9CM|HT|203.0|Multiple myeloma
C0026769|ICD9CM|AB|340|Multiple sclerosis
C0026769|ICD9CM|PT|340|Multiple sclerosis
C0026773|ICD9CM|PT|300.14|Dissociative identity disorder
C0026773|ICD9CM|AB|300.14|Dissociatve identity dis
C0026780|ICD9CM|HT|072|Mumps
C0026847|ICD9CM|HT|335.1|Spinal muscular atrophy
C0026847|ICD9CM|PT|335.10|Spinal muscular atrophy, unspecified
C0026847|ICD9CM|AB|335.10|Spinal muscl atrophy NOS
C0026848|ICD9CM|AB|359.9|Myopathy NOS
C0026848|ICD9CM|PT|359.9|Myopathy, unspecified
C0026849|ICD9CM|HT|359|Muscular dystrophies and other myopathies
C0026868|ICD9CM|AB|93.84|Music therapy
C0026868|ICD9CM|PT|93.84|Music therapy
C0026893|ICD9CM|PT|729.1|Myalgia and myositis, unspecified
C0026893|ICD9CM|AB|729.1|Myalgia and myositis NOS
C0026896|ICD9CM|HT|358.0|Myasthenia gravis
C0026897|ICD9CM|PT|358.1|Myasthenic syndromes in diseases classified elsewhere
C0026897|ICD9CM|AB|358.1|Myasthenia in oth dis
C0026918|ICD9CM|PT|031.9|Unspecified diseases due to mycobacteria
C0026918|ICD9CM|AB|031.9|Mycobacterial dis NOS
C0026946|ICD9CM|HT|110-118.99|MYCOSES
C0026948|ICD9CM|HT|202.1|Mycosis fungoides
C0026962|ICD9CM|PT|379.43|Mydriasis (persistent), not due to mydriatics
C0026962|ICD9CM|AB|379.43|Mydriasis not d/t mydrtc
C0026987|ICD9CM|PT|289.83|Myelofibrosis
C0026987|ICD9CM|AB|289.83|Myelofibrosis
C0026995|ICD9CM|AB|87.21|Contrast myelogram
C0026995|ICD9CM|PT|87.21|Contrast myelogram
C0027030|ICD9CM|AB|134.0|Myiasis
C0027030|ICD9CM|PT|134.0|Myiasis
C0027046|ICD9CM|AB|429.1|Myocardial degeneration
C0027046|ICD9CM|PT|429.1|Myocardial degeneration
C0027059|ICD9CM|AB|429.0|Myocarditis NOS
C0027059|ICD9CM|PT|429.0|Myocarditis, unspecified
C0027066|ICD9CM|AB|333.2|Myoclonus
C0027066|ICD9CM|PT|333.2|Myoclonus
C0027080|ICD9CM|AB|791.3|Myoglobinuria
C0027080|ICD9CM|PT|791.3|Myoglobinuria
C0027092|ICD9CM|AB|367.1|Myopia
C0027092|ICD9CM|PT|367.1|Myopia
C0027126|ICD9CM|PT|359.21|Myotonic muscular dystrophy
C0027126|ICD9CM|AB|359.21|Myotonic musclr dystrphy
C0027127|ICD9CM|PT|359.22|Myotonia congenita
C0027127|ICD9CM|AB|359.22|Myotonia congenita
C0027128|ICD9CM|AB|366.43|Myotonic cataract
C0027128|ICD9CM|PT|366.43|Myotonic cataract
C0027136|ICD9CM|AB|19.4|Myringoplasty
C0027136|ICD9CM|PT|19.4|Myringoplasty
C0027339|ICD9CM|HT|703|Diseases of nail
C0027339|ICD9CM|AB|703.9|Disease of nail NOS
C0027339|ICD9CM|PT|703.9|Unspecified disease of nail
C0027343|ICD9CM|AB|703.0|Ingrowing nail
C0027343|ICD9CM|PT|703.0|Ingrowing nail
C0027402|ICD9CM|PT|301.81|Narcissistic personality disorder
C0027402|ICD9CM|AB|301.81|Narcissistic personality
C0027404|ICD9CM|HT|347.0|Narcolepsy
C0027430|ICD9CM|HT|471|Nasal polyps
C0027430|ICD9CM|AB|471.9|Nasal polyp NOS
C0027430|ICD9CM|PT|471.9|Unspecified nasal polyp
C0027430|ICD9CM|AB|471.0|Polyp of nasal cavity
C0027430|ICD9CM|PT|471.0|Polyp of nasal cavity
C0027450|HL7V3.0|CSY|ICD9CMDiagnosiscodes|National Center for Health Statistics
C0027450|HL7V3.0|CSY|ICD9CMProcedurecodes|National Center for Health Statistics
C0027498|ICD9CM|HT|787.0|Nausea and vomiting
C0027498|ICD9CM|AB|787.01|Nausea with vomiting
C0027498|ICD9CM|PT|787.01|Nausea with vomiting
C0027529|ICD9CM|AB|126.1|Necator Americanus
C0027529|ICD9CM|PT|126.1|Necatoriasis due to necator americanus
C0027535|ICD9CM|AB|847.0|Sprain of neck
C0027535|ICD9CM|PT|847.0|Sprain of neck
C0027537|ICD9CM|AB|040.3|Necrobacillosis
C0027537|ICD9CM|PT|040.3|Necrobacillosis
C0027609|ICD9CM|PT|779.5|Drug withdrawal syndrome in newborn
C0027609|ICD9CM|AB|779.5|NB drug withdrawal syndr
C0027611|ICD9CM|PT|771.6|Neonatal conjunctivitis and dacryocystitis
C0027611|ICD9CM|AB|771.6|Neonatal conjunctivitis
C0027630|ICD9CM|PT|238.0|Neoplasm of uncertain behavior of bone and articular cartilage
C0027630|ICD9CM|AB|238.0|Unc behav neo bone
C0027632|ICD9CM|HT|238.7|Neoplasm of uncertain behavior of other lymphatic and hematopoietic tissues
C0027634|ICD9CM|PT|237.3|Neoplasm of uncertain behavior of paraganglia
C0027634|ICD9CM|AB|237.3|Unc behav neo paragang
C0027636|ICD9CM|PT|237.0|Neoplasm of uncertain behavior of pituitary gland and craniopharyngeal duct
C0027636|ICD9CM|AB|237.0|Unc behav neo pituitary
C0027638|ICD9CM|PT|238.6|Neoplasm of uncertain behavior of plasma cells
C0027638|ICD9CM|AB|238.6|Plasmacytoma NOS
C0027639|ICD9CM|PT|239.4|Neoplasm of unspecified nature of bladder
C0027639|ICD9CM|AB|239.4|Bladder neoplasm NOS
C0027641|ICD9CM|AB|239.3|Breast neoplasm NOS
C0027641|ICD9CM|PT|239.3|Neoplasm of unspecified nature of breast
C0027651|ICD9CM|HT|140-239.99|NEOPLASMS
C0027698|ICD9CM|HT|583|Nephritis and nephropathy, not specified as acute or chronic
C0027699|ICD9CM|PT|583.81|Nephritis and nephropathy, not specified as acute or chronic, in diseases classified elsewhere
C0027699|ICD9CM|AB|583.81|Nephritis NOS in oth dis
C0027700|ICD9CM|PT|583.2|Nephritis and nephropathy, not specified as acute or chronic, with lesion of membranoproliferative glomerulonephritis
C0027700|ICD9CM|AB|583.2|Membranoprolif nephr NOS
C0027701|ICD9CM|PT|583.1|Nephritis and nephropathy, not specified as acute or chronic, with lesion of membranous glomerulonephritis
C0027701|ICD9CM|AB|583.1|Membranous nephritis NOS
C0027702|MTH|PN|NOCODE|Nephritis NEC in ICD9CM_2014
C0027702|ICD9CM|HT|583.8|Nephritis and nephropathy, not specified as acute or chronic, with other specified pathological lesion in kidney
C0027702|ICD9CM|PT|583.89|Nephritis and nephropathy, not specified as acute or chronic, with other specified pathological lesion in kidney
C0027702|ICD9CM|AB|583.89|Nephritis NEC
C0027703|ICD9CM|PT|583.9|Nephritis and nephropathy, not specified as acute or chronic, with unspecified pathological lesion in kidney
C0027703|ICD9CM|AB|583.9|Nephritis NOS
C0027719|ICD9CM|AB|587|Renal sclerosis NOS
C0027719|ICD9CM|PT|587|Renal sclerosis, unspecified
C0027726|ICD9CM|HT|581|Nephrotic syndrome
C0027729|ICD9CM|HT|581.8|Nephrotic syndrome with other specified pathological lesion in kidney
C0027729|ICD9CM|PT|581.89|Nephrotic syndrome with other specified pathological lesion in kidney
C0027729|ICD9CM|AB|581.89|Nephrotic syndrome NEC
C0027730|ICD9CM|PT|581.9|Nephrotic syndrome with unspecified pathological lesion in kidney
C0027730|ICD9CM|AB|581.9|Nephrotic syndrome NOS
C0027732|ICD9CM|AB|55.51|Nephroureterectomy
C0027732|ICD9CM|PT|55.51|Nephroureterectomy
C0027765|ICD9CM|PT|349.9|Unspecified disorders of nervous system
C0027765|ICD9CM|AB|349.9|Cns disorder NOS
C0027769|ICD9CM|AB|799.21|Nervousness
C0027769|ICD9CM|PT|799.21|Nervousness
C0027804|ICD9CM|AB|300.5|Neurasthenia
C0027804|ICD9CM|PT|300.5|Neurasthenia
C0027821|ICD9CM|PT|306.2|Cardiovascular malfunction arising from mental factors
C0027821|ICD9CM|AB|306.2|Psychogen cardiovasc dis
C0027831|ICD9CM|PT|237.71|Neurofibromatosis, type 1 [von recklinghausen's disease]
C0027831|ICD9CM|AB|237.71|Neurofibromatosis type I
C0027832|ICD9CM|PT|237.72|Neurofibromatosis, type 2 [acoustic neurofibromatosis]
C0027832|ICD9CM|AB|237.72|Neurofibromatosis typ II
C0027849|ICD9CM|PT|333.92|Neuroleptic malignant syndrome
C0027849|ICD9CM|AB|333.92|Neuroleptic malgnt synd
C0027853|ICD9CM|AB|89.13|Neurologic examination
C0027853|ICD9CM|PT|89.13|Neurologic examination
C0027868|ICD9CM|HT|358|Myoneural disorders
C0027868|ICD9CM|AB|358.9|Myoneural disorders NOS
C0027868|ICD9CM|PT|358.9|Myoneural disorders, unspecified
C0027873|ICD9CM|AB|341.0|Neuromyelitis optica
C0027873|ICD9CM|PT|341.0|Neuromyelitis optica
C0027927|ICD9CM|HT|094|Neurosyphilis
C0027927|ICD9CM|AB|094.9|Neurosyphilis NOS
C0027927|ICD9CM|PT|094.9|Neurosyphilis, unspecified
C0027947|ICD9CM|HT|288.0|Neutropenia
C0027947|ICD9CM|AB|288.00|Neutropenia NOS
C0027947|ICD9CM|PT|288.00|Neutropenia, unspecified
C0028077|ICD9CM|HT|368.6|Night blindness
C0028077|ICD9CM|AB|368.60|Night blindness NOS
C0028077|ICD9CM|PT|368.60|Night blindness, unspecified
C0028271|ICD9CM|AB|528.1|Cancrum oris
C0028271|ICD9CM|PT|528.1|Cancrum oris
C0028283|ICD9CM|HT|283.1|Non-autoimmune hemolytic anemias
C0028283|ICD9CM|PT|283.10|Non-autoimmune hemolytic anemia, unspecified
C0028283|ICD9CM|AB|283.10|Nonauto hem anemia NOS
C0028315|ICD9CM|HT|793.9|Nonspecific abnormal findings on radiological and other examination of other sites of body
C0028431|ICD9CM|PT|738.0|Acquired deformity of nose
C0028431|ICD9CM|AB|738.0|Acq nose deformity
C0028734|ICD9CM|AB|788.43|Nocturia
C0028734|ICD9CM|PT|788.43|Nocturia
C0028738|ICD9CM|AB|379.50|Nystagmus NOS
C0028738|ICD9CM|PT|379.50|Nystagmus, unspecified
C0028754|ICD9CM|AB|278.00|Obesity NOS
C0028754|ICD9CM|PT|278.00|Obesity, unspecified
C0028756|ICD9CM|AB|278.01|Morbid obesity
C0028756|ICD9CM|PT|278.01|Morbid obesity
C0028768|ICD9CM|PT|300.3|Obsessive-compulsive disorders
C0028768|ICD9CM|AB|300.3|Obsessive-compulsive dis
C0028790|ICD9CM|HT|434|Occlusion of cerebral arteries
C0028790|ICD9CM|HT|434.9|Cerebral artery occlusion, unspecified
C0028840|ICD9CM|AB|365.04|Ocular hypertension
C0028840|ICD9CM|PT|365.04|Ocular hypertension
C0028841|ICD9CM|HT|360.3|Hypotony of eye
C0028841|ICD9CM|AB|360.30|Hypotony NOS, eye
C0028841|ICD9CM|PT|360.30|Hypotony of eye, unspecified
C0028850|ICD9CM|PT|378.9|Unspecified disorder of eye movements
C0028850|ICD9CM|AB|378.9|Eye movemnt disorder NOS
C0028856|ICD9CM|AB|781.93|Ocular torticollis
C0028856|ICD9CM|PT|781.93|Ocular torticollis
C0028960|ICD9CM|AB|606.1|Oligospermia
C0028960|ICD9CM|PT|606.1|Oligospermia
C0028962|ICD9CM|PT|788.5|Oliguria and anuria
C0028962|ICD9CM|AB|788.5|Oliguria & anuria
C0029001|ICD9CM|AB|125.3|Onchocerciasis
C0029001|ICD9CM|PT|125.3|Onchocerciasis
C0029077|ICD9CM|AB|360.11|Sympathetic uveitis
C0029077|ICD9CM|PT|360.11|Sympathetic uveitis
C0029090|ICD9CM|AB|16.21|Ophthalmoscopy
C0029090|ICD9CM|PT|16.21|Ophthalmoscopy
C0029095|ICD9CM|HT|305.5|Opioid abuse
C0029106|ICD9CM|AB|121.0|Opisthorchiasis
C0029106|ICD9CM|PT|121.0|Opisthorchiasis
C0029119|ICD9CM|AB|118|Opportunistic mycoses
C0029119|ICD9CM|PT|118|Opportunistic mycoses
C0029121|ICD9CM|PT|313.81|Oppositional defiant disorder
C0029121|ICD9CM|AB|313.81|Opposition defiant disor
C0029124|ICD9CM|HT|377.1|Optic atrophy
C0029124|ICD9CM|AB|377.10|Optic atrophy NOS
C0029124|ICD9CM|PT|377.10|Optic atrophy, unspecified
C0029125|ICD9CM|AB|377.16|Hereditary optic atrophy
C0029125|ICD9CM|PT|377.16|Hereditary optic atrophy
C0029128|ICD9CM|AB|377.21|Drusen of optic disc
C0029128|ICD9CM|PT|377.21|Drusen of optic disc
C0029134|ICD9CM|HT|377.3|Optic neuritis
C0029134|ICD9CM|AB|377.30|Optic neuritis NOS
C0029134|ICD9CM|PT|377.30|Optic neuritis, unspecified
C0029171|ICD9CM|PT|528.8|Oral submucosal fibrosis, including of tongue
C0029171|ICD9CM|AB|528.8|Oral submucosal fibrosis
C0029182|ICD9CM|PT|376.9|Unspecified disorder of orbit
C0029182|ICD9CM|HT|376|Disorders of the orbit
C0029182|ICD9CM|AB|376.9|Orbital disorder NOS
C0029188|ICD9CM|PT|62.61|Suture of laceration of testis
C0029188|ICD9CM|AB|62.61|Suture testicular lacer
C0029226|ICD9CM|PT|293.82|Psychotic disorder with hallucinations in conditions classified elsewhere
C0029226|ICD9CM|AB|293.82|Psy dis w halluc oth dis
C0029291|ICD9CM|HT|073|Ornithosis
C0029291|ICD9CM|AB|073.9|Ornithosis NOS
C0029291|ICD9CM|PT|073.9|Ornithosis, unspecified
C0029336|ICD9CM|AB|V58.5|Orthodontics aftercare
C0029336|ICD9CM|PT|V58.5|Orthodontics aftercare
C0029402|ICD9CM|HT|731|Osteitis deformans and osteopathies associated with other disorders classified elsewhere
C0029403|ICD9CM|PT|731.0|Osteitis deformans without mention of bone tumor
C0029403|ICD9CM|AB|731.0|Osteitis deformans NOS
C0029408|ICD9CM|HT|715.9|Osteoarthrosis, unspecified whether generalized or localized
C0029412|ICD9CM|AB|731.2|Hypertroph osteoarthrop
C0029412|ICD9CM|PT|731.2|Hypertrophic pulmonary osteoarthropathy
C0029421|ICD9CM|PT|732.7|Osteochondritis dissecans
C0029421|ICD9CM|AB|732.7|Osteochondrit dissecans
C0029434|ICD9CM|AB|756.51|Osteogenesis imperfecta
C0029434|ICD9CM|PT|756.51|Osteogenesis imperfecta
C0029442|ICD9CM|AB|268.2|Osteomalacia NOS
C0029442|ICD9CM|PT|268.2|Osteomalacia, unspecified
C0029443|ICD9CM|HT|730.2|Unspecified osteomyelitis
C0029443|ICD9CM|PT|730.20|Unspecified osteomyelitis, site unspecified
C0029443|ICD9CM|AB|730.20|Osteomyelitis NOS-unspec
C0029454|ICD9CM|AB|756.52|Osteopetrosis
C0029454|ICD9CM|PT|756.52|Osteopetrosis
C0029455|ICD9CM|AB|756.53|Osteopoikilosis
C0029455|ICD9CM|PT|756.53|Osteopoikilosis
C0029456|ICD9CM|HT|733.0|Osteoporosis
C0029456|ICD9CM|AB|733.00|Osteoporosis NOS
C0029456|ICD9CM|PT|733.00|Osteoporosis, unspecified
C0029459|ICD9CM|AB|733.01|Senile osteoporosis
C0029459|ICD9CM|PT|733.01|Senile osteoporosis
C0029480|ICD9CM|PT|39.29|Other (peripheral) vascular shunt or bypass
C0029480|ICD9CM|AB|39.29|Vasc shunt & bypass NEC
C0029481|ICD9CM|PT|790.6|Other abnormal blood chemistry
C0029481|ICD9CM|AB|790.6|Abn blood chemistry NEC
C0029482|ICD9CM|PT|133.8|Other acariasis
C0029482|ICD9CM|AB|133.8|Acariasis NEC
C0029483|ICD9CM|PT|E910.8|Other accidental drowning or submersion
C0029483|ICD9CM|AB|E910.8|Accidental drowning NEC
C0029484|ICD9CM|PT|E928.8|Other accidents
C0029484|ICD9CM|HT|E916-E928.9|OTHER ACCIDENTS
C0029484|ICD9CM|AB|E928.8|Accident NEC
C0029485|ICD9CM|PT|706.1|Other acne
C0029485|ICD9CM|AB|706.1|Acne NEC
C0029486|ICD9CM|PT|736.89|Other acquired deformity of other parts of limb
C0029486|ICD9CM|AB|736.89|Oth acq limb deformity
C0029487|ICD9CM|AB|99.92|Other acupuncture
C0029487|ICD9CM|PT|99.92|Other acupuncture
C0029488|ICD9CM|PT|308.3|Other acute reactions to stress
C0029488|ICD9CM|AB|308.3|Acute stress react NEC
C0029489|ICD9CM|PT|704.09|Other alopecia
C0029489|ICD9CM|AB|704.09|Alopecia NEC
C0029490|ICD9CM|HT|848|Other and ill-defined sprains and strains
C0029493|ICD9CM|PT|253.1|Other and unspecified anterior pituitary hyperfunction
C0029493|ICD9CM|AB|253.1|Ant pituit hyperfunc NEC
C0029495|ICD9CM|PT|245.8|Other and unspecified chronic thyroiditis
C0029495|ICD9CM|AB|245.8|Chr thyroiditis NEC/NOS
C0029496|ICD9CM|PT|286.9|Other and unspecified coagulation defects
C0029496|ICD9CM|AB|286.9|Coagulat defect NEC/NOS
C0029497|ICD9CM|PT|722.90|Other and unspecified disc disorder, unspecified region
C0029497|ICD9CM|AB|722.90|Disc dis NEC/NOS-unspec
C0029498|ICD9CM|PT|528.9|Other and unspecified diseases of the oral soft tissues
C0029498|ICD9CM|AB|528.9|Oral soft tissue dis NEC
C0029499|ICD9CM|PT|993.2|Other and unspecified effects of high altitude
C0029499|ICD9CM|AB|993.2|Eff high altitud NEC/NOS
C0029500|ICD9CM|HT|E928|Other and unspecified environmental and accidental causes
C0029505|ICD9CM|PT|959.4|Hand, except finger injury
C0029505|ICD9CM|AB|959.4|Hand injury NOS
C0029506|ICD9CM|PT|959.7|Knee, leg, ankle, and foot injury
C0029506|ICD9CM|AB|959.7|Lower leg injury NOS
C0029507|ICD9CM|PT|959.8|Other specified sites, including multiple injury
C0029507|ICD9CM|AB|959.8|Injury mlt site/site NEC
C0029508|ICD9CM|HT|959.1|Other and unspecified injury to trunk
C0029509|ICD9CM|PT|959.9|Unspecified site injury
C0029509|ICD9CM|AB|959.9|Injury-site NOS
C0029510|ICD9CM|PT|265.1|Other and unspecified manifestations of thiamine deficiency
C0029510|ICD9CM|AB|265.1|Thiamine defic NEC/NOS
C0029511|ICD9CM|PT|117.9|Other and unspecified mycoses
C0029511|ICD9CM|AB|117.9|Mycoses NEC & NOS
C0029512|ICD9CM|HT|558|Other and unspecified noninfectious gastroenteritis and colitis
C0029512|ICD9CM|PT|558.9|Other and unspecified noninfectious gastroenteritis and colitis
C0029512|ICD9CM|AB|558.9|Noninf gastroenterit NEC
C0029513|ICD9CM|PT|620.2|Other and unspecified ovarian cyst
C0029513|ICD9CM|AB|620.2|Ovarian cyst NEC/NOS
C0029514|ICD9CM|PT|696.5|Other and unspecified pityriasis
C0029514|ICD9CM|AB|696.5|Pityriasis NEC & NOS
C0029515|ICD9CM|PT|579.3|Other and unspecified postsurgical nonabsorption
C0029515|ICD9CM|AB|579.3|Intest postop nonabsorb
C0029516|ICD9CM|PT|298.8|Other and unspecified reactive psychosis
C0029516|ICD9CM|AB|298.8|React psychosis NEC/NOS
C0029519|ICD9CM|PT|414.19|Other aneurysm of heart
C0029519|ICD9CM|AB|414.19|Aneurysm of heart NEC
C0029520|ICD9CM|PT|747.49|Other anomalies of great veins
C0029520|ICD9CM|AB|747.49|Great vein anomaly NEC
C0029522|ICD9CM|PT|95.46|Other auditory and vestibular function tests
C0029522|ICD9CM|AB|95.46|Audit & vestib test NEC
C0029523|ICD9CM|PT|266.2|Other B-complex deficiencies
C0029523|ICD9CM|AB|266.2|B-complex defic NEC
C0029524|ICD9CM|HT|66.3|Other bilateral destruction or occlusion of fallopian tubes
C0029524|ICD9CM|PT|66.39|Other bilateral destruction or occlusion of fallopian tubes
C0029524|ICD9CM|AB|66.39|Bilat tubal destruct NEC
C0029525|ICD9CM|PT|733.29|Other bone cyst
C0029525|ICD9CM|AB|733.29|Bone cyst NEC
C0029526|ICD9CM|AB|33.23|Other bronchoscopy
C0029526|ICD9CM|PT|33.23|Other bronchoscopy
C0029527|ICD9CM|PT|023.8|Other brucellosis
C0029527|ICD9CM|AB|023.8|Brucellosis NEC
C0029528|ICD9CM|PT|727.3|Other bursitis
C0029528|ICD9CM|AB|727.3|Bursitis NEC
C0029531|ICD9CM|PT|366.8|Other cataract
C0029531|ICD9CM|AB|366.8|Cataract NEC
C0029534|ICD9CM|PT|334.3|Other cerebellar ataxia
C0029534|ICD9CM|AB|334.3|Cerebellar ataxia NEC
C0029535|ICD9CM|PT|74.99|Other cesarean section of unspecified type
C0029535|ICD9CM|AB|74.99|Cesarean section NOS
C0029537|ICD9CM|PT|786.59|Other chest pain
C0029537|ICD9CM|AB|786.59|Chest pain NEC
C0029538|ICD9CM|PT|87.54|Other cholangiogram
C0029538|ICD9CM|AB|87.54|Cholangiogram NEC
C0029539|ICD9CM|HT|575.1|Other cholecystitis
C0029540|MTH|PN|NOCODE|Cholecystostomy NEC in ICD9CM_2014
C0029540|ICD9CM|PT|51.03|Other cholecystostomy
C0029540|ICD9CM|AB|51.03|Cholecystostomy NEC
C0029541|ICD9CM|AB|03.29|Other chordotomy
C0029541|ICD9CM|PT|03.29|Other chordotomy
C0029542|ICD9CM|PT|333.5|Other choreas
C0029542|ICD9CM|AB|333.5|Chorea NEC
C0029543|ICD9CM|PT|372.14|Other chronic allergic conjunctivitis
C0029543|ICD9CM|AB|372.14|Chr allrg conjunctiv NEC
C0029544|ICD9CM|PT|491.8|Other chronic bronchitis
C0029544|ICD9CM|AB|491.8|Chronic bronchitis NEC
C0029545|ICD9CM|PT|571.49|Other chronic hepatitis
C0029545|ICD9CM|AB|571.49|Chronic hepatitis NEC
C0029546|ICD9CM|PT|571.8|Other chronic nonalcoholic liver disease
C0029546|ICD9CM|AB|571.8|Chronic liver dis NEC
C0029547|ICD9CM|HT|803.0|Other closed skull fracture without mention of intracranial injury
C0029548|ICD9CM|PT|368.59|Other color vision deficiencies
C0029548|ICD9CM|AB|368.59|Color deficiency NEC
C0029549|ICD9CM|PT|758.5|Other conditions due to autosomal anomalies
C0029549|ICD9CM|AB|758.5|Autosomal anomalies NEC
C0029550|ICD9CM|PT|758.81|Other conditions due to sex chromosome anomalies
C0029550|ICD9CM|AB|758.81|Oth cond due to sex chrm
C0029551|ICD9CM|HT|348.8|Other conditions of brain
C0029551|ICD9CM|HT|348|Other conditions of brain
C0029552|ICD9CM|PT|743.49|Other congenital anomalies of anterior segment
C0029552|ICD9CM|AB|743.49|Anom anter seg NEC-eye
C0029553|ICD9CM|PT|752.49|Other anomalies of cervix, vagina, and external female genitalia
C0029553|ICD9CM|AB|752.49|Cervix/fem gen anom NEC
C0029554|ICD9CM|PT|751.69|Other anomalies of gallbladder, bile ducts, and liver
C0029554|ICD9CM|AB|751.69|Biliary & liver anom NEC
C0029557|ICD9CM|PT|755.63|Other congenital deformity of hip (joint)
C0029557|ICD9CM|AB|755.63|Cong hip deformity NEC
C0029559|ICD9CM|PT|756.59|Other osteodystrophies
C0029559|ICD9CM|AB|756.59|Osteodystrophy NEC
C0029560|ICD9CM|PT|372.39|Other conjunctivitis
C0029560|ICD9CM|AB|372.39|Conjunctivitis NEC
C0029560|ICD9CM|HT|372.3|Other and unspecified conjunctivitis
C0029561|ICD9CM|PT|87.32|Other contrast bronchogram
C0029561|ICD9CM|AB|87.32|Contrast bronchogram NEC
C0029562|ICD9CM|PT|87.02|Other contrast radiogram of brain and skull
C0029562|ICD9CM|AB|87.02|Brain/skull contrst xray
C0029563|ICD9CM|PT|11.69|Other corneal transplant
C0029563|ICD9CM|AB|11.69|Corneal transplant NEC
C0029565|ICD9CM|PT|94.49|Other counseling
C0029565|ICD9CM|AB|94.49|Other counselling
C0029566|ICD9CM|AB|01.24|Other craniotomy
C0029566|ICD9CM|PT|01.24|Other craniotomy
C0029568|ICD9CM|PT|57.32|Other cystoscopy
C0029568|ICD9CM|AB|57.32|Cystoscopy NEC
C0029569|ICD9CM|PT|526.2|Other cysts of jaws
C0029569|ICD9CM|AB|526.2|Cysts of jaws NEC
C0029570|ICD9CM|PT|277.6|Other deficiencies of circulating enzymes
C0029570|ICD9CM|AB|277.6|Defic circul enzyme NEC
C0029571|ICD9CM|PT|333.0|Other degenerative diseases of the basal ganglia
C0029571|ICD9CM|AB|333.0|Degen basal ganglia NEC
C0029572|ICD9CM|PT|87.12|Other dental x-ray
C0029572|ICD9CM|AB|87.12|Dental x-ray NEC
C0029574|ICD9CM|HT|702|Other dermatoses
C0029575|ICD9CM|PT|V21.2|Other development of adolescence
C0029575|ICD9CM|AB|V21.2|Adolescence growth NEC
C0029577|ICD9CM|PT|12.29|Other diagnostic procedures on iris, ciliary body, sclera, and anterior chamber
C0029577|ICD9CM|AB|12.29|Ant segment dx proc NEC
C0029579|MTH|PN|NOCODE|OTHER LUNG DISEASE NEC in ICD9CM
C0029579|ICD9CM|PT|518.89|Other diseases of lung, not elsewhere classified
C0029579|ICD9CM|AB|518.89|Other lung disease NEC
C0029581|ICD9CM|PT|478.19|Other disease of nasal cavity and sinuses
C0029581|ICD9CM|HT|478.1|Other diseases of nasal cavity and sinuses
C0029581|ICD9CM|AB|478.19|Nasal & sinus dis NEC
C0029582|ICD9CM|HT|519|Other diseases of respiratory system
C0029582|ICD9CM|HT|510-519.99|OTHER DISEASES OF RESPIRATORY SYSTEM
C0029586|ICD9CM|HT|733|Other disorders of bone and cartilage
C0029586|ICD9CM|PT|733.99|Other disorders of bone and cartilage
C0029586|ICD9CM|HT|733.9|Other and unspecified disorders of bone and cartilage
C0029586|ICD9CM|AB|733.99|Bone & cartilage dis NEC
C0029587|ICD9CM|PT|307.59|Other disorders of eating
C0029587|ICD9CM|AB|307.59|Eating disorder NEC
C0029587|ICD9CM|HT|307.5|Other and unspecified disorders of eating
C0029588|ICD9CM|PT|312.39|Other disorders of impulse control
C0029588|ICD9CM|AB|312.39|Impulse control dis NEC
C0029590|ICD9CM|PT|379.39|Other disorders of lens
C0029590|ICD9CM|AB|379.39|Disorders of lens NEC
C0029591|ICD9CM|PT|272.8|Other disorders of lipoid metabolism
C0029591|ICD9CM|AB|272.8|Lipoid metabol dis NEC
C0029592|ICD9CM|PT|626.8|Other disorders of menstruation and other abnormal bleeding from female genital tract
C0029592|ICD9CM|AB|626.8|Menstrual disorder NEC
C0029593|ICD9CM|PT|253.6|Other disorders of neurohypophysis
C0029593|ICD9CM|AB|253.6|Neurohypophysis dis NEC
C0029594|ICD9CM|PT|273.8|Other disorders of plasma protein metabolism
C0029594|ICD9CM|AB|273.8|Dis plas protein met NEC
C0029595|ICD9CM|PT|277.2|Other disorders of purine and pyrimidine metabolism
C0029595|ICD9CM|AB|277.2|Purine/pyrimid dis NEC
C0029596|ICD9CM|HT|367.8|Other disorders of refraction and accommodation
C0029596|ICD9CM|PT|367.89|Other disorders of refraction and accommodation
C0029596|ICD9CM|AB|367.89|Refraction disorder NEC
C0029597|ICD9CM|PT|253.8|Other disorders of the pituitary and other syndromes of diencephalohypophyseal origin
C0029597|ICD9CM|AB|253.8|Pituitary disorder NEC
C0029600|ICD9CM|PT|77.39|Other division of bone, other bones
C0029600|ICD9CM|AB|77.39|Bone division NEC
C0029601|ICD9CM|PT|786.09|Other respiratory abnormalities
C0029601|ICD9CM|AB|786.09|Respiratory abnorm NEC
C0029603|ICD9CM|PT|958.8|Other early complications of trauma
C0029603|ICD9CM|AB|958.8|Early complic trauma NEC
C0029604|ICD9CM|HT|633.8|Other ectopic pregnancy
C0029605|ICD9CM|PT|99.62|Other electric countershock of heart
C0029605|ICD9CM|AB|99.62|Heart countershock NEC
C0029606|ICD9CM|PT|94.27|Other electroshock therapy
C0029606|ICD9CM|AB|94.27|Electroshock therapy NEC
C0029607|ICD9CM|PT|492.8|Other emphysema
C0029607|ICD9CM|AB|492.8|Emphysema NEC
C0029608|ICD9CM|PT|745.69|Other endocardial cushion defects
C0029608|ICD9CM|AB|745.69|Endocard cushion def NEC
C0029609|MTH|PN|NOCODE|Endocarditis NEC in ICD9CM_2014
C0029609|ICD9CM|AB|424.99|Endocarditis NEC
C0029609|ICD9CM|PT|424.99|Other endocarditis, valve unspecified
C0029610|ICD9CM|HT|360.1|Other endophthalmitis
C0029610|ICD9CM|PT|360.19|Other endophthalmitis
C0029610|ICD9CM|AB|360.19|Endophthalmitis NEC
C0029611|ICD9CM|PT|45.13|Other endoscopy of small intestine
C0029611|ICD9CM|AB|45.13|Sm bowel endoscopy NEC
C0029612|ICD9CM|HT|46.3|Other enterostomy
C0029612|ICD9CM|PT|46.39|Other enterostomy
C0029612|ICD9CM|AB|46.39|Enterostomy NEC
C0029613|ICD9CM|HT|38.6|Other excision of vessels
C0029614|ICD9CM|PT|03.09|Other exploration and decompression of spinal canal
C0029614|ICD9CM|AB|03.09|Spinal canal explor NEC
C0029616|ICD9CM|PT|351.8|Other facial nerve disorders
C0029616|ICD9CM|AB|351.8|Facial nerve dis NEC
C0029620|ICD9CM|PT|379.56|Other forms of nystagmus
C0029620|ICD9CM|AB|379.56|Nystagmus NEC
C0029622|MTH|PN|NOCODE|Gastroenterostomy NEC in ICD9CM_2014
C0029622|ICD9CM|AB|44.39|Gastroenterostomy NEC
C0029622|ICD9CM|PT|44.39|Other gastroenterostomy without gastrectomy
C0029623|MTH|PN|NOCODE|Gastroscopy NEC in ICD9CM_2014
C0029623|ICD9CM|PT|44.13|Other gastroscopy
C0029623|ICD9CM|AB|44.13|Gastroscopy NEC
C0029624|MTH|PN|NOCODE|Encounter for other specified contraceptive management in ICD9CM
C0029624|ICD9CM|PT|V25.09|Other general counseling and advice on contraceptive management
C0029624|ICD9CM|AB|V25.09|Contraceptive mangmt NEC
C0029625|ICD9CM|AB|780.99|Other general symptoms
C0029625|ICD9CM|HT|780.9|Other general symptoms
C0029625|ICD9CM|PT|780.99|Other general symptoms
C0029626|ICD9CM|PT|437.1|Other generalized ischemic cerebrovascular disease
C0029626|ICD9CM|AB|437.1|Ac cerebrovasc insuf NOS
C0029627|ICD9CM|PT|054.19|Other genital herpes
C0029627|ICD9CM|AB|054.19|Genital herpes NEC
C0029628|ICD9CM|AB|94.44|Other group therapy
C0029628|ICD9CM|PT|94.44|Other group therapy
C0029629|ICD9CM|PT|V20.1|Other healthy infant or child receiving care
C0029629|ICD9CM|AB|V20.1|Care of healthy chld NEC
C0029630|ICD9CM|AB|426.6|Other heart block
C0029630|ICD9CM|PT|426.6|Other heart block
C0029631|ICD9CM|AB|93.35|Other heat therapy
C0029631|ICD9CM|PT|93.35|Other heat therapy
C0029632|ICD9CM|PT|282.7|Other hemoglobinopathies
C0029632|ICD9CM|AB|282.7|Hemoglobinopathies NEC
C0029633|ICD9CM|PT|301.59|Other histrionic personality disorder
C0029633|ICD9CM|AB|301.59|Histrionic person NEC
C0029634|ICD9CM|AB|93.33|Other hydrotherapy
C0029634|ICD9CM|PT|93.33|Other hydrotherapy
C0029635|ICD9CM|AB|278.8|Other hyperalimentation
C0029635|ICD9CM|PT|278.8|Other hyperalimentation
C0029640|ICD9CM|PT|560.39|Other impaction of intestine
C0029640|ICD9CM|AB|560.39|Impaction intestine NEC
C0029641|ICD9CM|PT|34.09|Other incision of pleura
C0029641|ICD9CM|AB|34.09|Other pleural incision
C0029642|ICD9CM|PT|94.39|Other individual psychotherapy
C0029642|ICD9CM|AB|94.39|Individ psychotherap NEC
C0029644|ICD9CM|HT|720.8|Other inflammatory spondylopathies
C0029644|ICD9CM|PT|720.89|Other inflammatory spondylopathies
C0029644|ICD9CM|AB|720.89|Inflam spondylopathy NEC
C0029647|ICD9CM|PT|13.19|Other intracapsular extraction of lens
C0029647|ICD9CM|AB|13.19|Intracapsul lens ext NEC
C0029650|ICD9CM|PT|370.49|Other keratoconjunctivitis
C0029650|ICD9CM|AB|370.49|Keratoconjunctivitis NEC
C0029651|ICD9CM|PT|55.69|Other kidney transplantation
C0029651|ICD9CM|AB|55.69|Kidney transplant NEC
C0029652|ICD9CM|PT|737.39|Other kyphoscoliosis and scoliosis
C0029652|ICD9CM|AB|737.39|Scoliosis NEC
C0029653|ICD9CM|PT|737.19|Other kyphosis (acquired)
C0029653|ICD9CM|AB|737.19|Kyphosis NEC
C0029654|ICD9CM|PT|54.19|Other laparotomy
C0029654|ICD9CM|AB|54.19|Laparotomy NEC
C0029655|ICD9CM|HT|208.8|Other leukemia of unspecified cell type
C0029657|ICD9CM|PT|368.44|Other localized visual field defect
C0029657|ICD9CM|AB|368.44|Visual field defect NEC
C0029658|ICD9CM|PT|737.29|Other lordosis (acquired)
C0029658|ICD9CM|AB|737.29|Lordosis NEC
C0029659|ICD9CM|AB|457.1|Other lymphedema
C0029659|ICD9CM|PT|457.1|Other lymphedema
C0029660|ICD9CM|HT|204.8|Other lymphoid leukemia
C0029661|ICD9CM|PT|084.4|Other malaria
C0029661|ICD9CM|AB|084.4|Malaria NEC
C0029662|ICD9CM|HT|202.8|Other malignant lymphomas
C0029664|ICD9CM|PT|87.37|Other mammography
C0029664|ICD9CM|AB|87.37|Mammography NEC
C0029665|ICD9CM|PT|264.8|Other manifestations of vitamin A deficiency
C0029665|ICD9CM|AB|264.8|Vitamin A deficiency NEC
C0029666|ICD9CM|PT|14.74|Other mechanical vitrectomy
C0029666|ICD9CM|AB|14.74|Mech vitrectomy NEC
C0029667|ICD9CM|PT|066.3|Other mosquito-borne fever
C0029667|ICD9CM|AB|066.3|Mosquito-borne fever NEC
C0029668|ICD9CM|PT|372.03|Other mucopurulent conjunctivitis
C0029668|ICD9CM|AB|372.03|Mucopur conjunctivit NEC
C0029669|ICD9CM|HT|729.8|Other musculoskeletal symptoms referable to limbs
C0029669|ICD9CM|PT|729.89|Other musculoskeletal symptoms referable to limbs
C0029669|ICD9CM|AB|729.89|Muscskel sympt limb NEC
C0029670|ICD9CM|HT|205.8|Other myeloid leukemia
C0029672|ICD9CM|PT|368.69|Other night blindness
C0029672|ICD9CM|AB|368.69|Night blindness NEC
C0029673|ICD9CM|PT|457.8|Other noninfectious disorders of lymphatic channels
C0029673|ICD9CM|AB|457.8|Noninfect lymph dis NEC
C0029674|ICD9CM|PT|89.59|Other nonoperative cardiac and vascular measurements
C0029674|ICD9CM|AB|89.59|Nonop cardiac/vasc exam
C0029675|ICD9CM|PT|89.39|Other nonoperative measurements and examinations
C0029675|ICD9CM|AB|89.39|Nonoperative exams NEC
C0029676|ICD9CM|PT|95.49|Other nonoperative procedures related to hearing
C0029676|ICD9CM|AB|95.49|Non-op hearing proc NEC
C0029677|ICD9CM|PT|89.38|Other nonoperative respiratory measurements
C0029677|ICD9CM|AB|89.38|Respiratory measure NEC
C0029678|ICD9CM|PT|287.2|Other nonthrombocytopenic purpuras
C0029678|ICD9CM|AB|287.2|Purpura NOS
C0029679|ICD9CM|PT|537.3|Other obstruction of duodenum
C0029679|ICD9CM|AB|537.3|Duodenal obstruction NEC
C0029680|ICD9CM|HT|V62.2|Other occupational circumstances or maladjustment
C0029680|ICD9CM|PT|V62.29|Other occupational circumstances or maladjustment
C0029680|ICD9CM|AB|V62.29|Occupationl circumst NEC
C0029681|ICD9CM|PT|377.39|Other optic neuritis
C0029681|ICD9CM|AB|377.39|Optic neuritis NEC
C0029694|ICD9CM|PT|733.09|Other osteoporosis
C0029694|ICD9CM|AB|733.09|Osteoporosis NEC
C0029695|ICD9CM|HT|380.2|Other otitis externa
C0029696|ICD9CM|PT|387.8|Other otosclerosis
C0029696|ICD9CM|AB|387.8|Otosclerosis NEC
C0029697|ICD9CM|HT|256.3|Other ovarian failure
C0029697|ICD9CM|PT|256.39|Other ovarian failure
C0029697|ICD9CM|AB|256.39|Ovarian failure NEC
C0029698|ICD9CM|PT|273.2|Other paraproteinemias
C0029698|ICD9CM|AB|273.2|Paraproteinemia NEC
C0029699|ICD9CM|PT|V61.29|Other parent-child problems
C0029699|ICD9CM|AB|V61.29|Oth parent-child problem
C0029701|ICD9CM|HT|43.8|Other partial gastrectomy
C0029702|ICD9CM|HT|06.3|Other partial thyroidectomy
C0029702|ICD9CM|PT|06.39|Other partial thyroidectomy
C0029702|ICD9CM|AB|06.39|Part thyroidectomy NEC
C0029703|ICD9CM|PT|11.64|Other penetrating keratoplasty
C0029703|ICD9CM|AB|11.64|Perforat keratoplast NEC
C0029704|ICD9CM|AB|39.97|Other perfusion
C0029704|ICD9CM|PT|39.97|Other perfusion
C0029706|ICD9CM|PT|386.19|Other peripheral vertigo
C0029706|ICD9CM|HT|386.1|Other and unspecified peripheral vertigo
C0029706|ICD9CM|AB|386.19|Peripheral vertigo NEC
C0029707|ICD9CM|HT|301.8|Other personality disorders
C0029707|ICD9CM|PT|301.89|Other personality disorders
C0029707|ICD9CM|AB|301.89|Personality disorder NEC
C0029708|ICD9CM|AB|99.83|Other phototherapy
C0029708|ICD9CM|PT|99.83|Other phototherapy
C0029711|ICD9CM|PT|V50.1|Other plastic surgery for unacceptable cosmetic appearance
C0029711|ICD9CM|AB|V50.1|Plastic surgery NEC
C0029712|ICD9CM|PT|427.69|Other premature beats
C0029712|ICD9CM|AB|427.69|Premature beats NEC
C0029713|ICD9CM|HT|765.1|Other preterm infants
C0029713|ICD9CM|PT|765.10|Other preterm infants, unspecified [weight]
C0029713|ICD9CM|AB|765.10|Preterm infant NEC wtNOS
C0029715|ICD9CM|HT|658.8|Other problems associated with amniotic cavity and membranes
C0029715|ICD9CM|HT|658|Other problems associated with amniotic cavity and membranes
C0029716|MTH|PN|NOCODE|Prostatectomy NEC in ICD9CM_2014
C0029716|ICD9CM|HT|60.6|Other prostatectomy
C0029716|ICD9CM|PT|60.69|Other prostatectomy
C0029716|ICD9CM|AB|60.69|Prostatectomy NEC
C0029717|ICD9CM|PT|696.8|Other psoriasis and similar disorders
C0029717|ICD9CM|AB|696.8|Psorias related dis NEC
C0029718|ICD9CM|PT|94.29|Other psychiatric somatotherapy
C0029718|ICD9CM|AB|94.29|Psychiatr somatother NEC
C0029719|ICD9CM|PT|94.08|Other psychologic evaluation and testing
C0029719|ICD9CM|AB|94.08|Psychol eval & test NEC
C0029721|ICD9CM|PT|26.49|Other repair and plastic operations on salivary gland or duct
C0029721|ICD9CM|AB|26.49|Salivary repair NEC
C0029722|ICD9CM|HT|42.8|Other repair of esophagus
C0029722|ICD9CM|PT|42.89|Other repair of esophagus
C0029722|ICD9CM|AB|42.89|Esophageal repair NEC
C0029724|ICD9CM|HT|44.6|Other repair of stomach
C0029724|ICD9CM|PT|44.69|Other repair of stomach
C0029724|ICD9CM|AB|44.69|Gastric repair NEC
C0029725|ICD9CM|PT|39.59|Other repair of vessel
C0029725|ICD9CM|HT|39.5|Other repair of vessels
C0029725|ICD9CM|AB|39.59|Repair of vessel NEC
C0029729|ICD9CM|PT|743.56|Other retinal changes, congenital
C0029729|ICD9CM|AB|743.56|Cong retinal changes NEC
C0029730|ICD9CM|HT|398.9|Other and unspecified rheumatic heart diseases
C0029730|ICD9CM|PT|398.99|Other rheumatic heart diseases
C0029730|ICD9CM|HT|398|Other rheumatic heart disease
C0029730|ICD9CM|AB|398.99|Rheumatic heart dis NEC
C0029731|MTH|PN|NOCODE|Rhinoplasty NEC in ICD9CM_2014
C0029731|ICD9CM|PT|21.87|Other rhinoplasty
C0029731|ICD9CM|AB|21.87|Rhinoplasty NEC
C0029732|ICD9CM|PT|14.49|Other scleral buckling
C0029732|ICD9CM|AB|14.49|Scleral buckling NEC
C0029734|ICD9CM|PT|379.09|Other scleritis and episcleritis
C0029734|ICD9CM|AB|379.09|Scleritis NEC
C0029737|ICD9CM|PT|785.59|Other shock without mention of trauma
C0029737|ICD9CM|AB|785.59|Shock w/o trauma NEC
C0029739|ICD9CM|PT|86.69|Other skin graft to other sites
C0029739|ICD9CM|AB|86.69|Free skin graft NEC
C0029741|ICD9CM|PT|728.3|Other specific muscle disorders
C0029741|ICD9CM|AB|728.3|Muscle disorders NEC
C0029744|ICD9CM|PT|285.8|Other specified anemias
C0029744|ICD9CM|AB|285.8|Anemia NEC
C0029745|ICD9CM|HT|284.8|Other specified aplastic anemias
C0029746|ICD9CM|HT|716.8|Other specified arthropathy
C0029746|ICD9CM|HT|719.8|Other specified disorders of joint
C0029747|ICD9CM|PT|088.89|Other specified arthropod-borne diseases, other
C0029747|ICD9CM|HT|088.8|Other specified arthropod-borne diseases
C0029747|ICD9CM|AB|088.89|Oth arthropod-borne dis
C0029748|ICD9CM|PT|041.89|Other specified bacterial infections in conditions classified elsewhere and of unspecified site, other specified bacteria
C0029748|ICD9CM|HT|041.8|Other specified bacterial infections in conditions classified elsewhere and of unspecified site
C0029748|ICD9CM|AB|041.89|Oth specf bacteria
C0029751|ICD9CM|HT|093.8|Other specified cardiovascular syphilis
C0029751|ICD9CM|PT|093.89|Other specified cardiovascular syphilis
C0029751|ICD9CM|AB|093.89|Cardiovascular syph NEC
C0029752|ICD9CM|PT|598.8|Other specified causes of urethral stricture
C0029752|ICD9CM|AB|598.8|Urethral stricture NEC
C0029753|ICD9CM|PT|330.8|Other specified cerebral degenerations in childhood
C0029753|ICD9CM|AB|330.8|Cereb degen in child NEC
C0029754|ICD9CM|PT|123.8|Other specified cestode infection
C0029754|ICD9CM|AB|123.8|Cestode infection NEC
C0029758|ICD9CM|PT|750.4|Other specified anomalies of esophagus
C0029758|ICD9CM|AB|750.4|Esophageal anomaly NEC
C0029759|ICD9CM|PT|756.89|Other specified anomalies of muscle, tendon, fascia, and connective tissue
C0029759|ICD9CM|HT|756.8|Other specified congenital anomalies of muscle, tendon, fascia, and connective tissue
C0029759|ICD9CM|AB|756.89|Soft tissue anomaly NEC
C0029763|ICD9CM|PT|111.8|Other specified dermatomycoses
C0029763|ICD9CM|AB|111.8|Dermatomycoses NEC
C0029764|ICD9CM|HT|032.8|Other specified diphtheria
C0029764|ICD9CM|PT|032.89|Other specified diphtheria
C0029764|ICD9CM|AB|032.89|Diphtheria NEC
C0029767|ICD9CM|HT|078.8|Other specified diseases due to viruses and Chlamydiae
C0029768|ICD9CM|HT|289.8|Other specified diseases of blood and blood-forming organs
C0029768|ICD9CM|PT|289.89|Other specified diseases of blood and blood-forming organs
C0029768|ICD9CM|AB|289.89|Blood diseases NEC
C0029769|ICD9CM|PT|704.8|Other specified diseases of hair and hair follicles
C0029769|ICD9CM|AB|704.8|Hair diseases NEC
C0029770|ICD9CM|HT|521.8|Other specified diseases of hard tissues of teeth
C0029770|ICD9CM|PT|521.89|Other specific diseases of hard tissues of teeth
C0029770|ICD9CM|AB|521.89|Dis hard tiss teeth NEC
C0029771|ICD9CM|PT|577.8|Other specified diseases of pancreas
C0029771|ICD9CM|AB|577.8|Pancreatic disease NEC
C0029772|ICD9CM|HT|526.8|Other specified diseases of the jaws
C0029772|ICD9CM|PT|526.89|Other specified diseases of the jaws
C0029772|ICD9CM|AB|526.89|Jaw disease NEC
C0029773|ICD9CM|PT|527.8|Other specified diseases of the salivary glands
C0029773|ICD9CM|AB|527.8|Salivary gland dis NEC
C0029774|ICD9CM|PT|270.8|Other specified disorders of amino-acid metabolism
C0029774|ICD9CM|AB|270.8|Dis amino-acid metab NEC
C0029776|ICD9CM|PT|596.89|Other specified disorders of bladder
C0029776|ICD9CM|HT|596.8|Other specified disorders of bladder
C0029776|ICD9CM|AB|596.89|Disorders of bladder NEC
C0029777|ICD9CM|PT|271.8|Other specified disorders of carbohydrate transport and metabolism
C0029777|ICD9CM|AB|271.8|Dis carbohydr metab NEC
C0029781|ICD9CM|HT|593.8|Other specified disorders of kidney and ureter
C0029781|ICD9CM|PT|593.89|Other specified disorders of kidney and ureter
C0029781|ICD9CM|AB|593.89|Renal & ureteral dis NEC
C0029782|ICD9CM|HT|608.8|Other specified disorders of male genital organs
C0029782|ICD9CM|PT|608.89|Other specified disorders of male genital organs
C0029782|ICD9CM|AB|608.89|Male genital dis NEC
C0029784|ICD9CM|HT|349.8|Other specified disorders of nervous system
C0029784|ICD9CM|PT|349.89|Other specified disorders of nervous system
C0029784|ICD9CM|AB|349.89|Cns disorder NEC
C0029785|ICD9CM|HT|607.8|Other specified disorders of penis
C0029785|ICD9CM|PT|607.89|Other specified disorders of penis
C0029785|ICD9CM|AB|607.89|Disorder of penis NEC
C0029786|ICD9CM|HT|568.8|Other specified disorders of peritoneum
C0029786|ICD9CM|PT|568.89|Other specified disorders of peritoneum
C0029786|ICD9CM|AB|568.89|Peritoneal disorder NEC
C0029788|ICD9CM|PT|709.8|Other specified disorders of skin
C0029788|ICD9CM|AB|709.8|Skin disorders NEC
C0029790|ICD9CM|PT|525.8|Other specified disorders of the teeth and supporting structures
C0029790|ICD9CM|AB|525.8|Dental disorder NEC
C0029791|ICD9CM|HT|588.8|Other specified disorders resulting from impaired renal function
C0029791|ICD9CM|PT|588.89|Other specified disorders resulting from impaired renal function
C0029791|ICD9CM|AB|588.89|Impair ren funct dis NEC
C0029792|ICD9CM|PT|304.60|Other specified drug dependence, unspecified
C0029792|ICD9CM|HT|304.6|Other specified drug dependence
C0029792|ICD9CM|AB|304.60|Drug depend NEC-unspec
C0029793|ICD9CM|PT|259.8|Other specified endocrine disorders
C0029793|ICD9CM|AB|259.8|Endocrine disorders NEC
C0029794|ICD9CM|HT|695.8|Other specified erythematous conditions
C0029794|ICD9CM|PT|695.89|Other specified erythematous conditions
C0029794|ICD9CM|AB|695.89|Erythematous cond NEC
C0029795|ICD9CM|PT|V61.9|Unspecified family circumstance
C0029795|ICD9CM|AB|V61.9|Family circumstance NOS
C0029796|ICD9CM|PT|125.6|Other specified filariasis
C0029796|ICD9CM|AB|125.6|Filariasis NEC
C0029797|ICD9CM|PT|619.8|Other specified fistulas involving female genital tract
C0029797|ICD9CM|AB|619.8|Fem genital fistula NEC
C0029799|ICD9CM|HT|511.8|Other specified forms of pleural effusion, except tuberculous
C0029800|ICD9CM|HT|535.4|Other specified gastritis
C0029801|ICD9CM|HT|618.8|Other specified genital prolapse
C0029801|ICD9CM|PT|618.89|Other specified genital prolapse
C0029801|ICD9CM|AB|618.89|Genital prolapse NEC
C0029802|ICD9CM|HT|365.8|Other specified forms of glaucoma
C0029802|ICD9CM|AB|365.89|Glaucoma NEC
C0029802|ICD9CM|PT|365.89|Other specified glaucoma
C0029803|ICD9CM|PT|128.8|Other specified helminthiasis
C0029803|ICD9CM|AB|128.8|Helminthiasis NEC
C0029804|ICD9CM|PT|287.8|Other specified hemorrhagic conditions
C0029804|ICD9CM|AB|287.8|Hemorrhagic cond NEC
C0029805|ICD9CM|PT|701.8|Other specified hypertrophic and atrophic conditions of skin
C0029805|ICD9CM|AB|701.8|Skin hypertro/atroph NEC
C0029806|ICD9CM|PT|343.8|Other specified infantile cerebral palsy
C0029806|ICD9CM|AB|343.8|Cerebral palsy NEC
C0029807|ICD9CM|PT|614.8|Other specified inflammatory disease of female pelvic organs and tissues
C0029807|ICD9CM|AB|614.8|Fem pelv inflam dis NEC
C0029808|ICD9CM|PT|127.7|Other specified intestinal helminthiasis
C0029808|ICD9CM|AB|127.7|Intest helminthiasis NEC
C0029809|ICD9CM|PT|579.8|Other specified intestinal malabsorption
C0029809|ICD9CM|AB|579.8|Intest malabsorption NEC
C0029810|ICD9CM|PT|280.8|Other specified iron deficiency anemias
C0029810|ICD9CM|AB|280.8|Iron defic anemia NEC
C0029811|ICD9CM|PT|030.8|Other specified leprosy
C0029811|ICD9CM|AB|030.8|Leprosy NEC
C0029812|ICD9CM|HT|207|Other specified leukemia
C0029812|ICD9CM|HT|207.8|Other specified leukemia
C0029813|ICD9CM|PT|686.8|Other specified local infections of skin and subcutaneous tissue
C0029813|ICD9CM|AB|686.8|Local skin infection NEC
C0029815|ICD9CM|HT|036.8|Other specified meningococcal infections
C0029815|ICD9CM|PT|036.89|Other specified meningococcal infections
C0029815|ICD9CM|AB|036.89|Meningococcal infect NEC
C0029816|ICD9CM|PT|358.8|Other specified myoneural disorders
C0029816|ICD9CM|AB|358.8|Myoneural disorders NEC
C0029817|ICD9CM|HT|094.8|Other specified neurosyphilis
C0029817|ICD9CM|PT|094.89|Other specified neurosyphilis
C0029817|ICD9CM|AB|094.89|Neurosyphilis NEC
C0029818|ICD9CM|PT|049.8|Other specified non-arthropod-borne viral diseases of central nervous system
C0029818|ICD9CM|AB|049.8|Viral encephalitis NEC
C0029819|ICD9CM|PT|623.8|Other specified noninflammatory disorders of vagina
C0029819|ICD9CM|AB|623.8|Noninflam dis vagina NEC
C0029821|ICD9CM|PT|523.8|Other specified periodontal diseases
C0029821|ICD9CM|AB|523.8|Periodontal disease NEC
C0029822|ICD9CM|HT|443.8|Other specified peripheral vascular diseases
C0029823|ICD9CM|HT|567.8|Other specified peritonitis
C0029823|ICD9CM|PT|567.89|Other specified peritonitis
C0029823|ICD9CM|AB|567.89|Peritonitis NEC
C0029824|ICD9CM|PT|306.8|Other specified psychophysiological malfunction
C0029824|ICD9CM|AB|306.8|Psychogenic disorder NEC
C0029825|ICD9CM|HT|302.8|Other specified psychosexual disorders
C0029825|ICD9CM|PT|302.89|Other specified psychosexual disorders
C0029825|ICD9CM|AB|302.89|Psychosexual dis NEC
C0029826|ICD9CM|PT|003.8|Other specified salmonella infections
C0029826|ICD9CM|AB|003.8|Salmonella infection NEC
C0029827|ICD9CM|PT|120.8|Other specified schistosomiasis
C0029827|ICD9CM|AB|120.8|Schistosomiasis NEC
C0029829|ICD9CM|PT|848.8|Other specified sites of sprains and strains
C0029829|ICD9CM|AB|848.8|Sprain NEC
C0029830|ICD9CM|PT|104.8|Other specified spirochetal infections
C0029830|ICD9CM|AB|104.8|Spirochetal infect NEC
C0029831|ICD9CM|HT|378.7|Other specified strabismus
C0029832|ICD9CM|PT|063.8|Other specified tick-borne viral encephalitis
C0029832|ICD9CM|AB|063.8|Tick-borne enceph NEC
C0029833|ICD9CM|PT|121.8|Other specified trematode infections
C0029833|ICD9CM|AB|121.8|Trematode infection NEC
C0029834|ICD9CM|PT|350.8|Other specified trigeminal nerve disorders
C0029834|ICD9CM|AB|350.8|Trigeminal nerve dis NEC
C0029835|ICD9CM|PT|021.8|Other specified tularemia
C0029835|ICD9CM|AB|021.8|Tularemia NEC
C0029836|ICD9CM|HT|595.8|Other specified types of cystitis
C0029836|ICD9CM|PT|595.89|Other specified types of cystitis
C0029836|ICD9CM|AB|595.89|Cystitis NEC
C0029837|ICD9CM|PT|603.8|Other specified types of hydrocele
C0029837|ICD9CM|AB|603.8|Hydrocele NEC
C0029838|ICD9CM|PT|295.80|Other specified types of schizophrenia, unspecified
C0029838|ICD9CM|HT|295.8|Other specified types of schizophrenia
C0029838|ICD9CM|AB|295.80|Schizophrenia NEC-unspec
C0029839|ICD9CM|PT|708.8|Other specified urticaria
C0029839|ICD9CM|AB|708.8|Urticaria NEC
C0029840|ICD9CM|PT|099.8|Other specified venereal diseases
C0029840|ICD9CM|AB|099.8|Venereal disease NEC
C0029841|ICD9CM|PT|057.8|Other specified viral exanthemata
C0029841|ICD9CM|AB|057.8|Viral exanthemata NEC
C0029842|ICD9CM|PT|079.89|Other specified viral infection
C0029842|ICD9CM|AB|079.89|Oth specf viral infectn
C0029843|ICD9CM|PT|047.8|Other specified viral meningitis
C0029843|ICD9CM|AB|047.8|Viral meningitis NEC
C0029844|ICD9CM|PT|368.8|Other specified visual disturbances
C0029844|ICD9CM|AB|368.8|Visual disturbances NEC
C0029846|ICD9CM|PT|93.75|Other speech training and therapy
C0029846|ICD9CM|AB|93.75|Other speech therapy
C0029848|ICD9CM|PT|335.19|Other spinal muscular atrophy
C0029848|ICD9CM|AB|335.19|Spinal muscl atrophy NEC
C0029849|ICD9CM|PT|334.8|Other spinocerebellar diseases
C0029849|ICD9CM|AB|334.8|Spinocerebellar dis NEC
C0029851|ICD9CM|PT|33.39|Other surgical collapse of lung
C0029851|ICD9CM|AB|33.39|Surg collaps of lung NEC
C0029853|ICD9CM|PT|05.29|Other sympathectomy and ganglionectomy
C0029853|ICD9CM|AB|05.29|Other sympathectomy
C0029854|ICD9CM|PT|785.9|Other symptoms involving cardiovascular system
C0029854|ICD9CM|AB|785.9|Cardiovas sys symp NEC
C0029855|ICD9CM|HT|784.9|Other symptoms involving head and neck
C0029855|ICD9CM|PT|784.99|Other symptoms involving head and neck
C0029855|ICD9CM|AB|784.99|Head & neck symptoms NEC
C0029856|ICD9CM|PT|727.09|Other synovitis and tenosynovitis
C0029856|ICD9CM|AB|727.09|Synovitis NEC
C0029857|ICD9CM|PT|257.8|Other testicular dysfunction
C0029857|ICD9CM|AB|257.8|Testicular dysfunct NEC
C0029858|ICD9CM|PT|257.2|Other testicular hypofunction
C0029858|ICD9CM|AB|257.2|Testicular hypofunc NEC
C0029860|ICD9CM|AB|96.39|Other transanal enema
C0029860|ICD9CM|PT|96.39|Other transanal enema
C0029861|ICD9CM|PT|99.03|Other transfusion of whole blood
C0029861|ICD9CM|AB|99.03|Whole blood transfus NEC
C0029862|ICD9CM|PT|50.59|Other transplant of liver
C0029862|ICD9CM|AB|50.59|Liver transplant NEC
C0029863|ICD9CM|PT|85.34|Other unilateral subcutaneous mammectomy
C0029863|ICD9CM|AB|85.34|Unilat subq mammect NEC
C0029865|ICD9CM|PT|V61.7|Other unwanted pregnancy
C0029865|ICD9CM|AB|V61.7|Unwanted pregnancy NEC
C0029866|ICD9CM|PT|593.4|Other ureteric obstruction
C0029866|ICD9CM|AB|593.4|Ureteric obstruction NEC
C0029867|ICD9CM|HT|597.8|Other urethritis
C0029867|ICD9CM|PT|597.89|Other urethritis
C0029867|ICD9CM|AB|597.89|Urethritis NEC
C0029869|ICD9CM|PT|72.79|Other vacuum extraction
C0029869|ICD9CM|AB|72.79|Vacuum extract del NEC
C0029870|ICD9CM|PT|553.29|Other ventral hernia without mention of obstruction or gangrene
C0029870|ICD9CM|AB|553.29|Ventral hernia NEC
C0029871|ICD9CM|PT|077.8|Other viral conjunctivitis
C0029871|ICD9CM|AB|077.8|Viral conjunctivitis NEC
C0029872|ICD9CM|PT|379.24|Other vitreous opacities
C0029872|ICD9CM|AB|379.24|Vitreous opacities NEC
C0029874|ICD9CM|HT|88.1|Other x-ray of abdomen
C0029874|ICD9CM|PT|88.19|Other x-ray of abdomen
C0029874|ICD9CM|AB|88.19|Abdominal x-ray NEC
C0029875|ICD9CM|PT|87.17|Other x-ray of skull
C0029875|ICD9CM|AB|87.17|Skull x-ray NEC
C0029876|ICD9CM|HT|839|Other, multiple, and ill-defined dislocations
C0029882|ICD9CM|AB|382.9|Otitis media NOS
C0029882|ICD9CM|PT|382.9|Unspecified otitis media
C0029888|ICD9CM|AB|382.4|Suppur otitis media NOS
C0029888|ICD9CM|PT|382.4|Unspecified suppurative otitis media
C0029888|ICD9CM|HT|382|Suppurative and unspecified otitis media
C0029899|ICD9CM|HT|387|Otosclerosis
C0029899|ICD9CM|AB|387.9|Otosclerosis NOS
C0029899|ICD9CM|PT|387.9|Otosclerosis, unspecified
C0030193|ICD9CM|HT|338-338.99|PAIN
C0030196|ICD9CM|AB|729.5|Pain in limb
C0030196|ICD9CM|PT|729.5|Pain in limb
C0030197|ICD9CM|AB|379.91|Pain in or around eye
C0030197|ICD9CM|PT|379.91|Pain in or around eye
C0030232|ICD9CM|AB|782.61|Pallor
C0030232|ICD9CM|PT|782.61|Pallor
C0030252|ICD9CM|AB|785.1|Palpitations
C0030252|ICD9CM|PT|785.1|Palpitations
C0030275|ICD9CM|HT|52.8|Transplant of pancreas
C0030275|ICD9CM|PT|52.80|Pancreatic transplant, not otherwise specified
C0030275|ICD9CM|AB|52.80|Pancreat transplant NOS
C0030286|ICD9CM|AB|577.9|Pancreatic disease NOS
C0030286|ICD9CM|HT|577|Diseases of pancreas
C0030286|ICD9CM|PT|577.9|Unspecified disease of pancreas
C0030312|ICD9CM|HT|284.1|Pancytopenia
C0030326|ICD9CM|PT|729.30|Panniculitis, unspecified site
C0030326|ICD9CM|HT|729.3|Panniculitis, unspecified
C0030326|ICD9CM|AB|729.30|Panniculitis, unsp site
C0030332|ICD9CM|AB|360.02|Panophthalmitis
C0030332|ICD9CM|PT|360.02|Panophthalmitis
C0030343|ICD9CM|AB|360.12|Panuveitis
C0030343|ICD9CM|PT|360.12|Panuveitis
C0030353|ICD9CM|HT|377.0|Papilledema
C0030353|ICD9CM|AB|377.00|Papilledema NOS
C0030353|ICD9CM|AB|377.31|Optic papillitis
C0030353|ICD9CM|PT|377.31|Optic papillitis
C0030353|ICD9CM|PT|377.00|Papilledema, unspecified
C0030372|ICD9CM|AB|066.0|Phlebotomus fever
C0030372|ICD9CM|PT|066.0|Phlebotomus fever
C0030409|ICD9CM|AB|116.1|Paracoccidioidomycosis
C0030409|ICD9CM|PT|116.1|Paracoccidioidomycosis
C0030424|ICD9CM|AB|121.2|Paragonimiasis
C0030424|ICD9CM|PT|121.2|Paragonimiasis
C0030442|ICD9CM|AB|335.22|Progressive bulbar palsy
C0030442|ICD9CM|PT|335.22|Progressive bulbar palsy
C0030446|ICD9CM|AB|560.1|Paralytic ileus
C0030446|ICD9CM|PT|560.1|Paralytic ileus
C0030477|ICD9CM|PT|301.0|Paranoid personality disorder
C0030477|ICD9CM|AB|301.0|Paranoid personality
C0030484|ICD9CM|AB|297.2|Paraphrenia
C0030484|ICD9CM|PT|297.2|Paraphrenia
C0030486|ICD9CM|PT|344.1|Paraplegia
C0030486|ICD9CM|AB|344.1|Paraplegia NOS
C0030491|ICD9CM|AB|696.2|Parapsoriasis
C0030491|ICD9CM|PT|696.2|Parapsoriasis
C0030517|ICD9CM|PT|252.9|Unspecified disorder of parathyroid gland
C0030517|ICD9CM|AB|252.9|Parathyroid disorder NOS
C0030517|ICD9CM|HT|252|Disorders of parathyroid gland
C0030528|ICD9CM|AB|002.9|Paratyphoid fever NOS
C0030528|ICD9CM|PT|002.9|Paratyphoid fever, unspecified
C0030548|ICD9CM|PT|99.15|Parenteral infusion of concentrated nutritional substances
C0030548|ICD9CM|AB|99.15|Parent infus nutrit sub
C0030567|ICD9CM|HT|332|Parkinson's disease
C0030567|ICD9CM|AB|332.0|Paralysis agitans
C0030567|ICD9CM|PT|332.0|Paralysis agitans
C0030569|ICD9CM|AB|332.1|Secondary parkinsonism
C0030569|ICD9CM|PT|332.1|Secondary parkinsonism
C0030590|ICD9CM|PT|427.0|Paroxysmal supraventricular tachycardia
C0030590|ICD9CM|AB|427.0|Parox atrial tachycardia
C0030591|ICD9CM|PT|427.1|Paroxysmal ventricular tachycardia
C0030591|ICD9CM|AB|427.1|Parox ventric tachycard
C0030593|ICD9CM|AB|363.21|Pars planitis
C0030593|ICD9CM|PT|363.21|Pars planitis
C0030631|ICD9CM|PT|301.84|Passive-aggressive personality
C0030631|ICD9CM|AB|301.84|Passive-aggressiv person
C0030636|ICD9CM|AB|027.2|Pasteurellosis
C0030636|ICD9CM|PT|027.2|Pasteurellosis
C0030662|ICD9CM|AB|312.31|Pathological gambling
C0030662|ICD9CM|PT|312.31|Pathological gambling
C0030756|ICD9CM|AB|132.9|Pediculosis NOS
C0030756|ICD9CM|PT|132.9|Pediculosis, unspecified
C0030757|ICD9CM|PT|132.0|Pediculus capitis [head louse]
C0030757|ICD9CM|AB|132.0|Pediculus capitis
C0030758|ICD9CM|PT|132.1|Pediculus corporis [body louse]
C0030758|ICD9CM|AB|132.1|Pediculus corporis
C0030759|ICD9CM|AB|132.2|Phthirus pubis
C0030759|ICD9CM|PT|132.2|Phthirus pubis [pubic louse]
C0030764|ICD9CM|AB|302.2|Pedophilia
C0030764|ICD9CM|PT|302.2|Pedophilia
C0030783|ICD9CM|AB|265.2|Pellagra
C0030783|ICD9CM|PT|265.2|Pellagra
C0030788|ICD9CM|AB|68.8|Pelvic evisceration
C0030788|ICD9CM|PT|68.8|Pelvic evisceration
C0030796|ICD9CM|AB|88.25|Pelvimetry
C0030796|ICD9CM|PT|88.25|Pelvimetry
C0030804|ICD9CM|HT|694.6|Benign mucous membrane pemphigoid
C0030805|ICD9CM|AB|694.5|Pemphigoid
C0030805|ICD9CM|PT|694.5|Pemphigoid
C0030807|ICD9CM|AB|694.4|Pemphigus
C0030807|ICD9CM|PT|694.4|Pemphigus
C0030846|ICD9CM|HT|607|Disorders of penis
C0030846|ICD9CM|AB|607.9|Disorder of penis NOS
C0030846|ICD9CM|PT|607.9|Unspecified disorder of penis
C0030848|ICD9CM|AB|607.85|Peyronie's disease
C0030848|ICD9CM|PT|607.85|Peyronie's disease
C0030920|ICD9CM|HT|533|Peptic ulcer, site unspecified
C0030923|ICD9CM|HT|533.9|Peptic ulcer of unspecified site, unspecified as acute or chronic, without mention of hemorrhage or perforation
C0030924|ICD9CM|PT|533.90|Peptic ulcer of unspecified site, unspecified as acute or chronic, without mention of hemorrhage or perforation, without mention of obstruction
C0030924|ICD9CM|AB|533.90|Peptic ulcer NOS
C0030990|ICD9CM|PT|55.03|Percutaneous nephrostomy without fragmentation
C0030990|ICD9CM|AB|55.03|Percu nephrostm w/o frag
C0031036|ICD9CM|AB|446.0|Polyarteritis nodosa
C0031036|ICD9CM|PT|446.0|Polyarteritis nodosa
C0031042|ICD9CM|AB|37.31|Pericardiectomy
C0031042|ICD9CM|PT|37.31|Pericardiectomy
C0031048|ICD9CM|PT|423.2|Constrictive pericarditis
C0031048|ICD9CM|AB|423.2|Constrictiv pericarditis
C0031069|ICD9CM|PT|277.31|Familial Mediterranean fever
C0031069|ICD9CM|AB|277.31|Fam Mediterranean fever
C0031115|ICD9CM|PT|443.81|Peripheral angiopathy in diseases classified elsewhere
C0031115|ICD9CM|AB|443.81|Angiopathy in other dis
C0031139|ICD9CM|AB|54.98|Peritoneal dialysis
C0031139|ICD9CM|PT|54.98|Peritoneal dialysis
C0031142|ICD9CM|PT|568.9|Unspecified disorder of peritoneum
C0031142|ICD9CM|AB|568.9|Peritoneal disorder NOS
C0031144|ICD9CM|AB|568.82|Peritoneal effusion
C0031144|ICD9CM|PT|568.82|Peritoneal effusion (chronic)
C0031148|ICD9CM|AB|54.25|Peritoneal lavage
C0031148|ICD9CM|PT|54.25|Peritoneal lavage
C0031150|ICD9CM|AB|54.21|Laparoscopy
C0031150|ICD9CM|PT|54.21|Laparoscopy
C0031152|ICD9CM|PT|54.94|Creation of peritoneovascular shunt
C0031152|ICD9CM|AB|54.94|Creat peritoneovas shunt
C0031154|ICD9CM|AB|567.9|Peritonitis NOS
C0031154|ICD9CM|PT|567.9|Unspecified peritonitis
C0031157|ICD9CM|AB|475|Peritonsillar abscess
C0031157|ICD9CM|PT|475|Peritonsillar abscess
C0031190|ICD9CM|PT|747.83|Persistent fetal circulation
C0031190|ICD9CM|AB|747.83|Persistent fetal circ
C0031192|ICD9CM|AB|745.61|Ostium primum defect
C0031192|ICD9CM|PT|745.61|Ostium primum defect
C0031212|ICD9CM|HT|301|Personality disorders
C0031212|ICD9CM|AB|301.9|Personality disorder NOS
C0031212|ICD9CM|PT|301.9|Unspecified personality disorder
C0031315|ICD9CM|AB|353.6|Phantom limb (syndrome)
C0031315|ICD9CM|PT|353.6|Phantom limb (syndrome)
C0031345|ICD9CM|AB|478.20|Disease of pharynx NOS
C0031345|ICD9CM|PT|478.20|Unspecified disease of pharynx
C0031349|ICD9CM|HT|29.3|Excision or destruction of lesion or tissue of pharynx
C0031351|ICD9CM|PT|077.2|Pharyngoconjunctival fever
C0031351|ICD9CM|AB|077.2|Pharyngoconjunct fever
C0031485|ICD9CM|AB|270.1|Phenylketonuria - pku
C0031485|ICD9CM|PT|270.1|Phenylketonuria [PKU]
C0031545|ICD9CM|HT|88.6|Phlebography
C0031548|ICD9CM|AB|39.32|Suture of vein
C0031548|ICD9CM|PT|39.32|Suture of vein
C0031572|ICD9CM|AB|300.23|Social phobia
C0031572|ICD9CM|PT|300.23|Social phobia
C0031707|ICD9CM|PT|275.3|Disorders of phosphorus metabolism
C0031707|ICD9CM|AB|275.3|Dis phosphorus metabol
C0031809|ICD9CM|PT|89.7|General physical examination
C0031809|ICD9CM|AB|89.7|General physical exam
C0031873|ICD9CM|AB|307.52|Pica
C0031873|ICD9CM|PT|307.52|Pica
C0031880|ICD9CM|PT|278.03|Obesity hypoventilation syndrome
C0031880|ICD9CM|AB|278.03|Obesity hypovent synd
C0031925|ICD9CM|HT|685|Pilonidal cyst
C0031946|ICD9CM|HT|103|Pinta
C0031946|ICD9CM|AB|103.9|Pinta NOS
C0031946|ICD9CM|PT|103.9|Pinta, unspecified
C0032026|ICD9CM|AB|696.3|Pityriasis rosea
C0032026|ICD9CM|PT|696.3|Pityriasis rosea
C0032027|ICD9CM|AB|696.4|Pityriasis rubra pilaris
C0032027|ICD9CM|PT|696.4|Pityriasis rubra pilaris
C0032064|ICD9CM|HT|020|Plague
C0032064|ICD9CM|AB|020.9|Plague NOS
C0032064|ICD9CM|PT|020.9|Plague, unspecified
C0032134|ICD9CM|PT|99.71|Therapeutic plasmapheresis
C0032134|ICD9CM|AB|99.71|Therapeu plasmapheresis
C0032202|ICD9CM|PT|99.74|Therapeutic plateletpheresis
C0032202|ICD9CM|AB|99.74|Therapeu plateltpheresis
C0032216|ICD9CM|AB|94.36|Play psychotherapy
C0032216|ICD9CM|PT|94.36|Play psychotherapy
C0032221|ICD9CM|AB|89.58|Plethysmogram
C0032221|ICD9CM|PT|89.58|Plethysmogram
C0032227|ICD9CM|AB|511.9|Pleural effusion NOS
C0032227|ICD9CM|PT|511.9|Unspecified pleural effusion
C0032231|ICD9CM|HT|511|Pleurisy
C0032232|ICD9CM|PT|511.0|Pleurisy without mention of effusion or current tuberculosis
C0032232|ICD9CM|AB|511.0|Pleurisy w/o effus or TB
C0032238|ICD9CM|AB|074.1|Epidemic pleurodynia
C0032238|ICD9CM|PT|074.1|Epidemic pleurodynia
C0032272|ICD9CM|PT|041.2|Pneumococcus infection in conditions classified elsewhere and of unspecified site
C0032272|ICD9CM|AB|041.2|Pneumococcus infect NOS
C0032273|ICD9CM|AB|505|Pneumoconiosis NOS
C0032273|ICD9CM|PT|505|Pneumoconiosis, unspecified
C0032274|ICD9CM|PT|503|Pneumoconiosis due to other inorganic dust
C0032274|ICD9CM|AB|503|Inorg dust pneumocon NEC
C0032279|ICD9CM|AB|87.01|Pneumoencephalogram
C0032279|ICD9CM|PT|87.01|Pneumoencephalogram
C0032284|ICD9CM|HT|32.5|Pneumonectomy
C0032286|ICD9CM|HT|482.8|Pneumonia due to other specified bacteria
C0032286|ICD9CM|PT|482.89|Pneumonia due to other specified bacteria
C0032286|ICD9CM|AB|482.89|Pneumonia oth spcf bact
C0032287|ICD9CM|HT|483|Pneumonia due to other specified organism
C0032287|ICD9CM|PT|483.8|Pneumonia due to other specified organism
C0032287|ICD9CM|AB|483.8|Pneumon oth spec orgnsm
C0032302|ICD9CM|PT|483.0|Pneumonia due to mycoplasma pneumoniae
C0032302|ICD9CM|AB|483.0|Pneu mycplsm pneumoniae
C0032308|ICD9CM|HT|482.4|Pneumonia due to Staphylococcus
C0032308|ICD9CM|PT|482.40|Pneumonia due to Staphylococcus, unspecified
C0032308|ICD9CM|AB|482.40|Staphylococcal pneu NOS
C0032310|ICD9CM|HT|480|Viral pneumonia
C0032310|ICD9CM|AB|480.9|Viral pneumonia NOS
C0032310|ICD9CM|PT|480.9|Viral pneumonia, unspecified
C0032318|ICD9CM|PT|504|Pneumonopathy due to inhalation of other dust
C0032318|ICD9CM|AB|504|Dust pneumonopathy NEC
C0032328|ICD9CM|PT|33.32|Artificial pneumothorax for collapse of lung
C0032328|ICD9CM|AB|33.32|Pnemothorax-lung collaps
C0032371|ICD9CM|HT|045|Acute poliomyelitis
C0032371|ICD9CM|HT|045.9|Acute poliomyelitis, unspecified
C0032372|ICD9CM|HT|045.0|Acute paralytic poliomyelitis specified as bulbar
C0032460|ICD9CM|AB|256.4|Polycystic ovaries
C0032460|ICD9CM|PT|256.4|Polycystic ovaries
C0032463|ICD9CM|AB|238.4|Polycythemia vera
C0032463|ICD9CM|PT|238.4|Polycythemia vera
C0032533|ICD9CM|AB|725|Polymyalgia rheumatica
C0032533|ICD9CM|PT|725|Polymyalgia rheumatica
C0032617|ICD9CM|AB|788.42|Polyuria
C0032617|ICD9CM|PT|788.42|Polyuria
C0032633|ICD9CM|AB|705.81|Dyshidrosis
C0032633|ICD9CM|PT|705.81|Dyshidrosis
C0032650|ICD9CM|AB|727.51|Popliteal synovial cyst
C0032650|ICD9CM|PT|727.51|Synovial cyst of popliteal space
C0032708|ICD9CM|PT|277.1|Disorders of porphyrin metabolism
C0032708|ICD9CM|AB|277.1|Dis porphyrin metabolism
C0032763|ICD9CM|PT|564.2|Postgastric surgery syndromes
C0032763|ICD9CM|AB|564.2|Postgastric surgery synd
C0032776|ICD9CM|AB|627.1|Postmenopausal bleeding
C0032776|ICD9CM|PT|627.1|Postmenopausal bleeding
C0032781|ICD9CM|PT|784.91|Postnasal drip
C0032781|ICD9CM|AB|784.91|Postnasal drip
C0032792|ICD9CM|HT|998.0|Postoperative shock
C0032792|ICD9CM|AB|998.00|Postoperative shock, NOS
C0032792|ICD9CM|PT|998.00|Postoperative shock, unspecified
C0032797|ICD9CM|HT|666|Postpartum hemorrhage
C0032807|ICD9CM|HT|459.1|Postphlebitic syndrome
C0032811|ICD9CM|AB|V45.81|Aortocoronary bypass
C0032811|ICD9CM|PT|V45.81|Aortocoronary bypass status
C0032816|ICD9CM|HT|339.2|Post-traumatic headache
C0032816|ICD9CM|PT|339.20|Post-traumatic headache, unspecified
C0032816|ICD9CM|AB|339.20|Post-trauma headache NOS
C0032870|ICD9CM|AB|059.9|Poxvirus infection NOS
C0032870|ICD9CM|PT|059.9|Poxvirus infections, unspecified
C0032897|ICD9CM|PT|759.81|Prader-Willi syndrome
C0032897|ICD9CM|AB|759.81|Prader-willi syndrome
C0032962|ICD9CM|HT|646.9|Unspecified complication of pregnancy
C0032969|ICD9CM|PT|648.03|Diabetes mellitus of mother, complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C0032969|ICD9CM|AB|648.03|Diabetes-antepartum
C0032984|ICD9CM|HT|633.0|Abdominal pregnancy
C0032987|ICD9CM|HT|633|Ectopic pregnancy
C0032987|ICD9CM|HT|633.9|Unspecified ectopic pregnancy
C0032989|ICD9CM|HT|651.9|Unspecified multiple gestation
C0032989|ICD9CM|HT|651|Multiple gestation
C0032989|ICD9CM|PT|651.90|Unspecified multiple gestation, unspecified as to episode of care or not applicable
C0032989|ICD9CM|AB|651.90|Multi gestat NOS-unspec
C0032991|ICD9CM|HT|633.2|Ovarian pregnancy
C0032993|ICD9CM|HT|645.2|Prolonged pregnancy
C0032993|ICD9CM|HT|645.1|Post term pregnancy
C0032994|ICD9CM|HT|633.1|Tubal pregnancy
C0033036|ICD9CM|AB|427.61|Atrial premature beats
C0033036|ICD9CM|PT|427.61|Supraventricular premature beats
C0033038|ICD9CM|AB|302.75|Premature ejaculation
C0033038|ICD9CM|PT|302.75|Premature ejaculation
C0033074|ICD9CM|AB|388.01|Presbyacusis
C0033074|ICD9CM|PT|388.01|Presbyacusis
C0033075|ICD9CM|AB|367.4|Presbyopia
C0033075|ICD9CM|PT|367.4|Presbyopia
C0033117|ICD9CM|AB|607.3|Priapism
C0033117|ICD9CM|PT|607.3|Priapism
C0033132|ICD9CM|PT|334.2|Primary cerebellar degeneration
C0033132|ICD9CM|AB|334.2|Primary cerebellar degen
C0033359|ICD9CM|PT|056.01|Encephalomyelitis due to rubella
C0033359|ICD9CM|AB|056.01|Rubella encephalitis
C0033467|MTH|PN|NOCODE|Vaccination NEC in ICD9CM
C0033467|ICD9CM|PT|99.55|Prophylactic administration of vaccine against other diseases
C0033467|ICD9CM|AB|99.55|Vaccination NEC
C0033575|ICD9CM|AB|602.9|Prostatic disorder NOS
C0033575|ICD9CM|PT|602.9|Unspecified disorder of prostate
C0033581|ICD9CM|AB|601.9|Prostatitis NOS
C0033581|ICD9CM|HT|601|Inflammatory diseases of prostate
C0033581|ICD9CM|PT|601.9|Prostatitis, unspecified
C0033677|ICD9CM|PT|263.9|Unspecified protein-calorie malnutrition
C0033677|ICD9CM|AB|263.9|Protein-cal malnutr NOS
C0033687|ICD9CM|AB|791.0|Proteinuria
C0033687|ICD9CM|PT|791.0|Proteinuria
C0033698|ICD9CM|PT|041.6|Proteus (mirabilis) (morganii) infection in conditions classified elsewhere and of unspecified site
C0033698|ICD9CM|AB|041.6|Proteus infection NOS
C0033770|ICD9CM|AB|756.71|Prune belly syndrome
C0033770|ICD9CM|PT|756.71|Prune belly syndrome
C0033771|ICD9CM|AB|698.2|Prurigo
C0033771|ICD9CM|PT|698.2|Prurigo
C0033774|ICD9CM|PT|698.9|Unspecified pruritic disorder
C0033774|ICD9CM|AB|698.9|Pruritic disorder NOS
C0033775|ICD9CM|AB|698.0|Pruritus ani
C0033775|ICD9CM|PT|698.0|Pruritus ani
C0033777|ICD9CM|PT|698.1|Pruritus of genital organs
C0033777|ICD9CM|AB|698.1|Pruritus of genitalia
C0033790|ICD9CM|AB|335.23|Pseudobulbar palsy
C0033790|ICD9CM|PT|335.23|Pseudobulbar palsy
C0033816|ICD9CM|PT|041.7|Pseudomonas infection in conditions classified elsewhere and of unspecified site
C0033816|ICD9CM|AB|041.7|Pseudomonas infect NOS
C0033825|ICD9CM|PT|V43.1|Lens replaced by other means
C0033825|ICD9CM|AB|V43.1|Lens replacement NEC
C0033845|ICD9CM|AB|348.2|Pseudotumor cerebri
C0033845|ICD9CM|PT|348.2|Benign intracranial hypertension
C0033889|ICD9CM|AB|94.43|Psychodrama
C0033889|ICD9CM|PT|94.43|Psychodrama
C0033893|ICD9CM|AB|307.81|Tension headache
C0033893|ICD9CM|PT|307.81|Tension headache
C0033893|ICD9CM|AB|339.10|Tension headache NOS
C0033893|ICD9CM|HT|339.1|Tension type headache
C0033893|ICD9CM|PT|339.10|Tension type headache, unspecified
C0033905|ICD9CM|PT|94.02|Administration of psychologic test
C0033905|ICD9CM|AB|94.02|Psychologic test adminis
C0033936|ICD9CM|PT|291.9|Unspecified alcohol-induced mental disorders
C0033936|ICD9CM|AB|291.9|Alcohol mental disor NOS
C0033937|ICD9CM|HT|292.1|Drug-induced psychotic disorders
C0033948|ICD9CM|AB|302.73|Female orgasmic disorder
C0033948|ICD9CM|PT|302.73|Female orgasmic disorder
C0033950|ICD9CM|PT|302.72|Psychosexual dysfunction with inhibited sexual excitement
C0033950|ICD9CM|AB|302.72|Inhibited sex excitement
C0033951|ICD9CM|PT|302.79|Psychosexual dysfunction with other specified psychosexual dysfunctions
C0033951|ICD9CM|AB|302.79|Psychosexual dysfunc NEC
C0033953|ICD9CM|PT|302.9|Unspecified psychosexual disorder
C0033953|ICD9CM|AB|302.9|Psychosexual dis NOS
C0033975|ICD9CM|HT|290-299.99|PSYCHOSES
C0033975|ICD9CM|AB|298.9|Psychosis NOS
C0033975|ICD9CM|PT|298.9|Unspecified psychosis
C0034050|ICD9CM|PT|516.0|Pulmonary alveolar proteinosis
C0034050|ICD9CM|AB|516.0|Pul alveolar proteinosis
C0034066|ICD9CM|HT|415.1|Pulmonary embolism and infarction
C0034067|ICD9CM|HT|492|Emphysema
C0034068|ICD9CM|AB|518.3|Pulmonary eosinophilia
C0034068|ICD9CM|PT|518.3|Pulmonary eosinophilia
C0034076|ICD9CM|HT|518.5|Pulmonary insufficiency following trauma and surgery
C0034084|ICD9CM|PT|746.83|Infundibular pulmonic stenosis
C0034084|ICD9CM|AB|746.83|Infundib pulmon stenosis
C0034087|ICD9CM|AB|424.3|Pulmonary valve disorder
C0034087|ICD9CM|PT|424.3|Pulmonary valve disorders
C0034100|ICD9CM|PT|522.2|Pulp degeneration
C0034100|ICD9CM|AB|522.2|Tooth pulp degeneration
C0034103|ICD9CM|AB|522.0|Pulpitis
C0034103|ICD9CM|PT|522.0|Pulpitis
C0034152|ICD9CM|AB|287.0|Allergic purpura
C0034152|ICD9CM|PT|287.0|Allergic purpura
C0034186|ICD9CM|AB|590.80|Pyelonephritis NOS
C0034186|ICD9CM|PT|590.80|Pyelonephritis, unspecified
C0034212|ICD9CM|HT|686.0|Pyoderma
C0034212|ICD9CM|AB|686.00|Pyoderma NOS
C0034212|ICD9CM|PT|686.00|Pyoderma, unspecified
C0034214|ICD9CM|PT|686.1|Pyogenic granuloma of skin and subcutaneous tissue
C0034214|ICD9CM|AB|686.1|Pyogenic granuloma
C0034362|ICD9CM|AB|083.0|Q fever
C0034362|ICD9CM|PT|083.0|Q fever
C0034372|ICD9CM|PT|344.00|Quadriplegia, unspecified
C0034372|ICD9CM|AB|344.00|Quadriplegia, unspecifd
C0034494|ICD9CM|AB|071|Rabies
C0034494|ICD9CM|PT|071|Rabies
C0034525|ICD9CM|AB|990|Effects radiation NOS
C0034525|ICD9CM|PT|990|Effects of radiation, unspecified
C0034542|ICD9CM|PT|40.40|Radical neck dissection, not otherwise specified
C0034542|ICD9CM|AB|40.40|Rad neck dissection NOS
C0034543|ICD9CM|AB|522.8|Radicular cyst
C0034543|ICD9CM|PT|522.8|Radicular cyst
C0034606|ICD9CM|HT|92|Nuclear medicine
C0034668|ICD9CM|AB|E960.1|Rape
C0034668|ICD9CM|PT|E960.1|Rape
C0034686|ICD9CM|HT|026|Rat-bite fever
C0034686|ICD9CM|AB|026.9|Rat-bite fever NOS
C0034686|ICD9CM|PT|026.9|Unspecified rat-bite fever
C0034735|ICD9CM|AB|443.0|Raynaud's syndrome
C0034735|ICD9CM|PT|443.0|Raynaud's syndrome
C0034873|ICD9CM|AB|93.81|Recreational therapy
C0034873|ICD9CM|PT|93.81|Recreation therapy
C0034880|ICD9CM|AB|388.42|Hyperacusis
C0034880|ICD9CM|PT|388.42|Hyperacusis
C0034888|ICD9CM|AB|569.1|Rectal prolapse
C0034888|ICD9CM|PT|569.1|Rectal prolapse
C0034915|ICD9CM|PT|379.93|Redness or discharge of eye
C0034915|ICD9CM|AB|379.93|Redness/discharge of eye
C0034919|ICD9CM|PT|605|Redundant prepuce and phimosis
C0034919|ICD9CM|AB|605|Redun prepuce & phimosis
C0034931|ICD9CM|HT|337.2|Reflex sympathetic dystrophy
C0034931|ICD9CM|PT|337.20|Reflex sympathetic dystrophy, unspecified
C0034931|ICD9CM|AB|337.20|Unsp rflx sympth dystrph
C0034933|ICD9CM|AB|796.1|Abnormal reflex
C0034933|ICD9CM|PT|796.1|Abnormal reflex
C0034960|ICD9CM|AB|356.3|Refsum's disease
C0034960|ICD9CM|PT|356.3|Refsum's disease
C0034996|ICD9CM|PT|93.85|Vocational rehabilitation
C0034996|ICD9CM|AB|93.85|Vocational rehabilitat
C0035012|ICD9CM|AB|099.3|Reiter's disease
C0035012|ICD9CM|PT|099.3|Reiter's disease
C0035021|ICD9CM|HT|087|Relapsing fever
C0035021|ICD9CM|AB|087.9|Relapsing fever NOS
C0035021|ICD9CM|PT|087.9|Relapsing fever, unspecified
C0035022|ICD9CM|PT|087.1|Relapsing fever, tick-borne
C0035022|ICD9CM|AB|087.1|Tick-borne relaps fever
C0035058|ICD9CM|PT|62.41|Removal of both testes at same operative episode
C0035058|ICD9CM|AB|62.41|Remove both testes
C0035060|ICD9CM|HT|36.0|Removal of coronary artery obstruction
C0035078|ICD9CM|AB|586|Renal failure NOS
C0035078|ICD9CM|PT|586|Renal failure, unspecified
C0035086|ICD9CM|AB|588.0|Renal osteodystrophy
C0035086|ICD9CM|PT|588.0|Renal osteodystrophy
C0035204|ICD9CM|PT|519.9|Unspecified disease of respiratory system
C0035204|ICD9CM|HT|460-519.99|DISEASES OF THE RESPIRATORY SYSTEM
C0035204|ICD9CM|AB|519.9|Resp system disease NOS
C0035204|ICD9CM|AB|V12.60|Hx resp system dis NOS
C0035204|ICD9CM|PT|V12.60|Personal history of unspecified disease of respiratory system
C0035220|ICD9CM|PT|769|Respiratory distress syndrome in newborn
C0035220|ICD9CM|AB|769|Respiratory distress syn
C0035238|ICD9CM|HT|748|Anomalies of respiratory system, congenital
C0035238|ICD9CM|PT|748.9|Unspecified anomaly of respiratory system
C0035238|ICD9CM|AB|748.9|Respiratory anomaly NOS
C0035239|ICD9CM|HT|93.9|Respiratory therapy
C0035258|ICD9CM|AB|333.94|Restless legs syndrome
C0035258|ICD9CM|PT|333.94|Restless legs syndrome (RLS)
C0035305|ICD9CM|AB|361.9|Retinal detachment NOS
C0035305|ICD9CM|PT|361.9|Unspecified retinal detachment
C0035309|ICD9CM|AB|362.9|Retinal disorder NOS
C0035309|ICD9CM|PT|362.9|Unspecified retinal disorder
C0035312|ICD9CM|AB|362.57|Drusen (degenerative)
C0035312|ICD9CM|PT|362.57|Drusen (degenerative)
C0035317|ICD9CM|AB|362.81|Retinal hemorrhage
C0035317|ICD9CM|PT|362.81|Retinal hemorrhage
C0035320|ICD9CM|PT|362.16|Retinal neovascularization NOS
C0035320|ICD9CM|AB|362.16|Retinal neovascular NOS
C0035326|ICD9CM|HT|362.3|Retinal vascular occlusion
C0035326|ICD9CM|PT|362.30|Retinal vascular occlusion, unspecified
C0035326|ICD9CM|AB|362.30|Retinal vasc occlus NOS
C0035344|ICD9CM|AB|362.21|Retrolental fibroplasia
C0035344|ICD9CM|PT|362.21|Retrolental fibroplasia
C0035344|ICD9CM|AB|362.20|Retinoph prematurity NOS
C0035344|ICD9CM|PT|362.20|Retinopathy of prematurity, unspecified
C0035400|ICD9CM|AB|331.81|Reye's syndrome
C0035400|ICD9CM|PT|331.81|Reye's syndrome
C0035410|ICD9CM|AB|728.88|Rhabdomyolysis
C0035410|ICD9CM|PT|728.88|Rhabdomyolysis
C0035428|ICD9CM|HT|656.1|Rhesus isoimmunization affecting management of mother
C0035436|ICD9CM|HT|390-392.99|ACUTE RHEUMATIC FEVER
C0035439|ICD9CM|PT|398.90|Rheumatic heart disease, unspecified
C0035439|ICD9CM|AB|398.90|Rheumatic heart dis NOS
C0035440|ICD9CM|PT|391.9|Acute rheumatic heart disease, unspecified
C0035440|ICD9CM|AB|391.9|Ac rheumat hrt dis NOS
C0035445|ICD9CM|PT|729.0|Rheumatism, unspecified and fibrositis
C0035445|ICD9CM|AB|729.0|Rheumatism NOS
C0035468|ICD9CM|AB|040.1|Rhinoscleroma
C0035468|ICD9CM|PT|040.1|Rhinoscleroma
C0035469|ICD9CM|AB|117.0|Rhinosporidiosis
C0035469|ICD9CM|PT|117.0|Rhinosporidiosis
C0035519|ICD9CM|AB|86.82|Facial rhytidectomy
C0035519|ICD9CM|PT|86.82|Facial rhytidectomy
C0035528|ICD9CM|AB|266.0|Ariboflavinosis
C0035528|ICD9CM|PT|266.0|Ariboflavinosis
C0035585|ICD9CM|AB|083.9|Rickettsiosis NOS
C0035585|ICD9CM|PT|083.9|Rickettsiosis, unspecified
C0035597|ICD9CM|AB|083.2|Rickettsialpox
C0035597|ICD9CM|PT|083.2|Rickettsialpox
C0035622|ICD9CM|PT|48.23|Rigid proctosigmoidoscopy
C0035622|ICD9CM|AB|48.23|Rigid proctosigmoidoscpy
C0035849|ICD9CM|AB|23.70|Root canal NOS
C0035849|ICD9CM|PT|23.70|Root canal, not otherwise specified
C0035854|ICD9CM|AB|695.3|Rosacea
C0035854|ICD9CM|PT|695.3|Rosacea
C0035920|ICD9CM|HT|056|Rubella
C0035921|ICD9CM|AB|771.0|Congenital rubella
C0035921|ICD9CM|PT|771.0|Congenital rubella
C0035945|ICD9CM|AB|E007.2|Rugby
C0035945|ICD9CM|PT|E007.2|Activities involving rugby
C0035953|ICD9CM|AB|E001.1|Running
C0035953|ICD9CM|PT|E001.1|Activities involving running
C0036091|ICD9CM|AB|527.5|Sialolithiasis
C0036091|ICD9CM|PT|527.5|Sialolithiasis
C0036093|ICD9CM|HT|527|Diseases of the salivary glands
C0036093|ICD9CM|PT|527.9|Unspecified disease of the salivary glands
C0036093|ICD9CM|AB|527.9|Salivary gland dis NOS
C0036094|ICD9CM|AB|527.4|Salivary gland fistula
C0036094|ICD9CM|PT|527.4|Fistula of salivary gland
C0036114|ICD9CM|PT|003.0|Salmonella gastroenteritis
C0036114|ICD9CM|AB|003.0|Salmonella enteritis
C0036117|ICD9CM|AB|003.9|Salmonella infection NOS
C0036117|ICD9CM|PT|003.9|Salmonella infection, unspecified
C0036133|ICD9CM|PT|614.2|Salpingitis and oophoritis not specified as acute, subacute, or chronic
C0036133|ICD9CM|AB|614.2|Salpingo-oophoritis NOS
C0036136|ICD9CM|AB|66.02|Salpingostomy
C0036136|ICD9CM|PT|66.02|Salpingostomy
C0036202|ICD9CM|AB|135|Sarcoidosis
C0036202|ICD9CM|PT|135|Sarcoidosis
C0036220|ICD9CM|HT|176|Kaposi's sarcoma
C0036220|ICD9CM|AB|176.9|Kaposi's sarcoma NOS
C0036220|ICD9CM|PT|176.9|Kaposi's sarcoma, unspecified site
C0036221|ICD9CM|HT|202.6|Malignant mast cell tumors
C0036231|ICD9CM|AB|136.5|Sarcosporidiosis
C0036231|ICD9CM|PT|136.5|Sarcosporidiosis
C0036262|ICD9CM|AB|133.0|Scabies
C0036262|ICD9CM|PT|133.0|Scabies
C0036278|ICD9CM|PT|709.2|Scar conditions and fibrosis of skin
C0036278|ICD9CM|AB|709.2|Scar & fibrosis of skin
C0036285|ICD9CM|AB|034.1|Scarlet fever
C0036285|ICD9CM|PT|034.1|Scarlet fever
C0036310|ICD9CM|PT|732.0|Juvenile osteochondrosis of spine
C0036310|ICD9CM|AB|732.0|Juv osteochondros spine
C0036323|ICD9CM|AB|120.9|Schistosomiasis NOS
C0036323|ICD9CM|HT|120|Schistosomiasis [bilharziasis]
C0036323|ICD9CM|PT|120.9|Schistosomiasis, unspecified
C0036329|ICD9CM|AB|120.2|Schistosoma japonicum
C0036329|ICD9CM|PT|120.2|Schistosomiasis due to schistosoma japonicum
C0036330|ICD9CM|AB|120.1|Schistosoma mansoni
C0036330|ICD9CM|PT|120.1|Schistosomiasis due to schistosoma mansoni
C0036337|ICD9CM|HT|295.7|Schizoaffective disorder
C0036339|ICD9CM|HT|301.2|Schizoid personality disorder
C0036339|ICD9CM|AB|301.20|Schizoid personality NOS
C0036339|ICD9CM|PT|301.20|Schizoid personality disorder, unspecified
C0036341|ICD9CM|HT|295|Schizophrenic disorders
C0036341|ICD9CM|HT|295.9|Unspecified schizophrenia
C0036341|ICD9CM|PT|295.90|Unspecified schizophrenia, unspecified
C0036341|ICD9CM|AB|295.90|Schizophrenia NOS-unspec
C0036344|ICD9CM|HT|295.2|Catatonic type schizophrenia
C0036347|ICD9CM|HT|295.1|Disorganized type schizophrenia
C0036349|ICD9CM|HT|295.3|Paranoid type schizophrenia
C0036349|ICD9CM|PT|295.30|Paranoid type schizophrenia, unspecified
C0036349|ICD9CM|AB|295.30|Paranoid schizo-unspec
C0036351|ICD9CM|PT|295.60|Schizophrenic disorders, residual type, unspecified
C0036351|ICD9CM|HT|295.6|Residual type schizophrenic disorders
C0036351|ICD9CM|AB|295.60|Schizophr dis resid NOS
C0036358|ICD9CM|HT|295.4|Schizophreniform disorder
C0036363|ICD9CM|PT|301.22|Schizotypal personality disorder
C0036363|ICD9CM|AB|301.22|Schizotypal person dis
C0036391|ICD9CM|PT|359.23|Myotonic chondrodystrophy
C0036391|ICD9CM|AB|359.23|Myotonic chondrodystrphy
C0036396|ICD9CM|AB|724.3|Sciatica
C0036396|ICD9CM|PT|724.3|Sciatica
C0036415|ICD9CM|AB|778.1|Sclerema neonatorum
C0036415|ICD9CM|PT|778.1|Sclerema neonatorum
C0036416|ICD9CM|AB|379.00|Scleritis NOS
C0036416|ICD9CM|PT|379.00|Scleritis, unspecified
C0036420|ICD9CM|PT|701.0|Circumscribed scleroderma
C0036420|ICD9CM|AB|701.0|Circumscribe scleroderma
C0036421|ICD9CM|AB|710.1|Systemic sclerosis
C0036421|ICD9CM|PT|710.1|Systemic sclerosis
C0036440|ICD9CM|PT|737.30|Scoliosis [and kyphoscoliosis], idiopathic
C0036440|ICD9CM|AB|737.30|Idiopathic scoliosis
C0036464|ICD9CM|PT|V82.89|Special screening for other specified conditions
C0036464|ICD9CM|HT|V82.8|Screening for other specified conditions
C0036464|ICD9CM|AB|V82.89|Screen for condition NEC
C0036472|ICD9CM|AB|081.2|Scrub typhus
C0036472|ICD9CM|PT|081.2|Scrub typhus
C0036502|ICD9CM|HT|706|Diseases of sebaceous glands
C0036502|ICD9CM|PT|706.9|Unspecified disease of sebaceous glands
C0036502|ICD9CM|AB|706.9|Sebaceous gland dis NOS
C0036508|ICD9CM|HT|690.1|Seborrheic dermatitis
C0036508|ICD9CM|AB|706.3|Seborrhea
C0036508|ICD9CM|PT|706.3|Seborrhea
C0036508|ICD9CM|PT|690.10|Seborrheic dermatitis, unspecified
C0036508|ICD9CM|AB|690.10|Sebrrheic dermatitis NOS
C0036528|ICD9CM|PT|197.6|Secondary malignant neoplasm of retroperitoneum and peritoneum
C0036528|ICD9CM|AB|197.6|Sec mal neo peritoneum
C0036529|ICD9CM|PT|425.9|Secondary cardiomyopathy, unspecified
C0036529|ICD9CM|AB|425.9|Second cardiomyopath NOS
C0036550|ICD9CM|HT|305.4|Sedative, hypnotic or anxiolytic abuse
C0036552|ICD9CM|HT|304.1|Sedative, hypnotic or anxiolytic dependence
C0036646|ICD9CM|HT|366.1|Senile cataract
C0036646|ICD9CM|AB|366.10|Senile cataract NOS
C0036646|ICD9CM|PT|366.10|Senile cataract, unspecified
C0036647|ICD9CM|AB|371.41|Senile corneal changes
C0036647|ICD9CM|PT|371.41|Senile corneal changes
C0036654|ICD9CM|PT|797|Senility without mention of psychosis
C0036654|ICD9CM|AB|797|Senility w/o psychosis
C0036685|ICD9CM|PT|038.40|Septicemia due to gram-negative organism, unspecified
C0036685|ICD9CM|AB|038.40|Gram-neg septicemia NOS
C0036689|ICD9CM|PT|034.0|Streptococcal sore throat
C0036689|ICD9CM|AB|034.0|Strep sore throat
C0036690|ICD9CM|HT|038|Septicemia
C0036690|ICD9CM|AB|038.9|Septicemia NOS
C0036690|ICD9CM|PT|038.9|Unspecified septicemia
C0036857|ICD9CM|PT|318.1|Severe intellectual disabilities
C0036857|ICD9CM|AB|318.1|Sev intellect disability
C0036908|ICD9CM|AB|302.83|Sexual masochism
C0036908|ICD9CM|PT|302.83|Sexual masochism
C0036913|ICD9CM|AB|302.84|Sexual sadism
C0036913|ICD9CM|PT|302.84|Sexual sadism
C0036916|ICD9CM|AB|099.9|Venereal disease NOS
C0036916|ICD9CM|PT|099.9|Venereal disease, unspecified
C0036920|ICD9CM|HT|202.2|Sezary's disease
C0036939|ICD9CM|PT|297.3|Shared psychotic disorder
C0036939|ICD9CM|AB|297.3|Shared psychotic disord
C0036974|ICD9CM|AB|785.50|Shock NOS
C0036974|ICD9CM|PT|785.50|Shock, unspecified
C0036980|ICD9CM|AB|785.51|Cardiogenic shock
C0036980|ICD9CM|PT|785.51|Cardiogenic shock
C0036983|ICD9CM|AB|785.52|Septic shock
C0036983|ICD9CM|PT|785.52|Septic shock
C0036986|ICD9CM|AB|958.4|Traumatic shock
C0036986|ICD9CM|PT|958.4|Traumatic shock
C0037005|ICD9CM|HT|831|Dislocation of shoulder
C0037023|ICD9CM|AB|527.2|Sialoadenitis
C0037023|ICD9CM|PT|527.2|Sialoadenitis
C0037054|ICD9CM|AB|282.5|Sickle-cell trait
C0037054|ICD9CM|PT|282.5|Sickle-cell trait
C0037116|ICD9CM|PT|502|Pneumoconiosis due to other silica or silicates
C0037116|ICD9CM|AB|502|Silica pneumocon NEC
C0037158|ICD9CM|HT|240|Simple and unspecified goiter
C0037221|ICD9CM|AB|759.3|Situs inversus
C0037221|ICD9CM|PT|759.3|Situs inversus
C0037304|ICD9CM|HT|800-804.99|FRACTURE OF SKULL
C0037315|ICD9CM|AB|780.57|Sleep apnea NOS
C0037315|ICD9CM|PT|780.57|Unspecified sleep apnea
C0037317|ICD9CM|HT|780.5|Sleep disturbances
C0037317|ICD9CM|AB|780.50|Sleep disturbance NOS
C0037317|ICD9CM|PT|780.50|Sleep disturbance, unspecified
C0037354|ICD9CM|HT|050|Smallpox
C0037354|ICD9CM|AB|050.9|Smallpox NOS
C0037354|ICD9CM|PT|050.9|Smallpox, unspecified
C0037358|ICD9CM|AB|050.2|Modified smallpox
C0037358|ICD9CM|PT|050.2|Modified smallpox
C0037393|ICD9CM|AB|E007.5|Soccer
C0037393|ICD9CM|PT|E007.5|Activities involving soccer
C0037448|ICD9CM|HT|312.2|Socialized conduct disorder
C0037448|ICD9CM|PT|312.20|Socialized conduct disorder, unspecified
C0037448|ICD9CM|AB|312.20|Social conduct dis-unsp
C0037619|ICD9CM|AB|610.0|Solitary cyst of breast
C0037619|ICD9CM|PT|610.0|Solitary cyst of breast
C0037646|ICD9CM|HT|94.2|Psychiatric somatotherapy
C0037650|ICD9CM|HT|300.8|Somatoform disorders
C0037753|ICD9CM|AB|123.5|Sparganosis
C0037753|ICD9CM|PT|123.5|Sparganosis [larval diphyllobothriasis]
C0037763|ICD9CM|AB|728.85|Spasm of muscle
C0037763|ICD9CM|PT|728.85|Spasm of muscle
C0037769|ICD9CM|HT|345.6|Infantile spasms
C0037773|ICD9CM|PT|334.1|Hereditary spastic paraplegia
C0037773|ICD9CM|AB|334.1|Hered spastic paraplegia
C0037785|ICD9CM|HT|315|Specific delays in development
C0037856|ICD9CM|HT|608.2|Torsion of testis
C0037856|ICD9CM|AB|608.20|Torsion of testis NOS
C0037856|ICD9CM|PT|608.20|Torsion of testis, unspecified
C0037859|ICD9CM|AB|608.1|Spermatocele
C0037859|ICD9CM|PT|608.1|Spermatocele
C0037889|ICD9CM|AB|282.0|Hereditary spherocytosis
C0037889|ICD9CM|PT|282.0|Hereditary spherocytosis
C0037928|ICD9CM|AB|336.9|Spinal cord disease NOS
C0037928|ICD9CM|PT|336.9|Unspecified disease of spinal cord
C0037932|ICD9CM|HT|737|Curvature of spine
C0037935|ICD9CM|HT|81.0|Spinal fusion
C0037935|ICD9CM|AB|81.00|Spinal fusion NOS
C0037935|ICD9CM|PT|81.00|Spinal fusion, not otherwise specified
C0037944|ICD9CM|AB|724.00|Spinal stenosis NOS
C0037944|ICD9CM|PT|724.00|Spinal stenosis, unspecified region
C0037947|ICD9CM|HT|724.0|Spinal stenosis, other than cervical
C0037952|ICD9CM|HT|334|Spinocerebellar disease
C0037952|ICD9CM|PT|334.9|Spinocerebellar disease, unspecified
C0037952|ICD9CM|AB|334.9|Spinocerebellar dis NOS
C0037974|ICD9CM|PT|104.9|Spirochetal infection, unspecified
C0037974|ICD9CM|AB|104.9|Spirochetal infect NOS
C0037997|ICD9CM|AB|289.50|Spleen disease NOS
C0037997|ICD9CM|PT|289.50|Disease of spleen, unspecified
C0038002|ICD9CM|AB|789.2|Splenomegaly
C0038002|ICD9CM|PT|789.2|Splenomegaly
C0038006|ICD9CM|PT|41.95|Repair and plastic operations on spleen
C0038006|ICD9CM|AB|41.95|Repair of spleen
C0038012|ICD9CM|PT|720.9|Unspecified inflammatory spondylopathy
C0038012|ICD9CM|AB|720.9|Inflam spondylopathy NOS
C0038013|ICD9CM|AB|720.0|Ankylosing spondylitis
C0038013|ICD9CM|PT|720.0|Ankylosing spondylitis
C0038017|ICD9CM|AB|756.12|Spondylolisthesis
C0038017|ICD9CM|PT|756.12|Spondylolisthesis
C0038019|ICD9CM|HT|721.9|Spondylosis of unspecified site
C0038034|ICD9CM|AB|117.1|Sporotrichosis
C0038034|ICD9CM|PT|117.1|Sporotrichosis
C0038041|ICD9CM|AB|082.0|Spotted fevers
C0038041|ICD9CM|PT|082.0|Spotted fevers
C0038048|ICD9CM|HT|840-848.99|SPRAINS AND STRAINS OF JOINTS AND ADJACENT MUSCLES
C0038054|ICD9CM|AB|579.1|Tropical sprue
C0038054|ICD9CM|PT|579.1|Tropical sprue
C0038150|ICD9CM|HT|19.1|Stapedectomy
C0038153|ICD9CM|AB|19.0|Stapes mobilization
C0038153|ICD9CM|PT|19.0|Stapes mobilization
C0038157|ICD9CM|PT|008.41|Intestinal infection due to staphylococcus
C0038157|ICD9CM|AB|008.41|Staphylococc enteritis
C0038159|ICD9CM|PT|005.0|Staphylococcal food poisoning
C0038159|ICD9CM|AB|005.0|Staph food poisoning
C0038165|ICD9CM|AB|695.81|Ritter's disease
C0038165|ICD9CM|PT|695.81|Ritter's disease
C0038218|ICD9CM|PT|493.91|Asthma, unspecified type, with status asthmaticus
C0038218|ICD9CM|AB|493.91|Asthma w status asthmat
C0038273|ICD9CM|PT|307.3|Stereotypic movement disorder
C0038273|ICD9CM|AB|307.3|Stereotypic movement dis
C0038325|ICD9CM|PT|695.13|Stevens-Johnson syndrome
C0038325|ICD9CM|AB|695.13|Stevens-Johnson syndrome
C0038355|ICD9CM|AB|537.1|Gastric diverticulum
C0038355|ICD9CM|PT|537.1|Gastric diverticulum
C0038358|ICD9CM|HT|531|Gastric ulcer
C0038363|ICD9CM|AB|528.2|Oral aphthae
C0038363|ICD9CM|PT|528.2|Oral aphthae
C0038379|ICD9CM|AB|378.30|Heterotropia NOS
C0038379|ICD9CM|PT|378.30|Heterotropia, unspecified
C0038380|ICD9CM|HT|378|Strabismus and other disorders of binocular eye movements
C0038436|ICD9CM|PT|309.81|Posttraumatic stress disorder
C0038436|ICD9CM|AB|309.81|Posttraumatic stress dis
C0038437|ICD9CM|PT|625.6|Stress incontinence, female
C0038437|ICD9CM|AB|625.6|Fem stress incontinence
C0038449|ICD9CM|AB|447.1|Stricture of artery
C0038449|ICD9CM|PT|447.1|Stricture of artery
C0038450|ICD9CM|AB|786.1|Stridor
C0038450|ICD9CM|PT|786.1|Stridor
C0038463|ICD9CM|AB|127.2|Strongyloidiasis
C0038463|ICD9CM|PT|127.2|Strongyloidiasis
C0038522|ICD9CM|PT|046.2|Subacute sclerosing panencephalitis
C0038522|ICD9CM|AB|046.2|Subac scleros panenceph
C0038525|ICD9CM|AB|430|Subarachnoid hemorrhage
C0038525|ICD9CM|PT|430|Subarachnoid hemorrhage
C0038531|ICD9CM|PT|435.2|Subclavian steal syndrome
C0038531|ICD9CM|AB|435.2|Subclavian steal syndrom
C0038644|ICD9CM|PT|798.0|Sudden infant death syndrome
C0038644|ICD9CM|AB|798.0|Sudden infant death synd
C0038662|ICD9CM|PT|E953.9|Suicide and self-inflicted injury by unspecified means
C0038662|ICD9CM|PT|E958.9|Suicide and self-inflicted injury by unspecified means
C0038662|ICD9CM|AB|E958.9|Injury-NOS
C0038662|ICD9CM|AB|E953.9|Injury-strang/suff NOS
C0038814|ICD9CM|AB|692.71|Sunburn
C0038814|ICD9CM|PT|692.71|Sunburn
C0038824|ICD9CM|PT|918.1|Superficial injury of cornea
C0038824|ICD9CM|AB|918.1|Superficial inj cornea
C0038843|ICD9CM|PT|V22.1|Supervision of other normal pregnancy
C0038843|ICD9CM|AB|V22.1|Supervis oth normal preg
C0038897|ICD9CM|HT|35-39.99|OPERATIONS ON THE CARDIOVASCULAR SYSTEM
C0038898|ICD9CM|HT|42-54.99|OPERATIONS ON THE DIGESTIVE SYSTEM
C0038900|ICD9CM|HT|06-07.99|OPERATIONS ON THE ENDOCRINE SYSTEM
C0038902|ICD9CM|HT|65-71.99|OPERATIONS ON THE FEMALE GENITAL ORGANS
C0038986|ICD9CM|PT|705.9|Unspecified disorder of sweat glands
C0038986|ICD9CM|HT|705|Disorders of sweat glands
C0038986|ICD9CM|AB|705.9|Sweat gland disorder NOS
C0038992|ICD9CM|AB|078.2|Sweating fever
C0038992|ICD9CM|PT|078.2|Sweating fever
C0039003|ICD9CM|AB|E002.0|Swimming
C0039003|ICD9CM|PT|E002.0|Activities involving swimming
C0039038|ICD9CM|HT|05.2|Sympathectomy
C0039043|ICD9CM|PT|05.31|Injection of anesthetic into sympathetic nerve for analgesia
C0039043|ICD9CM|AB|05.31|Anesth inject symp nerve
C0039056|ICD9CM|AB|55.85|Symphysiotomy
C0039056|ICD9CM|PT|55.85|Symphysiotomy for horseshoe kidney
C0039070|ICD9CM|AB|780.2|Syncope and collapse
C0039070|ICD9CM|PT|780.2|Syncope and collapse
C0039075|ICD9CM|HT|755.1|Syndactyly
C0039104|ICD9CM|HT|727.0|Synovitis and tenosynovitis
C0039104|ICD9CM|AB|727.00|Synovitis NOS
C0039104|ICD9CM|PT|727.00|Synovitis and tenosynovitis, unspecified
C0039128|ICD9CM|AB|097.9|Syphilis NOS
C0039128|ICD9CM|PT|097.9|Syphilis, unspecified
C0039130|ICD9CM|HT|093|Cardiovascular syphilis
C0039130|ICD9CM|PT|093.9|Cardiovascular syphilis, unspecified
C0039130|ICD9CM|AB|093.9|Cardiovascular syph NOS
C0039131|ICD9CM|HT|090|Congenital syphilis
C0039131|ICD9CM|AB|090.9|Congenital syphilis NOS
C0039131|ICD9CM|PT|090.9|Congenital syphilis, unspecified
C0039133|ICD9CM|AB|097.1|Latent syphilis NOS
C0039133|ICD9CM|PT|097.1|Latent syphilis, unspecified
C0039145|ICD9CM|PT|336.0|Syringomyelia and syringobulbia
C0039145|ICD9CM|AB|336.0|Syringomyelia
C0039223|ICD9CM|AB|094.0|Tabes dorsalis
C0039223|ICD9CM|PT|094.0|Tabes dorsalis
C0039231|ICD9CM|AB|785.0|Tachycardia NOS
C0039231|ICD9CM|PT|785.0|Tachycardia, unspecified
C0039236|ICD9CM|PT|427.2|Paroxysmal tachycardia, unspecified
C0039236|ICD9CM|AB|427.2|Parox tachycardia NOS
C0039254|ICD9CM|AB|123.3|Taeniasis NOS
C0039254|ICD9CM|PT|123.3|Taeniasis, unspecified
C0039263|ICD9CM|AB|446.7|Takayasu's disease
C0039263|ICD9CM|PT|446.7|Takayasu's disease
C0039319|ICD9CM|AB|355.5|Tarsal tunnel syndrome
C0039319|ICD9CM|PT|355.5|Tarsal tunnel syndrome
C0039437|ICD9CM|AB|520.7|Teething syndrome
C0039437|ICD9CM|PT|520.7|Teething syndrome
C0039445|ICD9CM|PT|448.0|Hereditary hemorrhagic telangiectasia
C0039445|ICD9CM|AB|448.0|Heredit hemorr telangiec
C0039483|ICD9CM|AB|446.5|Giant cell arteritis
C0039483|ICD9CM|PT|446.5|Giant cell arteritis
C0039492|ICD9CM|AB|31.1|Temporary tracheostomy
C0039492|ICD9CM|PT|31.1|Temporary tracheostomy
C0039494|ICD9CM|HT|524.6|Temporomandibular joint disorders
C0039494|ICD9CM|PT|524.60|Temporomandibular joint disorders, unspecified
C0039494|ICD9CM|AB|524.60|TMJ disorders NOS
C0039516|ICD9CM|AB|726.32|Lateral epicondylitis
C0039516|ICD9CM|PT|726.32|Lateral epicondylitis
C0039585|ICD9CM|PT|259.51|Androgen insensitivity syndrome
C0039585|ICD9CM|HT|259.5|Androgen insensitivity syndrome
C0039585|ICD9CM|AB|259.51|Androgen insensitvty syn
C0039613|ICD9CM|AB|366.42|Tetanic cataract
C0039613|ICD9CM|PT|366.42|Tetanic cataract
C0039614|ICD9CM|AB|037|Tetanus
C0039614|ICD9CM|PT|037|Tetanus
C0039621|ICD9CM|AB|781.7|Tetany
C0039621|ICD9CM|PT|781.7|Tetany
C0039685|ICD9CM|AB|745.2|Tetralogy of fallot
C0039685|ICD9CM|PT|745.2|Tetralogy of fallot
C0039730|ICD9CM|HT|282.4|Thalassemias
C0039730|ICD9CM|AB|282.40|Thalassemia, unspecified
C0039730|ICD9CM|PT|282.40|Thalassemia, unspecified
C0039788|ICD9CM|PT|96.25|Therapeutic distention of bladder
C0039788|ICD9CM|AB|96.25|Therapeut distent bladd
C0039804|ICD9CM|PT|12.62|Thermocauterization of sclera with iridectomy
C0039804|ICD9CM|AB|12.62|Thermcaut scler w iridec
C0039810|ICD9CM|HT|88.8|Thermography
C0039812|ICD9CM|PT|88.89|Thermography of other sites
C0039812|ICD9CM|AB|88.89|Thermography NEC
C0039988|ICD9CM|AB|33.34|Thoracoplasty
C0039988|ICD9CM|PT|33.34|Thoracoplasty
C0039989|ICD9CM|PT|34.21|Transpleural thoracoscopy
C0039989|ICD9CM|AB|34.21|Transpleura thoracoscopy
C0039991|ICD9CM|AB|34.01|Incision of chest wall
C0039991|ICD9CM|PT|34.01|Incision of chest wall
C0040021|ICD9CM|PT|443.1|Thromboangiitis obliterans [Buerger's disease]
C0040021|ICD9CM|AB|443.1|Thromboangiit obliterans
C0040028|ICD9CM|PT|238.71|Essential thrombocythemia
C0040028|ICD9CM|AB|238.71|Essntial thrombocythemia
C0040034|ICD9CM|AB|287.5|Thrombocytopenia NOS
C0040034|ICD9CM|PT|287.5|Thrombocytopenia, unspecified
C0040038|ICD9CM|AB|453.9|Venous thrombosis NOS
C0040038|ICD9CM|PT|453.9|Other venous embolism and thrombosis of unspecified site
C0040071|ICD9CM|HT|07.8|Thymectomy
C0040071|ICD9CM|AB|07.80|Thymectomy NOS
C0040071|ICD9CM|PT|07.80|Thymectomy, not otherwise specified
C0040128|ICD9CM|PT|246.9|Unspecified disorder of thyroid
C0040128|ICD9CM|AB|246.9|Disorder of thyroid NOS
C0040128|ICD9CM|HT|240-246.99|DISORDERS OF THYROID GLAND
C0040147|ICD9CM|HT|245|Thyroiditis
C0040147|ICD9CM|AB|245.9|Thyroiditis NOS
C0040147|ICD9CM|PT|245.9|Thyroiditis, unspecified
C0040149|ICD9CM|AB|245.1|Subacute thyroiditis
C0040149|ICD9CM|PT|245.1|Subacute thyroiditis
C0040156|ICD9CM|HT|242|Thyrotoxicosis with or without goiter
C0040188|ICD9CM|AB|307.20|Tic disorder NOS
C0040188|ICD9CM|HT|307.2|Tics
C0040188|ICD9CM|PT|307.20|Tic disorder, unspecified
C0040199|ICD9CM|AB|066.1|Tick-borne fever
C0040199|ICD9CM|PT|066.1|Tick-borne fever
C0040213|ICD9CM|AB|733.6|Tietze's disease
C0040213|ICD9CM|PT|733.6|Tietze's disease
C0040249|ICD9CM|AB|111.2|Tinea blanca
C0040249|ICD9CM|PT|111.2|Tinea blanca
C0040259|ICD9CM|AB|110.4|Dermatophytosis of foot
C0040259|ICD9CM|PT|110.4|Dermatophytosis of foot
C0040262|ICD9CM|AB|111.0|Pityriasis versicolor
C0040262|ICD9CM|PT|111.0|Pityriasis versicolor
C0040264|ICD9CM|HT|388.3|Tinnitus
C0040264|ICD9CM|AB|388.30|Tinnitus NOS
C0040264|ICD9CM|PT|388.30|Tinnitus, unspecified
C0040335|ICD9CM|AB|V15.82|History of tobacco use
C0040335|ICD9CM|PT|V15.82|Personal history of tobacco use
C0040336|ICD9CM|AB|305.1|Tobacco use disorder
C0040336|ICD9CM|PT|305.1|Tobacco use disorder
C0040409|ICD9CM|PT|529.9|Unspecified condition of the tongue
C0040409|ICD9CM|AB|529.9|Tongue disorder NOS
C0040412|ICD9CM|AB|529.5|Plicated tongue
C0040412|ICD9CM|PT|529.5|Plicated tongue
C0040416|ICD9CM|AB|379.46|Tonic pupillary reaction
C0040416|ICD9CM|PT|379.46|Tonic pupillary reaction
C0040420|ICD9CM|AB|89.11|Tonometry
C0040420|ICD9CM|PT|89.11|Tonometry
C0040423|ICD9CM|AB|28.2|Tonsillectomy
C0040423|ICD9CM|PT|28.2|Tonsillectomy without adenoidectomy
C0040428|ICD9CM|HT|521.2|Abrasion of teeth
C0040433|ICD9CM|AB|524.31|Crowding of teeth
C0040433|ICD9CM|PT|524.31|Crowding of teeth
C0040436|ICD9CM|HT|521.3|Erosion of teeth
C0040440|ICD9CM|HT|23.1|Surgical removal of tooth
C0040451|ICD9CM|HT|521.4|Pathological tooth resorption
C0040457|ICD9CM|AB|520.1|Supernumerary teeth
C0040457|ICD9CM|PT|520.1|Supernumerary teeth
C0040485|ICD9CM|AB|723.5|Torticollis NOS
C0040485|ICD9CM|PT|723.5|Torticollis, unspecified
C0040507|ICD9CM|AB|50.4|Total hepatectomy
C0040507|ICD9CM|PT|50.4|Total hepatectomy
C0040508|ICD9CM|AB|81.51|Total hip replacement
C0040508|ICD9CM|PT|81.51|Total hip replacement
C0040511|ICD9CM|AB|52.6|Total pancreatectomy
C0040511|ICD9CM|PT|52.6|Total pancreatectomy
C0040517|ICD9CM|AB|307.23|Tourette's disorder
C0040517|ICD9CM|PT|307.23|Tourette's disorder
C0040528|ICD9CM|PT|988.2|Toxic effect of berries and other plants eaten as food
C0040528|ICD9CM|AB|988.2|Tox eff berry/plant NEC
C0040531|ICD9CM|PT|985.8|Toxic effect of other specified metals
C0040531|ICD9CM|AB|985.8|Toxic effect metals NEC
C0040533|ICD9CM|PT|989.5|Toxic effect of venom
C0040533|ICD9CM|AB|989.5|Toxic effect venom
C0040543|ICD9CM|PT|91.85|Microscopic examination of specimen from other site, toxicology
C0040543|ICD9CM|AB|91.85|Toxicology NEC
C0040553|ICD9CM|AB|128.0|Toxocariasis
C0040553|ICD9CM|PT|128.0|Toxocariasis
C0040558|ICD9CM|HT|130|Toxoplasmosis
C0040558|ICD9CM|AB|130.9|Toxoplasmosis NOS
C0040558|ICD9CM|PT|130.9|Toxoplasmosis, unspecified
C0040585|ICD9CM|PT|67.61|Suture of laceration of cervix
C0040585|ICD9CM|AB|67.61|Suture cervical lacerat
C0040588|ICD9CM|PT|530.84|Tracheoesophageal fistula
C0040588|ICD9CM|AB|530.84|Tracheoesophageal fstula
C0040592|ICD9CM|HT|076|Trachoma
C0040592|ICD9CM|AB|076.9|Trachoma NOS
C0040592|ICD9CM|PT|076.9|Trachoma, unspecified
C0040630|ICD9CM|PT|302.50|Trans-sexualism with unspecified sexual history
C0040630|ICD9CM|AB|302.50|Trans-sexualism NOS
C0040694|ICD9CM|PT|99.07|Transfusion of other serum
C0040694|ICD9CM|AB|99.07|Serum transfusion NEC
C0040701|ICD9CM|HT|309|Adjustment reaction
C0040701|ICD9CM|AB|309.9|Adjustment reaction NOS
C0040701|ICD9CM|PT|309.9|Unspecified adjustment reaction
C0040702|ICD9CM|AB|307.21|Transient tic disorder
C0040702|ICD9CM|PT|307.21|Transient tic disorder
C0040750|ICD9CM|PT|V42.4|Bone replaced by transplant
C0040750|ICD9CM|AB|V42.4|Bone transplant status
C0040761|ICD9CM|HT|745.1|Transposition of great vessels
C0040761|ICD9CM|PT|745.10|Complete transposition of great vessels
C0040761|ICD9CM|AB|745.10|Compl transpos great ves
C0040765|ICD9CM|HT|302.5|Trans-sexualism
C0040769|ICD9CM|PT|57.0|Transurethral clearance of bladder
C0040769|ICD9CM|AB|57.0|Tu bladder clearance
C0040771|ICD9CM|HT|60.2|Transurethral prostatectomy
C0040774|ICD9CM|AB|302.3|Transvestic fetishism
C0040774|ICD9CM|PT|302.3|Transvestic fetishism
C0040793|ICD9CM|AB|958.5|Traumatic anuria
C0040793|ICD9CM|PT|958.5|Traumatic anuria
C0040798|ICD9CM|PT|728.12|Traumatic myositis ossificans
C0040798|ICD9CM|AB|728.12|Traum myositis ossifican
C0040799|ICD9CM|PT|958.7|Traumatic subcutaneous emphysema
C0040799|ICD9CM|AB|958.7|Traum subcutan emphysema
C0040820|ICD9CM|AB|121.9|Trematode infection NOS
C0040820|ICD9CM|PT|121.9|Trematode infection, unspecified
C0040830|ICD9CM|AB|083.1|Trench fever
C0040830|ICD9CM|PT|083.1|Trench fever
C0040896|ICD9CM|AB|124|Trichinosis
C0040896|ICD9CM|PT|124|Trichinosis
C0040921|ICD9CM|HT|131|Trichomoniasis
C0040921|ICD9CM|AB|131.9|Trichomoniasis NOS
C0040921|ICD9CM|PT|131.9|Trichomoniasis, unspecified
C0040926|ICD9CM|PT|131.8|Trichomoniasis of other specified sites
C0040926|ICD9CM|AB|131.8|Trichomoniasis NEC
C0040928|ICD9CM|HT|131.0|Urogenital trichomoniasis
C0040928|ICD9CM|PT|131.00|Urogenital trichomoniasis, unspecified
C0040928|ICD9CM|AB|131.00|Urogenital trichomon NOS
C0040948|ICD9CM|AB|127.6|Trichostrongyliasis
C0040948|ICD9CM|PT|127.6|Trichostrongyliasis
C0040997|ICD9CM|AB|350.1|Trigeminal neuralgia
C0040997|ICD9CM|PT|350.1|Trigeminal neuralgia
C0041188|ICD9CM|AB|040.81|Tropical pyomyositis
C0041188|ICD9CM|PT|040.81|Tropical pyomyositis
C0041207|ICD9CM|AB|745.0|Common truncus
C0041207|ICD9CM|PT|745.0|Common truncus
C0041227|ICD9CM|HT|086|Trypanosomiasis
C0041227|ICD9CM|AB|086.9|Trypanosomiasis NOS
C0041227|ICD9CM|PT|086.9|Trypanosomiasis, unspecified
C0041228|ICD9CM|AB|086.5|African trypanosoma NOS
C0041228|ICD9CM|PT|086.5|African trypanosomiasis, unspecified
C0041232|ICD9CM|AB|086.3|Gambian trypanosomiasis
C0041232|ICD9CM|PT|086.3|Gambian trypanosomiasis
C0041233|ICD9CM|PT|086.4|Rhodesian trypanosomiasis
C0041233|ICD9CM|AB|086.4|Rhodesian trypanosomias
C0041296|ICD9CM|HT|010-018.99|TUBERCULOSIS
C0041300|ICD9CM|HT|017|Tuberculosis of other organs
C0041301|ICD9CM|HT|017.9|Tuberculosis of other specified organs
C0041301|ICD9CM|AB|017.90|TB of organ NEC-unspec
C0041301|ICD9CM|PT|017.90|Tuberculosis of other specified organs, unspecified
C0041315|ICD9CM|HT|012.3|Tuberculous laryngitis
C0041318|ICD9CM|HT|013.0|Tuberculous meningitis
C0041318|ICD9CM|AB|013.00|TB meningitis-unspec
C0041318|ICD9CM|PT|013.00|Tuberculous meningitis, unspecified
C0041321|ICD9CM|HT|018|Miliary tuberculosis
C0041321|ICD9CM|HT|018.9|Unspecified miliary tuberculosis
C0041321|ICD9CM|AB|018.90|Miliary TB NOS-unspec
C0041321|ICD9CM|PT|018.90|Miliary tuberculosis, unspecified, unspecified
C0041322|ICD9CM|HT|017.3|Tuberculosis of eye
C0041322|ICD9CM|AB|017.30|TB of eye-unspec
C0041322|ICD9CM|PT|017.30|Tuberculosis of eye, unspecified
C0041324|ICD9CM|HT|015.9|Tuberculosis of unspecified bones and joints
C0041324|ICD9CM|HT|015|Tuberculosis of bones and joints
C0041325|ICD9CM|HT|014.0|Tuberculous peritonitis
C0041326|ICD9CM|HT|012.0|Tuberculous pleurisy
C0041326|ICD9CM|AB|012.00|TB pleurisy-unspec
C0041326|ICD9CM|PT|012.00|Tuberculous pleurisy, unspecified
C0041327|ICD9CM|HT|011|Pulmonary tuberculosis
C0041327|ICD9CM|HT|011.9|Unspecified pulmonary tuberculosis
C0041327|ICD9CM|AB|011.90|Pulmonary TB NOS-unspec
C0041327|ICD9CM|PT|011.90|Pulmonary tuberculosis, unspecified, unspecified
C0041328|ICD9CM|HT|016.0|Tuberculosis of kidney
C0041328|ICD9CM|AB|016.00|TB of kidney-unspec
C0041328|ICD9CM|PT|016.00|Tuberculosis of kidney, unspecified
C0041330|ICD9CM|AB|015.00|TB of vertebra-unspec
C0041330|ICD9CM|HT|015.0|Tuberculosis of vertebral column
C0041330|ICD9CM|PT|015.00|Tuberculosis of vertebral column, unspecified
C0041331|ICD9CM|HT|017.7|Tuberculosis of spleen
C0041332|ICD9CM|HT|016.3|Tuberculosis of other urinary organs
C0041333|ICD9CM|HT|016|Tuberculosis of genitourinary system
C0041333|ICD9CM|HT|016.9|Genitourinary tuberculosis, unspecified
C0041336|ICD9CM|HT|011.4|Tuberculous fibrosis of lung
C0041336|ICD9CM|AB|011.40|TB lung fibrosis-unspec
C0041336|ICD9CM|PT|011.40|Tuberculous fibrosis of lung, unspecified
C0041341|ICD9CM|AB|759.5|Tuberous sclerosis
C0041341|ICD9CM|PT|759.5|Tuberous sclerosis
C0041351|ICD9CM|HT|021|Tularemia
C0041351|ICD9CM|AB|021.9|Tularemia NOS
C0041351|ICD9CM|PT|021.9|Unspecified tularemia
C0041364|ICD9CM|PT|277.88|Tumor lysis syndrome
C0041364|ICD9CM|AB|277.88|Tumor lysis syndrome
C0041423|ICD9CM|HT|V33|Twin birth, unspecified whether mate liveborn or stillborn
C0041428|ICD9CM|AB|759.4|Conjoined twins
C0041428|ICD9CM|PT|759.4|Conjoined twins
C0041466|ICD9CM|AB|002.0|Typhoid fever
C0041466|ICD9CM|PT|002.0|Typhoid fever
C0041471|ICD9CM|AB|081.9|Typhus NOS
C0041471|ICD9CM|PT|081.9|Typhus, unspecified
C0041472|ICD9CM|PT|081.0|Murine (endemic) typhus
C0041472|ICD9CM|AB|081.0|Murine typhus
C0041473|ICD9CM|PT|080|Louse-borne (epidemic) typhus
C0041473|ICD9CM|AB|080|Louse-borne typhus
C0041618|ICD9CM|HT|88.7|Diagnostic ultrasound
C0041620|ICD9CM|HT|00.0|Therapeutic ultrasound
C0041626|ICD9CM|PT|99.82|Ultraviolet light therapy
C0041626|ICD9CM|AB|99.82|Ultraviolet light therap
C0041636|ICD9CM|PT|553.1|Umbilical hernia without mention of obstruction or gangrene
C0041636|ICD9CM|AB|553.1|Umbilical hernia
C0041665|ICD9CM|HT|312.0|Undersocialized conduct disorder, aggressive type
C0041667|ICD9CM|AB|783.22|Underweight
C0041667|ICD9CM|PT|783.22|Underweight
C0041672|ICD9CM|PT|300.82|Undifferentiated somatoform disorder
C0041672|ICD9CM|AB|300.82|Undiff somatoform disrdr
C0041684|ICD9CM|AB|07.22|Unilateral adrenalectomy
C0041684|ICD9CM|PT|07.22|Unilateral adrenalectomy
C0041685|ICD9CM|PT|85.47|Unilateral extended radical mastectomy
C0041685|ICD9CM|AB|85.47|Unil ext rad mastectomy
C0041687|ICD9CM|HT|65.3|Unilateral oophorectomy
C0041688|ICD9CM|PT|553.00|Femoral hernia without mention of obstruction of gangrene, unilateral or unspecified(not specified as recurrent)
C0041688|ICD9CM|AB|553.00|Unilat femoral hernia
C0041690|ICD9CM|PT|85.45|Unilateral radical mastectomy
C0041690|ICD9CM|AB|85.45|Unilat radical mastectom
C0041691|ICD9CM|PT|53.00|Unilateral repair of inguinal hernia, not otherwise specified
C0041691|ICD9CM|AB|53.00|Unilat ing hern rep NOS
C0041692|ICD9CM|HT|65.4|Unilateral salpingo-oophorectomy
C0041782|ICD9CM|AB|281.9|Deficiency anemia NOS
C0041782|ICD9CM|PT|281.9|Unspecified deficiency anemia
C0041784|ICD9CM|PT|736.00|Unspecified deformity of forearm, excluding fingers
C0041784|ICD9CM|AB|736.00|Forearm deformity NOS
C0041785|ICD9CM|HT|710|Diffuse diseases of connective tissue
C0041785|ICD9CM|PT|710.9|Unspecified diffuse connective tissue disease
C0041785|ICD9CM|AB|710.9|Diff connect tis dis NOS
C0041792|ICD9CM|HT|077.9|Unspecified diseases of conjunctiva due to viruses and Chlamydiae
C0041806|ICD9CM|PT|279.9|Unspecified disorder of immune mechanism
C0041806|ICD9CM|HT|279|Disorders involving the immune mechanism
C0041806|ICD9CM|AB|279.9|Immune mechanism dis NOS
C0041825|ICD9CM|PT|384.9|Unspecified disorder of tympanic membrane
C0041825|ICD9CM|AB|384.9|Dis tympanic memb NOS
C0041827|ICD9CM|PT|626.9|Unspecified disorders of menstruation and other abnormal bleeding from female genital tract
C0041827|ICD9CM|HT|626|Disorders of menstruation and other abnormal bleeding from female genital tract
C0041827|ICD9CM|AB|626.9|Menstrual disorder NOS
C0041831|ICD9CM|PT|E947.9|Unspecified drug or medicinal substance causing adverse effects in therapeutic use
C0041831|ICD9CM|AB|E947.9|Adv eff medicinal NOS
C0041834|ICD9CM|PT|695.9|Unspecified erythematous condition
C0041834|ICD9CM|HT|695|Erythematous conditions
C0041834|ICD9CM|AB|695.9|Erythematous cond NOS
C0041841|ICD9CM|HT|535.5|Unspecified gastritis and gastroduodenitis
C0041844|ICD9CM|AB|455.6|Hemorrhoids NOS
C0041844|ICD9CM|PT|455.6|Unspecified hemorrhoids without mention of complication
C0041847|ICD9CM|PT|701.9|Unspecified hypertrophic and atrophic conditions of skin
C0041847|ICD9CM|AB|701.9|Skin hypertro/atroph NOS
C0041849|ICD9CM|PT|136.9|Unspecified infectious and parasitic diseases
C0041849|ICD9CM|HT|001-139.99|INFECTIOUS AND PARASITIC DISEASES
C0041849|ICD9CM|AB|136.9|Infect/parasite dis NOS
C0041857|ICD9CM|PT|300.9|Unspecified nonpsychotic mental disorder
C0041857|ICD9CM|AB|300.9|Nonpsychotic disord NOS
C0041862|ICD9CM|PT|310.9|Unspecified nonpsychotic mental disorder following organic brain damage
C0041862|ICD9CM|AB|310.9|Nonpsychot brain syn NOS
C0041866|ICD9CM|PT|V42.9|Unspecified organ or tissue replaced by transplant
C0041866|ICD9CM|HT|V42|Organ or tissue replaced by transplant
C0041866|ICD9CM|AB|V42.9|Transplant status NOS
C0041876|ICD9CM|PT|306.9|Unspecified psychophysiological malfunction
C0041876|ICD9CM|AB|306.9|Psychogenic disorder NOS
C0041880|ICD9CM|PT|V65.9|Unspecified reason for consultation
C0041880|ICD9CM|AB|V65.9|Reason for consult NOS
C0041881|ICD9CM|PT|506.9|Unspecified respiratory conditions due to fumes and vapors
C0041881|ICD9CM|AB|506.9|Fum/vapor resp cond NOS
C0041887|ICD9CM|PT|848.9|Unspecified site of sprain and strain
C0041887|ICD9CM|AB|848.9|Sprain NOS
C0041889|ICD9CM|PT|625.9|Unspecified symptom associated with female genital organs
C0041889|ICD9CM|AB|625.9|Fem genital symptoms NOS
C0041893|ICD9CM|PT|553.20|Ventral, unspecified, hernia without mention of obstruction or gangrene
C0041893|ICD9CM|AB|553.20|Ventral hernia NOS
C0041952|ICD9CM|AB|592.1|Calculus of ureter
C0041952|ICD9CM|PT|592.1|Calculus of ureter
C0041953|ICD9CM|AB|59.8|Ureteral catheterization
C0041953|ICD9CM|PT|59.8|Ureteral catheterization
C0041970|ICD9CM|AB|599.1|Urethral fistula
C0041970|ICD9CM|PT|599.1|Urethral fistula
C0041979|ICD9CM|PT|58.41|Suture of laceration of urethra
C0041979|ICD9CM|AB|58.41|Suture urethral lacerat
C0042023|ICD9CM|AB|788.41|Urinary frequency
C0042023|ICD9CM|PT|788.41|Urinary frequency
C0042024|ICD9CM|HT|788.3|Urinary incontinence
C0042024|ICD9CM|AB|788.30|Urinary incontinence NOS
C0042024|ICD9CM|PT|788.30|Urinary incontinence, unspecified
C0042029|ICD9CM|PT|599.0|Urinary tract infection, site not specified
C0042029|ICD9CM|AB|599.0|Urin tract infection NOS
C0042033|ICD9CM|PT|619.0|Urinary-genital tract fistula, female
C0042033|ICD9CM|AB|619.0|Urin-genital fistul, fem
C0042075|ICD9CM|PT|599.9|Unspecified disorder of urethra and urinary tract
C0042075|ICD9CM|AB|599.9|Urinary tract dis NOS
C0042109|ICD9CM|HT|708|Urticaria
C0042109|ICD9CM|AB|708.9|Urticaria NOS
C0042109|ICD9CM|PT|708.9|Urticaria, unspecified
C0042131|ICD9CM|AB|621.9|Disorder of uterus NOS
C0042131|ICD9CM|PT|621.9|Unspecified disorder of uterus
C0042133|ICD9CM|HT|218|Uterine leiomyoma
C0042133|ICD9CM|AB|218.9|Uterine leiomyoma NOS
C0042133|ICD9CM|PT|218.9|Leiomyoma of uterus, unspecified
C0042170|ICD9CM|AB|364.24|Vogt-koyanagi syndrome
C0042170|ICD9CM|PT|364.24|Vogt-koyanagi syndrome
C0042170|ICD9CM|AB|363.22|Harada's disease
C0042170|ICD9CM|PT|363.22|Harada's disease
C0042199|ICD9CM|PT|99.31|Vaccination against cholera
C0042199|ICD9CM|AB|99.31|Cholera vaccination
C0042200|ICD9CM|AB|99.52|Influenza vaccination
C0042200|ICD9CM|PT|99.52|Prophylactic vaccination against influenza
C0042201|ICD9CM|AB|99.45|Measles vaccination
C0042201|ICD9CM|PT|99.45|Vaccination against measles
C0042202|ICD9CM|PT|99.46|Vaccination against mumps
C0042202|ICD9CM|AB|99.46|Mumps vaccination
C0042203|ICD9CM|AB|99.37|Pertussis vaccination
C0042203|ICD9CM|PT|99.37|Vaccination against pertussis
C0042204|ICD9CM|AB|99.34|Plague vaccination
C0042204|ICD9CM|PT|99.34|Vaccination against plague
C0042205|ICD9CM|AB|99.44|Rabies vaccination
C0042205|ICD9CM|PT|99.44|Vaccination against rabies
C0042206|ICD9CM|AB|99.47|Rubella vaccination
C0042206|ICD9CM|PT|99.47|Vaccination against rubella
C0042207|ICD9CM|PT|99.42|Vaccination against smallpox
C0042207|ICD9CM|AB|99.42|Smallpox vaccination
C0042225|ICD9CM|HT|72.7|Vacuum extraction
C0042237|ICD9CM|PT|184.0|Malignant neoplasm of vagina
C0042237|ICD9CM|AB|184.0|Malign neopl vagina
C0042266|ICD9CM|AB|306.51|Psychogenic vaginismus
C0042266|ICD9CM|PT|306.51|Psychogenic vaginismus
C0042268|ICD9CM|HT|616.1|Vaginitis and vulvovaginitis
C0042268|ICD9CM|AB|616.10|Vaginitis NOS
C0042268|ICD9CM|PT|616.10|Vaginitis and vulvovaginitis, unspecified
C0042273|ICD9CM|PT|44.02|Highly selective vagotomy
C0042273|ICD9CM|AB|44.02|Highly select vagotomy
C0042275|ICD9CM|AB|44.01|Truncal vagotomy
C0042275|ICD9CM|PT|44.01|Truncal vagotomy
C0042341|ICD9CM|AB|456.4|Scrotal varices
C0042341|ICD9CM|PT|456.4|Scrotal varices
C0042347|ICD9CM|PT|454.1|Varicose veins of lower extremities with inflammation
C0042347|ICD9CM|AB|454.1|Leg varicosity w inflam
C0042370|ICD9CM|PT|372.74|Vascular abnormalities of conjunctiva
C0042370|ICD9CM|AB|372.74|Conjunctiva vasc anomaly
C0042374|ICD9CM|PT|608.83|Vascular disorders of male genital organs
C0042374|ICD9CM|AB|608.83|Male gen vascul dis NEC
C0042387|ICD9CM|AB|63.73|Vasectomy
C0042387|ICD9CM|PT|63.73|Vasectomy
C0042416|ICD9CM|AB|63.6|Vasotomy
C0042416|ICD9CM|PT|63.6|Vasotomy
C0042421|ICD9CM|AB|63.82|Postop vas reconstruct
C0042421|ICD9CM|PT|63.82|Reconstruction of surgically divided vas deferens
C0042477|ICD9CM|PT|E905.0|Venomous snakes and lizards causing poisoning and toxic reactions
C0042477|ICD9CM|AB|E905.0|Venomous snake bite
C0042478|ICD9CM|AB|E905.1|Venomous spider bite
C0042478|ICD9CM|PT|E905.1|Venomous spiders causing poisoning and toxic reactions
C0042485|ICD9CM|AB|459.81|Venous insufficiency NOS
C0042485|ICD9CM|PT|459.81|Venous (peripheral) insufficiency, unspecified
C0042505|ICD9CM|HT|553.2|Ventral hernia without mention of obstruction or gangrene
C0042510|ICD9CM|AB|427.41|Ventricular fibrillation
C0042510|ICD9CM|PT|427.41|Ventricular fibrillation
C0042517|ICD9CM|HT|02.2|Ventriculostomy
C0042548|ICD9CM|PT|078.12|Plantar wart
C0042548|ICD9CM|AB|078.12|Plantar wart
C0042568|ICD9CM|PT|435.3|Vertebrobasilar artery syndrome
C0042568|ICD9CM|AB|435.3|Vertbrobaslr artery synd
C0042580|ICD9CM|HT|593.7|Vesicoureteral reflux
C0042588|ICD9CM|AB|608.0|Seminal vesiculitis
C0042588|ICD9CM|PT|608.0|Seminal vesiculitis
C0042609|ICD9CM|PT|24.91|Extension or deepening of buccolabial or lingual sulcus
C0042609|ICD9CM|AB|24.91|Exten buccolabial/sulcus
C0042721|ICD9CM|HT|070|Viral hepatitis
C0042749|ICD9CM|AB|790.8|Viremia NOS
C0042749|ICD9CM|PT|790.8|Viremia, unspecified
C0042818|ICD9CM|AB|368.13|Visual discomfort
C0042818|ICD9CM|PT|368.13|Visual discomfort
C0042825|ICD9CM|AB|95.05|Visual field study
C0042825|ICD9CM|PT|95.05|Visual field study
C0042835|ICD9CM|PT|89.37|Vital capacity determination
C0042835|ICD9CM|AB|89.37|Vital capacity determin
C0042842|ICD9CM|HT|264|Vitamin A deficiency
C0042842|ICD9CM|AB|264.9|Vitamin A deficiency NOS
C0042842|ICD9CM|PT|264.9|Unspecified vitamin A deficiency
C0042850|ICD9CM|AB|266.9|Vitamin b deficiency NOS
C0042850|ICD9CM|PT|266.9|Unspecified vitamin B deficiency
C0042850|ICD9CM|HT|266|Deficiency of B-complex components
C0042870|ICD9CM|HT|268|Vitamin D deficiency
C0042870|ICD9CM|AB|268.9|Vitamin D deficiency NOS
C0042870|ICD9CM|PT|268.9|Unspecified vitamin D deficiency
C0042880|ICD9CM|PT|269.0|Deficiency of vitamin K
C0042880|ICD9CM|AB|269.0|Deficiency of vitamin k
C0042900|ICD9CM|AB|709.01|Vitiligo
C0042900|ICD9CM|PT|709.01|Vitiligo
C0042904|ICD9CM|AB|360.04|Vitreous abscess
C0042904|ICD9CM|PT|360.04|Vitreous abscess
C0042909|ICD9CM|AB|379.23|Vitreous hemorrhage
C0042909|ICD9CM|PT|379.23|Vitreous hemorrhage
C0042928|ICD9CM|AB|478.30|Vocal cord paralysis NOS
C0042928|ICD9CM|PT|478.30|Paralysis of vocal cords or larynx, unspecified
C0042951|ICD9CM|PT|958.6|Volkmann's ischemic contracture
C0042951|ICD9CM|AB|958.6|Volkmann's isch contract
C0042961|ICD9CM|PT|560.2|Volvulus
C0042961|ICD9CM|AB|560.2|Volvulus of intestine
C0042974|ICD9CM|PT|286.4|Von Willebrand's disease
C0042974|ICD9CM|AB|286.4|Von willebrand's disease
C0042979|ICD9CM|AB|302.82|Voyeurism
C0042979|ICD9CM|PT|302.82|Voyeurism
C0043102|ICD9CM|AB|100.0|Leptospiros icterohem
C0043102|ICD9CM|PT|100.0|Leptospirosis icterohemorrhagica
C0043116|ICD9CM|PT|335.0|Werdnig-Hoffmann disease
C0043116|ICD9CM|AB|335.0|Werdnig-hoffmann disease
C0043124|ICD9CM|HT|066.4|West Nile fever
C0043124|ICD9CM|AB|066.40|West Nile Fever NOS
C0043124|ICD9CM|PT|066.40|West Nile Fever, unspecified
C0043144|ICD9CM|AB|786.07|Wheezing
C0043144|ICD9CM|PT|786.07|Wheezing
C0043167|ICD9CM|AB|033.0|Bordetella pertussis
C0043167|ICD9CM|PT|033.0|Whooping cough due to bordetella pertussis [B. pertussis]
C0043168|ICD9CM|HT|033|Whooping cough
C0043168|ICD9CM|AB|033.9|Whooping cough NOS
C0043168|ICD9CM|PT|033.9|Whooping cough, unspecified organism
C0043170|ICD9CM|PT|033.8|Whooping cough due to other specified organism
C0043170|ICD9CM|AB|033.8|Whooping cough NEC
C0043194|ICD9CM|AB|279.12|Wiskott-aldrich syndrome
C0043194|ICD9CM|PT|279.12|Wiskott-aldrich syndrome
C0043261|ICD9CM|AB|E008.1|Wrestling
C0043261|ICD9CM|PT|E008.1|Activities involving wrestling
C0043299|ICD9CM|HT|87|Diagnostic Radiology
C0043348|ICD9CM|PT|87.36|Xerography of breast
C0043348|ICD9CM|AB|87.36|Breast xerography
C0043349|ICD9CM|AB|375.15|Tear film insuffic NOS
C0043349|ICD9CM|PT|375.15|Tear film insufficiency, unspecified
C0043384|ICD9CM|PT|059.22|Yaba monkey tumor virus
C0043384|ICD9CM|AB|059.22|Yaba monkey tumor virus
C0043388|ICD9CM|HT|102|Yaws
C0043388|ICD9CM|AB|102.9|Yaws NOS
C0043388|ICD9CM|PT|102.9|Yaws, unspecified
C0043395|ICD9CM|HT|060|Yellow fever
C0043395|ICD9CM|AB|060.9|Yellow fever NOS
C0043395|ICD9CM|PT|060.9|Yellow fever, unspecified
C0043397|ICD9CM|AB|060.0|Sylvatic yellow fever
C0043397|ICD9CM|PT|060.0|Sylvatic yellow fever
C0043398|ICD9CM|AB|060.1|Urban yellow fever
C0043398|ICD9CM|PT|060.1|Urban yellow fever
C0043541|ICD9CM|AB|117.7|Zygomycosis
C0043541|ICD9CM|PT|117.7|Zygomycosis [Phycomycosis or Mucormycosis]
C0079102|ICD9CM|HT|434.0|Cerebral thrombosis
C0079157|ICD9CM|PT|742.2|Congenital reduction deformities of brain
C0079157|ICD9CM|AB|742.2|Reduction deform, brain
C0079229|ICD9CM|PT|88.73|Diagnostic ultrasound of other sites of thorax
C0079229|ICD9CM|AB|88.73|Dx ultrasound-thorax NEC
C0079774|ICD9CM|HT|202.7|Peripheral T-cell lymphoma
C0079801|ICD9CM|AB|E008.4|Martial arts
C0079801|ICD9CM|PT|E008.4|Activities involving martial arts
C0079924|ICD9CM|HT|658.0|Oligohydramnios
C0079953|ICD9CM|PT|12.59|Other facilitation of intraocular circulation
C0079953|ICD9CM|AB|12.59|Facilit intraoc circ NEC
C0079954|ICD9CM|HT|728.7|Other fibromatoses of muscle, ligament, and fascia
C0079954|ICD9CM|PT|728.79|Other fibromatoses of muscle, ligament, and fascia
C0079954|ICD9CM|AB|728.79|Fibromatoses NEC
C0079955|ICD9CM|HT|200.8|Other named variants of lymphosarcoma and reticulosarcoma
C0079956|ICD9CM|AB|06.89|Other parathyroidectomy
C0079956|ICD9CM|PT|06.89|Other parathyroidectomy
C0079957|ICD9CM|PT|694.8|Other specified bullous dermatoses
C0079957|ICD9CM|AB|694.8|Bullous dermatoses NEC
C0079989|ICD9CM|HT|06.8|Parathyroidectomy
C0080032|ICD9CM|PT|511.81|Malignant pleural effusion
C0080032|ICD9CM|AB|511.81|Malignant pleural effusn
C0080099|ICD9CM|AB|V62.6|Refusal of treatment
C0080099|ICD9CM|PT|V62.6|Refusal of treatment for reasons of religion or conscience
C0080102|ICD9CM|PT|93.89|Rehabilitation, not elsewhere classified
C0080102|ICD9CM|AB|93.89|Rehabilitation NEC
C0080174|ICD9CM|AB|756.17|Spina bifida occulta
C0080174|ICD9CM|PT|756.17|Spina bifida occulta
C0080178|ICD9CM|HT|741|Spina bifida
C0080233|ICD9CM|PT|525.10|Acquired absence of teeth, unspecified
C0080233|ICD9CM|AB|525.10|Acq absence of teeth NOS
C0080253|ICD9CM|PT|04.6|Transposition of cranial and peripheral nerves
C0080253|ICD9CM|AB|04.6|Periph nerve transposit
C0080274|ICD9CM|HT|788.2|Retention of urine
C0080274|ICD9CM|AB|788.20|Retention urine NOS
C0080274|ICD9CM|PT|788.20|Retention of urine, unspecified
C0080276|ICD9CM|HT|580-629.99|DISEASES OF THE GENITOURINARY SYSTEM
C0085084|ICD9CM|HT|335.2|Motor neuron disease
C0085096|ICD9CM|PT|443.9|Peripheral vascular disease, unspecified
C0085096|ICD9CM|AB|443.9|Periph vascular dis NOS
C0085109|ICD9CM|HT|370.6|Corneal neovascularization
C0085109|ICD9CM|PT|370.60|Corneal neovascularization, unspecified
C0085109|ICD9CM|AB|370.60|Cornea neovasculariz NOS
C0085160|ICD9CM|AB|705.83|Hidradenitis
C0085160|ICD9CM|PT|705.83|Hidradenitis
C0085179|ICD9CM|PT|710.5|Eosinophilia myalgia syndrome
C0085179|ICD9CM|AB|710.5|Eosinophilia myalgia snd
C0085198|ICD9CM|AB|42.40|Esophagectomy NOS
C0085198|ICD9CM|HT|42.4|Excision of esophagus
C0085198|ICD9CM|PT|42.40|Esophagectomy, not otherwise specified
C0085222|ICD9CM|AB|567.31|Psoas muscle abscess
C0085222|ICD9CM|PT|567.31|Psoas muscle abscess
C0085273|ICD9CM|AB|057.0|Erythema infectiosum
C0085273|ICD9CM|PT|057.0|Erythema infectiosum (fifth disease)
C0085290|ICD9CM|AB|38.94|Venous cutdown
C0085290|ICD9CM|PT|38.94|Venous cutdown
C0085292|ICD9CM|AB|333.91|Stiff-man syndrome
C0085292|ICD9CM|PT|333.91|Stiff-man syndrome
C0085315|ICD9CM|PT|130.0|Meningoencephalitis due to toxoplasmosis
C0085315|ICD9CM|AB|130.0|Toxoplasm meningoenceph
C0085388|ICD9CM|HT|013.2|Tuberculoma of brain
C0085388|ICD9CM|AB|013.20|Tuberculoma brain-unspec
C0085388|ICD9CM|PT|013.20|Tuberculoma of brain, unspecified
C0085399|ICD9CM|HT|082.4|Ehrlichiosis
C0085399|ICD9CM|AB|082.40|Ehrlichiosis NOS
C0085399|ICD9CM|PT|082.40|Ehrlichiosis, unspecified
C0085413|ICD9CM|PT|753.13|Polycystic kidney, autosomal dominant
C0085413|ICD9CM|AB|753.13|Polycyst kid-autosom dom
C0085436|ICD9CM|AB|321.0|Cryptococcal meningitis
C0085436|ICD9CM|PT|321.0|Cryptococcal meningitis
C0085437|ICD9CM|HT|320|Bacterial meningitis
C0085437|ICD9CM|AB|320.9|Bacterial meningitis NOS
C0085437|ICD9CM|PT|320.9|Meningitis due to unspecified bacterium
C0085543|ICD9CM|HT|345.7|Epilepsia partialis continua
C0085548|ICD9CM|PT|753.14|Polycystic kidney, autosomal recessive
C0085548|ICD9CM|AB|753.14|Polycyst kid-autosom rec
C0085574|ICD9CM|HT|719.3|Palindromic rheumatism
C0085574|ICD9CM|PT|719.30|Palindromic rheumatism, site unspecified
C0085574|ICD9CM|AB|719.30|Palindrom rheum-unspec
C0085578|ICD9CM|PT|282.46|Thalassemia minor
C0085578|ICD9CM|AB|282.46|Thalassemia minor
C0085580|ICD9CM|HT|401|Essential hypertension
C0085580|ICD9CM|AB|401.9|Hypertension NOS
C0085580|ICD9CM|PT|401.9|Unspecified essential hypertension
C0085584|ICD9CM|AB|348.30|Encephalopathy NOS
C0085584|ICD9CM|PT|348.30|Encephalopathy, unspecified
C0085584|ICD9CM|HT|348.3|Encephalopathy, not elsewhere classified
C0085592|ICD9CM|AB|992.2|Heat cramps
C0085592|ICD9CM|PT|992.2|Heat cramps
C0085602|ICD9CM|AB|783.5|Polydipsia
C0085602|ICD9CM|PT|783.5|Polydipsia
C0085606|ICD9CM|AB|788.63|Urgency of urination
C0085606|ICD9CM|PT|788.63|Urgency of urination
C0085614|ICD9CM|PT|426.11|First degree atrioventricular block
C0085614|ICD9CM|AB|426.11|Atriovent block-1st degr
C0085615|ICD9CM|PT|426.4|Right bundle branch block
C0085615|ICD9CM|AB|426.4|Rt bundle branch block
C0085619|ICD9CM|AB|786.02|Orthopnea
C0085619|ICD9CM|PT|786.02|Orthopnea
C0085622|ICD9CM|AB|344.5|Monoplegia NOS
C0085622|ICD9CM|PT|344.5|Unspecified monoplegia
C0085633|ICD9CM|AB|799.24|Emotional lability
C0085633|ICD9CM|PT|799.24|Emotional lability
C0085639|ICD9CM|AB|E888.9|Fall NOS
C0085639|ICD9CM|PT|E888.9|Unspecified fall
C0085648|ICD9CM|AB|727.40|Synovial cyst NOS
C0085648|ICD9CM|PT|727.40|Synovial cyst, unspecified
C0085652|ICD9CM|AB|686.01|Pyoderma gangrenosum
C0085652|ICD9CM|PT|686.01|Pyoderma gangrenosum
C0085655|ICD9CM|AB|710.4|Polymyositis
C0085655|ICD9CM|PT|710.4|Polymyositis
C0085663|ICD9CM|PT|288.64|Plasmacytosis
C0085663|ICD9CM|AB|288.64|Plasmacytosis
C0085669|ICD9CM|HT|208.0|Leukemia of unspecified cell type, acute
C0085677|ICD9CM|AB|357.5|Alcoholic polyneuropathy
C0085677|ICD9CM|PT|357.5|Alcoholic polyneuropathy
C0085690|ICD9CM|AB|373.12|Hordeolum internum
C0085690|ICD9CM|PT|373.12|Hordeolum internum
C0085693|ICD9CM|HT|540|Acute appendicitis
C0085694|ICD9CM|AB|575.11|Chronic cholecystitis
C0085694|ICD9CM|PT|575.11|Chronic cholecystitis
C0085696|ICD9CM|AB|601.1|Chronic prostatitis
C0085696|ICD9CM|PT|601.1|Chronic prostatitis
C0085697|ICD9CM|HT|590.0|Chronic pyelonephritis
C0085700|ICD9CM|AB|733.92|Chondromalacia
C0085700|ICD9CM|PT|733.92|Chondromalacia
C0085704|ICD9CM|AB|54.11|Exploratory laparotomy
C0085704|ICD9CM|PT|54.11|Exploratory laparotomy
C0085762|ICD9CM|HT|305.0|Alcohol abuse
C0085762|ICD9CM|PT|305.00|Alcohol abuse, unspecified
C0085762|ICD9CM|AB|305.00|Alcohol abuse-unspec
C0085932|ICD9CM|HT|694|Bullous dermatoses
C0085932|ICD9CM|AB|694.9|Bullous dermatoses NOS
C0085932|ICD9CM|PT|694.9|Unspecified bullous dermatoses
C0085988|ICD9CM|HT|653.4|Fetopelvic disproportion
C0085990|ICD9CM|AB|42.11|Cervical esophagostomy
C0085990|ICD9CM|PT|42.11|Cervical esophagostomy
C0086227|ICD9CM|AB|127.4|Enterobiasis
C0086227|ICD9CM|PT|127.4|Enterobiasis
C0086438|ICD9CM|AB|279.00|Hypogammaglobulinem NOS
C0086438|ICD9CM|PT|279.00|Hypogammaglobulinemia, unspecified
C0086511|ICD9CM|AB|81.54|Total knee replacement
C0086511|ICD9CM|PT|81.54|Total knee replacement
C0086541|ICD9CM|PT|085.1|Cutaneous leishmaniasis, urban
C0086541|ICD9CM|AB|085.1|Cutan leishmanias urban
C0086543|ICD9CM|HT|366|Cataract
C0086543|ICD9CM|AB|366.9|Cataract NOS
C0086543|ICD9CM|PT|366.9|Unspecified cataract
C0086588|ICD9CM|AB|261|Nutritional marasmus
C0086588|ICD9CM|PT|261|Nutritional marasmus
C0086692|ICD9CM|HT|210-229.99|BENIGN NEOPLASMS
C0086692|ICD9CM|AB|229.9|Benign neoplasm NOS
C0086692|ICD9CM|PT|229.9|Benign neoplasm of unspecified site
C0086809|ICD9CM|PT|704.41|Pilar cyst
C0086809|ICD9CM|AB|704.41|Pilar cyst
C0086818|ICD9CM|AB|99.05|Platelet transfusion
C0086818|ICD9CM|PT|99.05|Transfusion of platelets
C0086981|ICD9CM|AB|710.2|Sicca syndrome
C0086981|ICD9CM|PT|710.2|Sicca syndrome
C0087123|ICD9CM|HT|20.0|Myringotomy
C0149504|ICD9CM|AB|349.82|Toxic encephalopathy
C0149504|ICD9CM|PT|349.82|Toxic encephalopathy
C0149505|ICD9CM|AB|375.01|Acute dacryoadenitis
C0149505|ICD9CM|PT|375.01|Acute dacryoadenitis
C0149506|ICD9CM|AB|375.42|Chronic dacryocystitis
C0149506|ICD9CM|PT|375.42|Chronic dacryocystitis
C0149507|ICD9CM|AB|376.01|Orbital cellulitis
C0149507|ICD9CM|PT|376.01|Orbital cellulitis
C0149508|ICD9CM|HT|381.6|Obstruction of Eustachian tube
C0149508|ICD9CM|PT|381.60|Obstruction of Eustachian tube, unspecified
C0149508|ICD9CM|AB|381.60|Obstr eustach tube NOS
C0149512|ICD9CM|HT|461|Acute sinusitis
C0149512|ICD9CM|AB|461.9|Acute sinusitis NOS
C0149512|ICD9CM|PT|461.9|Acute sinusitis, unspecified
C0149513|ICD9CM|HT|464.1|Acute tracheitis
C0149514|ICD9CM|AB|466.0|Acute bronchitis
C0149514|ICD9CM|PT|466.0|Acute bronchitis
C0149516|ICD9CM|HT|473|Chronic sinusitis
C0149516|ICD9CM|AB|473.9|Chronic sinusitis NOS
C0149516|ICD9CM|PT|473.9|Unspecified sinusitis (chronic)
C0149517|ICD9CM|AB|474.00|Chronic tonsillitis
C0149517|ICD9CM|PT|474.00|Chronic tonsillitis
C0149518|ICD9CM|HT|535.0|Acute gastritis
C0149519|ICD9CM|PT|571.41|Chronic persistent hepatitis
C0149519|ICD9CM|AB|571.41|Chr persistent hepatitis
C0149520|ICD9CM|AB|575.0|Acute cholecystitis
C0149520|ICD9CM|PT|575.0|Acute cholecystitis
C0149521|ICD9CM|AB|577.1|Chronic pancreatitis
C0149521|ICD9CM|PT|577.1|Chronic pancreatitis
C0149523|ICD9CM|AB|595.0|Acute cystitis
C0149523|ICD9CM|PT|595.0|Acute cystitis
C0149524|ICD9CM|AB|601.0|Acute prostatitis
C0149524|ICD9CM|PT|601.0|Acute prostatitis
C0149525|ICD9CM|AB|602.0|Calculus of prostate
C0149525|ICD9CM|PT|602.0|Calculus of prostate
C0149526|ICD9CM|AB|708.0|Allergic urticaria
C0149526|ICD9CM|PT|708.0|Allergic urticaria
C0149530|ICD9CM|AB|746.86|Congenital heart block
C0149530|ICD9CM|PT|746.86|Congenital heart block
C0149531|ICD9CM|HT|808|Fracture of pelvis
C0149532|ICD9CM|PT|935.1|Foreign body in esophagus
C0149532|ICD9CM|AB|935.1|Foreign body esophagus
C0149533|ICD9CM|AB|39.98|Hemorrhage control NOS
C0149533|ICD9CM|PT|39.98|Control of hemorrhage, not otherwise specified
C0149534|ICD9CM|AB|96.52|Irrigation of ear
C0149534|ICD9CM|PT|96.52|Irrigation of ear
C0149627|ICD9CM|PT|222.1|Benign neoplasm of penis
C0149627|ICD9CM|AB|222.1|Benign neoplasm penis
C0149649|ICD9CM|HT|445|Atheroembolism
C0149654|ICD9CM|PT|312.9|Unspecified disturbance of conduct
C0149654|ICD9CM|AB|312.9|Conduct disturbance NOS
C0149707|ICD9CM|AB|608.82|Hematospermia
C0149707|ICD9CM|PT|608.82|Hematospermia
C0149771|ICD9CM|AB|618.04|Rectocele
C0149771|ICD9CM|PT|618.04|Rectocele
C0149823|ICD9CM|PT|536.1|Acute dilatation of stomach
C0149823|ICD9CM|AB|536.1|Ac dilation of stomach
C0149825|ICD9CM|AB|474.12|Hypertrophy adenoids
C0149825|ICD9CM|PT|474.12|Hypertrophy of adenoids alone
C0149870|ICD9CM|PT|727.04|Radial styloid tenosynovitis
C0149870|ICD9CM|AB|727.04|Radial styloid tenosynov
C0149881|ICD9CM|HT|604|Orchitis and epididymitis
C0149881|ICD9CM|PT|604.90|Orchitis and epididymitis, unspecified
C0149881|ICD9CM|AB|604.90|Orchitis/epididymit NOS
C0149882|ICD9CM|AB|530.12|Acute esophagitis
C0149882|ICD9CM|PT|530.12|Acute esophagitis
C0149896|ICD9CM|AB|274.01|Acute gouty arthropathy
C0149896|ICD9CM|PT|274.01|Acute gouty arthropathy
C0149931|ICD9CM|HT|346|Migraine
C0149931|ICD9CM|HT|346.9|Migraine, unspecified
C0149966|ICD9CM|PT|098.6|Gonococcal infection of pharynx
C0149966|ICD9CM|AB|098.6|Gonococcal infec pharynx
C0149977|ICD9CM|AB|832.2|Nursemaid's elbow
C0149977|ICD9CM|PT|832.2|Nursemaid's elbow
C0149985|ICD9CM|AB|091.9|Secondary syphilis NOS
C0149985|ICD9CM|PT|091.9|Unspecified secondary syphilis
C0150042|ICD9CM|PT|788.91|Functional urinary incontinence
C0150042|ICD9CM|AB|788.91|Fnctnl urinary incontnce
C0150045|ICD9CM|AB|788.31|Urge incontinence
C0150045|ICD9CM|PT|788.31|Urge incontinence
C0150055|ICD9CM|HT|338.2|Chronic pain
C0150260|ICD9CM|PT|01.10|Intracranial pressure monitoring
C0150260|ICD9CM|AB|01.10|Intracran pressure montr
C0150411|ICD9CM|PT|89.65|Measurement of systemic arterial blood gases
C0150411|ICD9CM|AB|89.65|Arterial bld gas measure
C0150460|ICD9CM|PT|89.61|Systemic arterial pressure monitoring
C0150460|ICD9CM|AB|89.61|Arterial pressure monit
C0151295|ICD9CM|AB|354.5|Mononeuritis multiplex
C0151295|ICD9CM|PT|354.5|Mononeuritis multiplex
C0151436|ICD9CM|HT|446.2|Hypersensitivity angiitis
C0151436|ICD9CM|PT|446.20|Hypersensitivity angiitis, unspecified
C0151436|ICD9CM|AB|446.20|Hypersensit angiitis NOS
C0151482|ICD9CM|AB|281.2|Folate-deficiency anemia
C0151482|ICD9CM|PT|281.2|Folate-deficiency anemia
C0151511|ICD9CM|AB|611.4|Atrophy of breast
C0151511|ICD9CM|PT|611.4|Atrophy of breast
C0151517|ICD9CM|PT|426.0|Atrioventricular block, complete
C0151517|ICD9CM|AB|426.0|Atriovent block complete
C0151526|ICD9CM|HT|644.2|Early onset of delivery
C0151583|ICD9CM|PT|792.0|Nonspecific abnormal findings in cerebrospinal fluid
C0151583|ICD9CM|AB|792.0|Abn fnd-cerebrospinal fl
C0151601|ICD9CM|AB|372.73|Conjunctival edema
C0151601|ICD9CM|PT|372.73|Conjunctival edema
C0151620|ICD9CM|PT|437.2|Hypertensive encephalopathy
C0151620|ICD9CM|AB|437.2|Hypertens encephalopathy
C0151632|ICD9CM|PT|790.1|Elevated sedimentation rate
C0151632|ICD9CM|AB|790.1|Elevated sediment rate
C0151699|ICD9CM|PT|432.9|Unspecified intracranial hemorrhage
C0151699|ICD9CM|AB|432.9|Intracranial hemorr NOS
C0151731|ICD9CM|AB|573.4|Hepatic infarction
C0151731|ICD9CM|PT|573.4|Hepatic infarction
C0151744|ICD9CM|HT|410-414.99|ISCHEMIC HEART DISEASE
C0151766|ICD9CM|PT|794.8|Nonspecific abnormal results of function study of liver
C0151766|ICD9CM|AB|794.8|Abn liver function study
C0151779|ICD9CM|PT|172.9|Melanoma of skin, site unspecified
C0151779|ICD9CM|HT|172|Malignant melanoma of skin
C0151779|ICD9CM|AB|172.9|Malig melanoma skin NOS
C0151844|ICD9CM|AB|370.06|Perforated corneal ulcer
C0151844|ICD9CM|PT|370.06|Perforated corneal ulcer
C0151907|ICD9CM|HT|709.0|Dyschromia
C0151907|ICD9CM|AB|709.00|Dyschromia, unspecified
C0151907|ICD9CM|PT|709.00|Dyschromia, unspecified
C0151970|ICD9CM|HT|530.2|Ulcer of esophagus
C0151971|ICD9CM|AB|569.82|Ulceration of intestine
C0151971|ICD9CM|PT|569.82|Ulceration of intestine
C0152020|ICD9CM|AB|536.3|Gastroparesis
C0152020|ICD9CM|PT|536.3|Gastroparesis
C0152026|ICD9CM|AB|362.18|Retinal vasculitis
C0152026|ICD9CM|PT|362.18|Retinal vasculitis
C0152032|ICD9CM|PT|788.64|Urinary hesitancy
C0152032|ICD9CM|AB|788.64|Urinary hesitancy
C0152061|ICD9CM|PT|087.0|Relapsing fever, louse-borne
C0152061|ICD9CM|AB|087.0|Louse-borne relaps fever
C0152062|ICD9CM|AB|026.0|Spirillary fever
C0152062|ICD9CM|PT|026.0|Spirillary fever
C0152063|ICD9CM|AB|026.1|Streptobacillary fever
C0152063|ICD9CM|PT|026.1|Streptobacillary fever
C0152066|ICD9CM|AB|116.2|Lobomycosis
C0152066|ICD9CM|PT|116.2|Lobomycosis
C0152067|ICD9CM|AB|111.1|Tinea nigra
C0152067|ICD9CM|PT|111.1|Tinea nigra
C0152068|ICD9CM|PT|122.4|Echinococcus granulosus infection, unspecified
C0152068|ICD9CM|AB|122.4|Echinococc granul NOS
C0152069|ICD9CM|PT|122.7|Echinococcus multilocularis infection, unspecified
C0152069|ICD9CM|AB|122.7|Echinococc multiloc NOS
C0152070|ICD9CM|AB|125.1|Malayan filariasis
C0152070|ICD9CM|PT|125.1|Malayan filariasis
C0152071|ICD9CM|AB|121.6|Heterophyiasis
C0152071|ICD9CM|PT|121.6|Heterophyiasis
C0152072|ICD9CM|AB|084.3|Ovale malaria
C0152072|ICD9CM|PT|084.3|Ovale malaria
C0152073|ICD9CM|PT|123.2|Taenia saginata infection
C0152073|ICD9CM|AB|123.2|Taenia saginata infect
C0152074|ICD9CM|PT|085.3|Cutaneous leishmaniasis, Ethiopian
C0152074|ICD9CM|AB|085.3|Cutan leishmanias ethiop
C0152077|ICD9CM|AB|246.1|Dyshormonogenic goiter
C0152077|ICD9CM|PT|246.1|Dyshormonogenic goiter
C0152078|ICD9CM|PT|625.5|Pelvic congestion syndrome
C0152078|ICD9CM|AB|625.5|Pelvic congestion synd
C0152079|ICD9CM|PT|620.6|Broad ligament laceration syndrome
C0152079|ICD9CM|AB|620.6|Broad ligament lacer syn
C0152083|ICD9CM|HT|716.4|Transient arthropathy
C0152083|ICD9CM|PT|716.40|Transient arthropathy, site unspecified
C0152083|ICD9CM|AB|716.40|Trans arthropathy-unspec
C0152084|ICD9CM|PT|714.4|Chronic postrheumatic arthropathy
C0152084|ICD9CM|AB|714.4|Chr postrheum arthritis
C0152085|ICD9CM|PT|711.30|Postdysenteric arthropathy, site unspecified
C0152085|ICD9CM|HT|711.3|Postdysenteric arthropathy
C0152085|ICD9CM|AB|711.30|Dysenter arthrit-unspec
C0152086|ICD9CM|HT|716.1|Traumatic arthropathy
C0152086|ICD9CM|PT|716.10|Traumatic arthropathy, site unspecified
C0152086|ICD9CM|AB|716.10|Traum arthropathy-unspec
C0152087|ICD9CM|HT|712|Crystal arthropathies
C0152087|ICD9CM|HT|712.9|Unspecified crystal arthropathy
C0152087|ICD9CM|PT|712.90|Unspecified crystal arthropathy, site unspecified
C0152087|ICD9CM|AB|712.90|Cryst arthrop NOS-unspec
C0152088|ICD9CM|AB|721.7|Traumatic spondylopathy
C0152088|ICD9CM|PT|721.7|Traumatic spondylopathy
C0152089|ICD9CM|PT|722.80|Postlaminectomy syndrome, unspecified region
C0152089|ICD9CM|HT|722.8|Postlaminectomy syndrome
C0152089|ICD9CM|AB|722.80|Postlaminectomy synd NOS
C0152090|ICD9CM|AB|720.1|Spinal enthesopathy
C0152090|ICD9CM|PT|720.1|Spinal enthesopathy
C0152091|ICD9CM|HT|732|Osteochondropathies
C0152091|ICD9CM|AB|732.9|Osteochondropathy NOS
C0152091|ICD9CM|PT|732.9|Unspecified osteochondropathy
C0152091|ICD9CM|PT|733.90|Disorder of bone and cartilage, unspecified
C0152091|ICD9CM|AB|733.90|Bone & cartilage dis NOS
C0152092|ICD9CM|PT|694.2|Juvenile dermatitis herpetiformis
C0152092|ICD9CM|AB|694.2|Juven dermat herpetiform
C0152093|ICD9CM|AB|728.5|Hypermobility syndrome
C0152093|ICD9CM|PT|728.5|Hypermobility syndrome
C0152094|ICD9CM|AB|279.13|Nezelof's syndrome
C0152094|ICD9CM|PT|279.13|Nezelof's syndrome
C0152095|ICD9CM|AB|758.1|Patau's syndrome
C0152095|ICD9CM|PT|758.1|Patau's syndrome
C0152096|ICD9CM|AB|758.2|Edwards' syndrome
C0152096|ICD9CM|PT|758.2|Edwards' syndrome
C0152097|ICD9CM|AB|519.4|Disorders of diaphragm
C0152097|ICD9CM|PT|519.4|Disorders of diaphragm
C0152099|ICD9CM|PT|576.0|Postcholecystectomy syndrome
C0152099|ICD9CM|AB|576.0|Postcholecystectomy synd
C0152101|ICD9CM|PT|746.7|Hypoplastic left heart syndrome
C0152101|ICD9CM|AB|746.7|Hypoplas left heart synd
C0152102|ICD9CM|PT|416.1|Kyphoscoliotic heart disease
C0152102|ICD9CM|AB|416.1|Kyphoscoliotic heart dis
C0152105|ICD9CM|HT|402|Hypertensive heart disease
C0152105|ICD9CM|HT|402.9|Unspecified hypertensive heart disease
C0152107|ICD9CM|PT|411.0|Postmyocardial infarction syndrome
C0152107|ICD9CM|AB|411.0|Post MI syndrome
C0152108|ICD9CM|AB|495.3|Suberosis
C0152108|ICD9CM|PT|495.3|Suberosis
C0152109|ICD9CM|PT|335.11|Kugelberg-Welander disease
C0152109|ICD9CM|AB|335.11|Kugelberg-welander dis
C0152110|ICD9CM|AB|355.1|Meralgia paresthetica
C0152110|ICD9CM|PT|355.1|Meralgia paresthetica
C0152112|ICD9CM|PT|377.04|Foster-Kennedy syndrome
C0152112|ICD9CM|AB|377.04|Foster-kennedy syndrome
C0152113|ICD9CM|HT|392|Rheumatic chorea
C0152115|ICD9CM|AB|333.82|Orofacial dyskinesia
C0152115|ICD9CM|PT|333.82|Orofacial dyskinesia
C0152116|ICD9CM|AB|333.83|Spasmodic torticollis
C0152116|ICD9CM|PT|333.83|Spasmodic torticollis
C0152124|ICD9CM|AB|298.2|Reactive confusion
C0152124|ICD9CM|PT|298.2|Reactive confusion
C0152125|ICD9CM|AB|298.3|Acute paranoid reaction
C0152125|ICD9CM|PT|298.3|Acute paranoid reaction
C0152126|ICD9CM|PT|298.4|Psychogenic paranoid psychosis
C0152126|ICD9CM|AB|298.4|Psychogen paranoid psych
C0152128|ICD9CM|AB|292.0|Drug withdrawal
C0152128|ICD9CM|PT|292.0|Drug withdrawal
C0152129|ICD9CM|PT|292.2|Pathological drug intoxication
C0152129|ICD9CM|AB|292.2|Pathologic drug intox
C0152131|ICD9CM|AB|363.31|Solar retinopathy
C0152131|ICD9CM|PT|363.31|Solar retinopathy
C0152132|ICD9CM|AB|362.11|Hypertensive retinopathy
C0152132|ICD9CM|PT|362.11|Hypertensive retinopathy
C0152134|ICD9CM|PT|378.86|Internuclear ophthalmoplegia
C0152134|ICD9CM|AB|378.86|Internucl ophthalmopleg
C0152135|ICD9CM|PT|376.22|Exophthalmic ophthalmoplegia
C0152135|ICD9CM|AB|376.22|Exophthalm ophthalmopleg
C0152136|ICD9CM|AB|365.12|Low tension glaucoma
C0152136|ICD9CM|PT|365.12|Low tension open-angle glaucoma
C0152137|ICD9CM|AB|365.51|Phacolytic glaucoma
C0152137|ICD9CM|PT|365.51|Phacolytic glaucoma
C0152138|ICD9CM|PT|364.22|Glaucomatocyclitic crises
C0152138|ICD9CM|AB|364.22|Glaucomatocyclit crises
C0152144|ICD9CM|PT|992.4|Heat exhaustion due to salt depletion
C0152144|ICD9CM|AB|992.4|Heat exhaust-salt deple
C0152145|ICD9CM|AB|992.6|Heat fatigue, transient
C0152145|ICD9CM|PT|992.6|Heat fatigue, transient
C0152149|ICD9CM|AB|625.2|Mittelschmerz
C0152149|ICD9CM|PT|625.2|Mittelschmerz
C0152150|ICD9CM|HT|651.0|Twin pregnancy
C0152151|ICD9CM|HT|651.1|Triplet pregnancy
C0152152|ICD9CM|HT|651.2|Quadruplet pregnancy
C0152154|ICD9CM|HT|662.1|Prolonged labor, unspecified
C0152154|ICD9CM|HT|662|Long labor
C0152156|ICD9CM|HT|660|Obstructed labor
C0152156|ICD9CM|HT|660.9|Unspecified obstructed labor
C0152158|ICD9CM|HT|676.4|Failure of lactation
C0152158|ICD9CM|PT|676.40|Failure of lactation, unspecified as to episode of care or not applicable
C0152158|ICD9CM|AB|676.40|Lactation fail-unspec
C0152159|ICD9CM|HT|661.0|Primary uterine inertia
C0152163|ICD9CM|AB|537.81|Pylorospasm
C0152163|ICD9CM|PT|537.81|Pylorospasm
C0152165|ICD9CM|AB|536.2|Persistent vomiting
C0152165|ICD9CM|PT|536.2|Persistent vomiting
C0152166|ICD9CM|AB|579.4|Pancreatic steatorrhea
C0152166|ICD9CM|PT|579.4|Pancreatic steatorrhea
C0152167|ICD9CM|AB|564.6|Anal spasm
C0152167|ICD9CM|PT|564.6|Anal spasm
C0152168|ICD9CM|PT|576.5|Spasm of sphincter of Oddi
C0152168|ICD9CM|AB|576.5|Spasm sphincter of oddi
C0152169|ICD9CM|AB|788.0|Renal colic
C0152169|ICD9CM|PT|788.0|Renal colic
C0152171|ICD9CM|PT|416.0|Primary pulmonary hypertension
C0152171|ICD9CM|AB|416.0|Prim pulm hypertension
C0152172|ICD9CM|AB|413.0|Angina decubitus
C0152172|ICD9CM|PT|413.0|Angina decubitus
C0152173|ICD9CM|AB|427.42|Ventricular flutter
C0152173|ICD9CM|PT|427.42|Ventricular flutter
C0152174|ICD9CM|AB|307.80|Psychogenic pain NOS
C0152174|ICD9CM|PT|307.80|Psychogenic pain, site unspecified
C0152177|ICD9CM|HT|350|Trigeminal nerve disorders
C0152177|ICD9CM|PT|350.9|Trigeminal nerve disorder, unspecified
C0152177|ICD9CM|AB|350.9|Trigeminal nerve dis NOS
C0152179|ICD9CM|PT|352.3|Disorders of pneumogastric [10th] nerve
C0152179|ICD9CM|AB|352.3|Pneumogastric nerve dis
C0152180|ICD9CM|AB|352.4|Accessory nerve disorder
C0152180|ICD9CM|PT|352.4|Disorders of accessory [11th] nerve
C0152181|ICD9CM|PT|352.5|Disorders of hypoglossal [12th] nerve
C0152181|ICD9CM|AB|352.5|Hypoglossal nerve dis
C0152183|ICD9CM|PT|301.3|Explosive personality disorder
C0152183|ICD9CM|AB|301.3|Explosive personality
C0152186|ICD9CM|AB|302.1|Zoophilia
C0152186|ICD9CM|PT|302.1|Zoophilia
C0152187|ICD9CM|HT|368.0|Amblyopia ex anopsia
C0152189|ICD9CM|AB|368.02|Deprivation amblyopia
C0152189|ICD9CM|PT|368.02|Deprivation amblyopia
C0152190|ICD9CM|AB|368.03|Refractive amblyopia
C0152190|ICD9CM|PT|368.03|Refractive amblyopia
C0152191|ICD9CM|AB|368.41|Central scotoma
C0152191|ICD9CM|PT|368.41|Scotoma involving central area
C0152192|ICD9CM|PT|368.42|Scotoma of blind spot area
C0152192|ICD9CM|AB|368.42|Scotoma of blind spot
C0152193|ICD9CM|AB|367.21|Regular astigmatism
C0152193|ICD9CM|PT|367.21|Regular astigmatism
C0152194|ICD9CM|AB|367.22|Irregular astigmatism
C0152194|ICD9CM|PT|367.22|Irregular astigmatism
C0152196|ICD9CM|AB|367.53|Spasm of accommodation
C0152196|ICD9CM|PT|367.53|Spasm of accommodation
C0152197|ICD9CM|PT|367.52|Total or complete internal ophthalmoplegia
C0152197|ICD9CM|AB|367.52|Tot intern ophthalmopleg
C0152198|ICD9CM|HT|367.5|Disorders of accommodation
C0152200|ICD9CM|AB|368.54|Achromatopsia
C0152200|ICD9CM|PT|368.54|Achromatopsia
C0152202|ICD9CM|AB|368.62|Acquired night blindness
C0152202|ICD9CM|PT|368.62|Acquired night blindness
C0152204|ICD9CM|AB|378.01|Monocular esotropia
C0152204|ICD9CM|PT|378.01|Monocular esotropia
C0152205|ICD9CM|AB|378.05|Alternating esotropia
C0152205|ICD9CM|PT|378.05|Alternating esotropia
C0152206|ICD9CM|AB|378.11|Monocular exotropia
C0152206|ICD9CM|PT|378.11|Monocular exotropia
C0152207|ICD9CM|AB|378.15|Alternating exotropia
C0152207|ICD9CM|PT|378.15|Alternating exotropia
C0152208|ICD9CM|AB|378.32|Hypotropia
C0152208|ICD9CM|PT|378.32|Hypotropia
C0152209|ICD9CM|AB|378.33|Cyclotropia
C0152209|ICD9CM|PT|378.33|Cyclotropia
C0152210|ICD9CM|HT|378.2|Intermittent heterotropia
C0152210|ICD9CM|PT|378.20|Intermittent heterotropia, unspecified
C0152210|ICD9CM|AB|378.20|Intermit heterotrop NOS
C0152211|ICD9CM|PT|378.21|Intermittent esotropia, monocular
C0152211|ICD9CM|AB|378.21|Intermit monoc esotropia
C0152212|ICD9CM|PT|378.22|Intermittent esotropia, alternating
C0152212|ICD9CM|AB|378.22|Intermit altrn esotropia
C0152213|ICD9CM|PT|378.23|Intermittent exotropia, monocular
C0152213|ICD9CM|AB|378.23|Intermit monoc exotropia
C0152214|ICD9CM|PT|378.24|Intermittent exotropia, alternating
C0152214|ICD9CM|AB|378.24|Intermit altrn exotropia
C0152216|ICD9CM|AB|378.41|Esophoria
C0152216|ICD9CM|PT|378.41|Esophoria
C0152217|ICD9CM|AB|378.42|Exophoria
C0152217|ICD9CM|PT|378.42|Exophoria
C0152218|ICD9CM|AB|378.43|Vertical heterophoria
C0152218|ICD9CM|PT|378.43|Vertical heterophoria
C0152219|ICD9CM|AB|378.44|Cyclophoria
C0152219|ICD9CM|PT|378.44|Cyclophoria
C0152220|ICD9CM|AB|378.45|Alternating hyperphoria
C0152220|ICD9CM|PT|378.45|Alternating hyperphoria
C0152221|ICD9CM|HT|378.5|Paralytic strabismus
C0152221|ICD9CM|AB|378.50|Paralytic strabismus NOS
C0152221|ICD9CM|PT|378.50|Paralytic strabismus, unspecified
C0152223|ICD9CM|HT|378.6|Mechanical strabismus
C0152223|ICD9CM|PT|378.60|Mechanical strabismus, unspecified
C0152223|ICD9CM|AB|378.60|Mechanical strabism NOS
C0152225|ICD9CM|AB|379.52|Latent nystagmus
C0152225|ICD9CM|PT|379.52|Latent nystagmus
C0152226|ICD9CM|HT|374.2|Lagophthalmos
C0152226|ICD9CM|AB|374.20|Lagophthalmos NOS
C0152226|ICD9CM|PT|374.20|Lagophthalmos, unspecified
C0152227|ICD9CM|HT|375.2|Epiphora
C0152227|ICD9CM|AB|375.20|Epiphora NOS
C0152227|ICD9CM|PT|375.20|Epiphora, unspecified as to cause
C0152228|ICD9CM|AB|388.41|Diplacusis
C0152228|ICD9CM|PT|388.41|Diplacusis
C0152229|ICD9CM|AB|798.9|Unattended death
C0152229|ICD9CM|PT|798.9|Unattended death
C0152230|ICD9CM|AB|708.5|Cholinergic urticaria
C0152230|ICD9CM|PT|708.5|Cholinergic urticaria
C0152234|ICD9CM|AB|740.2|Iniencephaly
C0152234|ICD9CM|PT|740.2|Iniencephaly
C0152235|ICD9CM|PT|754.40|Genu recurvatum
C0152235|ICD9CM|AB|754.40|Cong genu recurvatum
C0152236|ICD9CM|AB|754.60|Talipes valgus
C0152236|ICD9CM|PT|754.60|Talipes valgus
C0152238|ICD9CM|AB|745.7|Cor biloculare
C0152238|ICD9CM|PT|745.7|Cor biloculare
C0152239|ICD9CM|PT|748.61|Congenital bronchiectasis
C0152239|ICD9CM|AB|748.61|Congen bronchiectasis
C0152240|ICD9CM|AB|752.35|Septate uterus
C0152240|ICD9CM|PT|752.35|Septate uterus
C0152240|ICD9CM|AB|752.2|Doubling of uterus
C0152240|ICD9CM|PT|752.2|Doubling of uterus
C0152242|ICD9CM|AB|492.0|Emphysematous bleb
C0152242|ICD9CM|PT|492.0|Emphysematous bleb
C0152243|ICD9CM|AB|611.5|Galactocele
C0152243|ICD9CM|PT|611.5|Galactocele
C0152244|ICD9CM|AB|733.22|Aneurysmal bone cyst
C0152244|ICD9CM|PT|733.22|Aneurysmal bone cyst
C0152245|ICD9CM|AB|788.8|Extravasation of urine
C0152245|ICD9CM|PT|788.8|Extravasation of urine
C0152246|ICD9CM|AB|364.76|Iridodialysis
C0152246|ICD9CM|PT|364.76|Iridodialysis
C0152247|ICD9CM|AB|599.3|Urethral caruncle
C0152247|ICD9CM|PT|599.3|Urethral caruncle
C0152249|ICD9CM|AB|706.0|Acne varioliformis
C0152249|ICD9CM|PT|706.0|Acne varioliformis
C0152250|ICD9CM|AB|453.1|Thrombophlebitis migrans
C0152250|ICD9CM|PT|453.1|Thrombophlebitis migrans
C0152251|ICD9CM|AB|695.0|Toxic erythema
C0152251|ICD9CM|PT|695.0|Toxic erythema
C0152252|ICD9CM|AB|364.72|Anterior synechiae
C0152252|ICD9CM|PT|364.72|Anterior synechiae of iris
C0152253|ICD9CM|AB|364.71|Posterior synechiae
C0152253|ICD9CM|PT|364.71|Posterior synechiae of iris
C0152255|ICD9CM|AB|372.51|Pinguecula
C0152255|ICD9CM|PT|372.51|Pinguecula
C0152256|ICD9CM|AB|733.03|Disuse osteoporosis
C0152256|ICD9CM|PT|733.03|Disuse osteoporosis
C0152258|ICD9CM|AB|366.18|Hypermature cataract
C0152258|ICD9CM|PT|366.18|Hypermature cataract
C0152259|ICD9CM|HT|366.3|Cataract secondary to ocular disorders
C0152260|ICD9CM|AB|366.51|Soemmering's ring
C0152260|ICD9CM|PT|366.51|Soemmering's ring
C0152262|ICD9CM|AB|595.81|Cystitis cystica
C0152262|ICD9CM|PT|595.81|Cystitis cystica
C0152263|ICD9CM|AB|733.5|Osteitis condensans
C0152263|ICD9CM|PT|733.5|Osteitis condensans
C0152264|ICD9CM|AB|289.6|Familial polycythemia
C0152264|ICD9CM|PT|289.6|Familial polycythemia
C0152266|ICD9CM|HT|201.6|Hodgkin's disease, mixed cellularity
C0152267|ICD9CM|HT|201.7|Hodgkin's disease, lymphocytic depletion
C0152268|ICD9CM|HT|201.5|Hodgkin's disease, nodular sclerosis
C0152271|ICD9CM|HT|204.2|Lymphoid leukemia, subacute
C0152272|ICD9CM|HT|207.1|Chronic erythremia
C0152275|ICD9CM|HT|206.2|Monocytic leukemia, subacute
C0152413|ICD9CM|PT|480.1|Pneumonia due to respiratory syncytial virus
C0152413|ICD9CM|AB|480.1|Resp syncyt viral pneum
C0152415|ICD9CM|AB|750.0|Tongue tie
C0152415|ICD9CM|PT|750.0|Tongue tie
C0152417|ICD9CM|PT|746.3|Congenital stenosis of aortic valve
C0152417|ICD9CM|AB|746.3|Cong aorta valv stenosis
C0152419|ICD9CM|AB|747.11|Interrupt of aortic arch
C0152419|ICD9CM|PT|747.11|Interruption of aortic arch
C0152421|ICD9CM|AB|744.22|Macrotia
C0152421|ICD9CM|PT|744.22|Macrotia
C0152422|ICD9CM|AB|743.35|Congenital aphakia
C0152422|ICD9CM|PT|743.35|Congenital aphakia
C0152423|ICD9CM|AB|744.23|Microtia
C0152423|ICD9CM|PT|744.23|Microtia
C0152424|ICD9CM|AB|745.3|Common ventricle
C0152424|ICD9CM|PT|745.3|Common ventricle
C0152426|ICD9CM|AB|740.1|Craniorachischisis
C0152426|ICD9CM|PT|740.1|Craniorachischisis
C0152427|ICD9CM|HT|755.0|Polydactyly
C0152427|ICD9CM|AB|755.00|Polydactyly NOS
C0152427|ICD9CM|PT|755.00|Polydactyly, unspecified digits
C0152429|ICD9CM|AB|750.22|Accessory salivary gland
C0152429|ICD9CM|PT|750.22|Accessory salivary gland
C0152430|ICD9CM|AB|755.61|Congenital coxa valga
C0152430|ICD9CM|PT|755.61|Coxa valga, congenital
C0152431|ICD9CM|AB|755.62|Congenital coxa vara
C0152431|ICD9CM|PT|755.62|Coxa vara, congenital
C0152432|ICD9CM|PT|754.44|Congenital bowing of unspecified long bones of leg
C0152432|ICD9CM|AB|754.44|Cong bowing leg NOS
C0152436|ICD9CM|AB|752.42|Imperforate hymen
C0152436|ICD9CM|PT|752.42|Imperforate hymen
C0152437|ICD9CM|HT|674.4|Placental polyp
C0152438|ICD9CM|PT|755.52|Congenital elevation of scapula
C0152438|ICD9CM|AB|755.52|Cong elevation-scapula
C0152439|ICD9CM|AB|361.10|Retinoschisis NOS
C0152439|ICD9CM|PT|361.10|Retinoschisis, unspecified
C0152440|ICD9CM|AB|371.73|Corneal staphyloma
C0152440|ICD9CM|PT|371.73|Corneal staphyloma
C0152441|ICD9CM|AB|755.54|Madelung's deformity
C0152441|ICD9CM|PT|755.54|Madelung's deformity
C0152442|ICD9CM|AB|610.4|Mammary duct ectasia
C0152442|ICD9CM|PT|610.4|Mammary duct ectasia
C0152443|ICD9CM|AB|599.2|Urethral diverticulum
C0152443|ICD9CM|PT|599.2|Urethral diverticulum
C0152444|ICD9CM|AB|742.53|Hydromyelia
C0152444|ICD9CM|PT|742.53|Hydromyelia
C0152445|ICD9CM|AB|575.3|Hydrops of gallbladder
C0152445|ICD9CM|PT|575.3|Hydrops of gallbladder
C0152447|ICD9CM|AB|788.7|Urethral discharge
C0152447|ICD9CM|PT|788.7|Urethral discharge
C0152448|ICD9CM|AB|681.01|Felon
C0152448|ICD9CM|PT|681.01|Felon
C0152450|ICD9CM|AB|517.1|Rheumatic pneumonia
C0152450|ICD9CM|PT|517.1|Rheumatic pneumonia
C0152451|ICD9CM|HT|582|Chronic glomerulonephritis
C0152452|ICD9CM|AB|423.1|Adhesive pericarditis
C0152452|ICD9CM|PT|423.1|Adhesive pericarditis
C0152453|ICD9CM|AB|611.2|Fissure of nipple
C0152453|ICD9CM|PT|611.2|Fissure of nipple
C0152454|ICD9CM|AB|372.63|Symblepharon
C0152454|ICD9CM|PT|372.63|Symblepharon
C0152455|ICD9CM|AB|371.45|Keratomalacia NOS
C0152455|ICD9CM|PT|371.45|Keratomalacia NOS
C0152456|ICD9CM|PT|575.6|Cholesterolosis of gallbladder
C0152456|ICD9CM|AB|575.6|Gb cholesterolosis
C0152457|ICD9CM|PT|371.14|Kayser-Fleischer ring
C0152457|ICD9CM|AB|371.14|Kayser-fleischer ring
C0152458|ICD9CM|AB|360.44|Leucocoria
C0152458|ICD9CM|PT|360.44|Leucocoria
C0152459|ICD9CM|AB|701.3|Striae atrophicae
C0152459|ICD9CM|PT|701.3|Striae atrophicae
C0152460|ICD9CM|PT|607.81|Balanitis xerotica obliterans
C0152460|ICD9CM|AB|607.81|Balanitis xerotica oblit
C0152461|ICD9CM|HT|42.0|Esophagotomy
C0152462|ICD9CM|HT|16.0|Orbitotomy
C0152463|ICD9CM|HT|34.5|Pleurectomy
C0152485|ICD9CM|HT|003|Other salmonella infections
C0152486|ICD9CM|AB|003.1|Salmonella septicemia
C0152486|ICD9CM|PT|003.1|Salmonella septicemia
C0152487|ICD9CM|HT|003.2|Localized salmonella infections
C0152487|ICD9CM|PT|003.20|Localized salmonella infection, unspecified
C0152487|ICD9CM|AB|003.20|Local salmonella inf NOS
C0152488|ICD9CM|AB|003.21|Salmonella meningitis
C0152488|ICD9CM|PT|003.21|Salmonella meningitis
C0152489|ICD9CM|AB|003.22|Salmonella pneumonia
C0152489|ICD9CM|PT|003.22|Salmonella pneumonia
C0152490|ICD9CM|AB|003.23|Salmonella arthritis
C0152490|ICD9CM|PT|003.23|Salmonella arthritis
C0152491|ICD9CM|AB|003.24|Salmonella osteomyelitis
C0152491|ICD9CM|PT|003.24|Salmonella osteomyelitis
C0152492|ICD9CM|PT|003.29|Other localized salmonella infections
C0152492|ICD9CM|AB|003.29|Local salmonella inf NEC
C0152493|ICD9CM|PT|004.8|Other specified shigella infections
C0152493|ICD9CM|AB|004.8|Shigella infection NEC
C0152496|ICD9CM|PT|005.3|Food poisoning due to other Clostridia
C0152496|ICD9CM|AB|005.3|Food pois: clostrid NEC
C0152497|ICD9CM|PT|005.4|Food poisoning due to Vibrio parahaemolyticus
C0152497|ICD9CM|AB|005.4|Food pois: v. parahaem
C0152498|ICD9CM|HT|005.8|Other bacterial food poisoning
C0152498|ICD9CM|PT|005.89|Other bacterial food poisoning
C0152498|ICD9CM|HT|005|Other food poisoning (bacterial)
C0152498|ICD9CM|AB|005.89|Bact food poisoning NEC
C0152500|ICD9CM|PT|006.1|Chronic intestinal amebiasis without mention of abscess
C0152500|ICD9CM|AB|006.1|Chr amebiasis w/o absces
C0152501|ICD9CM|PT|006.2|Amebic nondysenteric colitis
C0152501|ICD9CM|AB|006.2|Amebic nondysent colitis
C0152502|ICD9CM|AB|006.4|Amebic lung abscess
C0152502|ICD9CM|PT|006.4|Amebic lung abscess
C0152503|ICD9CM|AB|006.5|Amebic brain abscess
C0152503|ICD9CM|PT|006.5|Amebic brain abscess
C0152505|ICD9CM|PT|006.8|Amebic infection of other sites
C0152505|ICD9CM|AB|006.8|Amebic infection NEC
C0152506|ICD9CM|HT|007|Other protozoal intestinal diseases
C0152507|ICD9CM|PT|007.8|Other specified protozoal intestinal diseases
C0152507|ICD9CM|AB|007.8|Protozoal intest dis NEC
C0152511|ICD9CM|PT|008.1|Intestinal infection due to arizona group of paracolon bacilli
C0152511|ICD9CM|AB|008.1|Arizona enteritis
C0152513|ICD9CM|PT|008.3|Intestinal infection due to proteus (mirabilis) (morganii)
C0152513|ICD9CM|AB|008.3|Proteus enteritis
C0152515|ICD9CM|PT|008.42|Intestinal infection due to pseudomonas
C0152515|ICD9CM|AB|008.42|Pseudomonas enteritis
C0152516|ICD9CM|AB|008.5|Bacterial enteritis NOS
C0152516|ICD9CM|PT|008.5|Bacterial enteritis, unspecified
C0152517|ICD9CM|HT|008.6|Enteritis due to specified virus
C0152518|ICD9CM|HT|008|Intestinal infections due to other organisms
C0152519|ICD9CM|HT|009|Ill-defined intestinal infections
C0152522|ICD9CM|PT|009.3|Diarrhea of presumed infectious origin
C0152522|ICD9CM|AB|009.3|Diarrhea of infect orig
C0152531|ICD9CM|HT|010.1|Tuberculous pleurisy in primary progressive tuberculosis
C0152532|ICD9CM|PT|010.11|Tuberculous pleurisy in primary progressive tuberculosis, bacteriological or histological examination not done
C0152532|ICD9CM|AB|010.11|Prim TB pleurisy-no exam
C0152533|ICD9CM|PT|010.12|Tuberculous pleurisy in primary progressive tuberculosis, bacteriological or histological examination unknown (at present)
C0152533|ICD9CM|AB|010.12|Prim TB pleur-exam unkn
C0152534|ICD9CM|PT|010.13|Tuberculous pleurisy in primary progressive tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152534|ICD9CM|AB|010.13|Prim TB pleuris-micro dx
C0152535|ICD9CM|PT|010.14|Tuberculous pleurisy in primary progressive tuberculosis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152535|ICD9CM|AB|010.14|Prim TB pleurisy-cult dx
C0152536|ICD9CM|PT|010.15|Tuberculous pleurisy in primary progressive tuberculosis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152536|ICD9CM|AB|010.15|Prim TB pleuris-histo dx
C0152537|ICD9CM|PT|010.16|Tuberculous pleurisy in primary progressive tuberculosis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152537|ICD9CM|AB|010.16|Prim TB pleuris-oth test
C0152538|ICD9CM|HT|010.8|Other primary progressive tuberculosis
C0152539|ICD9CM|PT|010.81|Other primary progressive tuberculosis, bacteriological or histological examination not done
C0152539|ICD9CM|AB|010.81|Prim prog TB NEC-no exam
C0152540|ICD9CM|PT|010.82|Other primary progressive tuberculosis, bacteriological or histological examination unknown (at present)
C0152540|ICD9CM|AB|010.82|Prim pr TB NEC-exam unkn
C0152541|ICD9CM|PT|010.83|Other primary progressive tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152541|ICD9CM|AB|010.83|Prim prg TB NEC-micro dx
C0152542|ICD9CM|PT|010.84|Other primary progressive tuberculosis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152542|ICD9CM|AB|010.84|Prim prog TB NEC-cult dx
C0152543|ICD9CM|PT|010.85|Other primary progressive tuberculosis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152543|ICD9CM|AB|010.85|Prim prg TB NEC-histo dx
C0152544|ICD9CM|PT|010.86|Other primary progressive tuberculosis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152544|ICD9CM|AB|010.86|Prim prg TB NEC-oth test
C0152545|ICD9CM|HT|010|Primary tuberculous infection
C0152545|ICD9CM|HT|010.0|Primary tuberculous infection
C0152546|ICD9CM|PT|010.91|Primary tuberculous infection, unspecified, bacteriological or histological examination not done
C0152546|ICD9CM|AB|010.91|Primary TB NOS-no exam
C0152547|ICD9CM|PT|010.92|Primary tuberculous infection, unspecified, bacteriological or histological examination unknown (at present)
C0152547|ICD9CM|AB|010.92|Primary TB NOS-exam unkn
C0152548|ICD9CM|PT|010.93|Primary tuberculous infection, unspecified, tubercle bacilli found (in sputum) by microscopy
C0152548|ICD9CM|AB|010.93|Primary TB NOS-micro dx
C0152549|ICD9CM|PT|010.94|Primary tuberculous infection, unspecified, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152549|ICD9CM|AB|010.94|Primary TB NOS-cult dx
C0152550|ICD9CM|PT|010.95|Primary tuberculous infection, unspecified, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152550|ICD9CM|AB|010.95|Primary TB NOS-histo dx
C0152551|ICD9CM|PT|010.96|Primary tuberculous infection, unspecified, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152551|ICD9CM|AB|010.96|Primary TB NOS-oth test
C0152552|ICD9CM|HT|011.0|Tuberculosis of lung, infiltrative
C0152552|ICD9CM|AB|011.00|TB lung infiltr-unspec
C0152552|ICD9CM|PT|011.00|Tuberculosis of lung, infiltrative, unspecified
C0152553|ICD9CM|PT|011.01|Tuberculosis of lung, infiltrative, bacteriological or histological examination not done
C0152553|ICD9CM|AB|011.01|TB lung infiltr-no exam
C0152554|ICD9CM|PT|011.02|Tuberculosis of lung, infiltrative, bacteriological or histological examination unknown (at present)
C0152554|ICD9CM|AB|011.02|TB lung infiltr-exm unkn
C0152555|ICD9CM|PT|011.03|Tuberculosis of lung, infiltrative, tubercle bacilli found (in sputum) by microscopy
C0152555|ICD9CM|AB|011.03|TB lung infiltr-micro dx
C0152556|ICD9CM|PT|011.04|Tuberculosis of lung, infiltrative, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152556|ICD9CM|AB|011.04|TB lung infiltr-cult dx
C0152557|ICD9CM|PT|011.05|Tuberculosis of lung, infiltrative, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152557|ICD9CM|AB|011.05|TB lung infiltr-histo dx
C0152558|ICD9CM|PT|011.06|Tuberculosis of lung, infiltrative, tubercle bacilli not found bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152558|ICD9CM|AB|011.06|TB lung infiltr-oth test
C0152559|ICD9CM|HT|011.1|Tuberculosis of lung, nodular
C0152559|ICD9CM|AB|011.10|TB lung nodular-unspec
C0152559|ICD9CM|PT|011.10|Tuberculosis of lung, nodular, unspecified
C0152560|ICD9CM|PT|011.11|Tuberculosis of lung, nodular, bacteriological or histological examination not done
C0152560|ICD9CM|AB|011.11|TB lung nodular-no exam
C0152561|ICD9CM|PT|011.12|Tuberculosis of lung, nodular, bacteriological or histological examination unknown (at present)
C0152561|ICD9CM|AB|011.12|TB lung nodul-exam unkn
C0152562|ICD9CM|PT|011.13|Tuberculosis of lung, nodular, tubercle bacilli found (in sputum) by microscopy
C0152562|ICD9CM|AB|011.13|TB lung nodular-micro dx
C0152563|ICD9CM|PT|011.14|Tuberculosis of lung, nodular, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152563|ICD9CM|AB|011.14|TB lung nodular-cult dx
C0152564|ICD9CM|PT|011.15|Tuberculosis of lung, nodular, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152564|ICD9CM|AB|011.15|TB lung nodular-histo dx
C0152565|ICD9CM|PT|011.16|Tuberculosis of lung, nodular, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152565|ICD9CM|AB|011.16|TB lung nodular-oth test
C0152566|ICD9CM|HT|011.2|Tuberculosis of lung with cavitation
C0152566|ICD9CM|AB|011.20|TB lung w cavity-unspec
C0152566|ICD9CM|PT|011.20|Tuberculosis of lung with cavitation, unspecified
C0152567|ICD9CM|PT|011.21|Tuberculosis of lung with cavitation, bacteriological or histological examination not done
C0152567|ICD9CM|AB|011.21|TB lung w cavity-no exam
C0152568|ICD9CM|PT|011.22|Tuberculosis of lung with cavitation, bacteriological or histological examination unknown (at present)
C0152568|ICD9CM|AB|011.22|TB lung cavity-exam unkn
C0152569|ICD9CM|PT|011.23|Tuberculosis of lung with cavitation, tubercle bacilli found (in sputum) by microscopy
C0152569|ICD9CM|AB|011.23|TB lung w cavit-micro dx
C0152570|ICD9CM|PT|011.24|Tuberculosis of lung with cavitation, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152570|ICD9CM|AB|011.24|TB lung w cavity-cult dx
C0152571|ICD9CM|PT|011.25|Tuberculosis of lung with cavitation, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152571|ICD9CM|AB|011.25|TB lung w cavit-histo dx
C0152572|ICD9CM|PT|011.26|Tuberculosis of lung with cavitation, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152572|ICD9CM|AB|011.26|TB lung w cavit-oth test
C0152573|ICD9CM|HT|011.3|Tuberculosis of bronchus
C0152573|ICD9CM|AB|011.30|TB of bronchus-unspec
C0152573|ICD9CM|PT|011.30|Tuberculosis of bronchus, unspecified
C0152574|ICD9CM|PT|011.31|Tuberculosis of bronchus, bacteriological or histological examination not done
C0152574|ICD9CM|AB|011.31|TB of bronchus-no exam
C0152575|ICD9CM|PT|011.32|Tuberculosis of bronchus, bacteriological or histological examination unknown (at present)
C0152575|ICD9CM|AB|011.32|TB of bronchus-exam unkn
C0152576|ICD9CM|PT|011.33|Tuberculosis of bronchus, tubercle bacilli found (in sputum) by microscopy
C0152576|ICD9CM|AB|011.33|TB of bronchus-micro dx
C0152577|ICD9CM|PT|011.34|Tuberculosis of bronchus, tubercle bacilli not found (in sputum) by microscopy, but found in bacterial culture
C0152577|ICD9CM|AB|011.34|TB of bronchus-cult dx
C0152578|ICD9CM|PT|011.35|Tuberculosis of bronchus, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152578|ICD9CM|AB|011.35|TB of bronchus-histo dx
C0152579|ICD9CM|PT|011.36|Tuberculosis of bronchus, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152579|ICD9CM|AB|011.36|TB of bronchus-oth test
C0152580|ICD9CM|PT|011.41|Tuberculous fibrosis of lung, bacteriological or histological examination not done
C0152580|ICD9CM|AB|011.41|TB lung fibrosis-no exam
C0152581|ICD9CM|PT|011.42|Tuberculous fibrosis of lung, bacteriological or histological examination unknown (at present)
C0152581|ICD9CM|AB|011.42|TB lung fibros-exam unkn
C0152582|ICD9CM|PT|011.43|Tuberculous fibrosis of lung, tubercle bacilli found (in sputum) by microscopy
C0152582|ICD9CM|AB|011.43|TB lung fibros-micro dx
C0152583|ICD9CM|PT|011.44|Tuberculous fibrosis of lung, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152583|ICD9CM|AB|011.44|TB lung fibrosis-cult dx
C0152584|ICD9CM|PT|011.45|Tuberculous fibrosis of lung, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152584|ICD9CM|AB|011.45|TB lung fibros-histo dx
C0152585|ICD9CM|PT|011.46|Tuberculous fibrosis of lung, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152585|ICD9CM|AB|011.46|TB lung fibros-oth test
C0152586|ICD9CM|HT|011.5|Tuberculous bronchiectasis
C0152586|ICD9CM|AB|011.50|TB bronchiectasis-unspec
C0152586|ICD9CM|PT|011.50|Tuberculous bronchiectasis, unspecified
C0152587|ICD9CM|PT|011.51|Tuberculous bronchiectasis, bacteriological or histological examination not done
C0152587|ICD9CM|AB|011.51|TB bronchiect-no exam
C0152588|ICD9CM|PT|011.52|Tuberculous bronchiectasis, bacteriological or histological examination unknown (at present)
C0152588|ICD9CM|AB|011.52|TB bronchiect-exam unkn
C0152589|ICD9CM|PT|011.53|Tuberculous bronchiectasis, tubercle bacilli found (in sputum) by microscopy
C0152589|ICD9CM|AB|011.53|TB bronchiect-micro dx
C0152590|ICD9CM|PT|011.54|Tuberculous bronchiectasis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152590|ICD9CM|AB|011.54|TB bronchiect-cult dx
C0152591|ICD9CM|PT|011.55|Tuberculous bronchiectasis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152591|ICD9CM|AB|011.55|TB bronchiect-histo dx
C0152592|ICD9CM|PT|011.56|Tuberculous bronchiectasis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152592|ICD9CM|AB|011.56|TB bronchiect-oth test
C0152594|ICD9CM|PT|011.61|Tuberculous pneumonia [any form], bacteriological or histological examination not done
C0152594|ICD9CM|AB|011.61|TB pneumonia-no exam
C0152595|ICD9CM|PT|011.62|Tuberculous pneumonia [any form], bacteriological or histological examination unknown (at present)
C0152595|ICD9CM|AB|011.62|TB pneumonia-exam unkn
C0152596|ICD9CM|PT|011.63|Tuberculous pneumonia [any form], tubercle bacilli found (in sputum) by microscopy
C0152596|ICD9CM|AB|011.63|TB pneumonia-micro dx
C0152597|ICD9CM|PT|011.64|Tuberculous pneumonia [any form], tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152597|ICD9CM|AB|011.64|TB pneumonia-cult dx
C0152598|ICD9CM|PT|011.65|Tuberculous pneumonia [any form], tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152598|ICD9CM|AB|011.65|TB pneumonia-histo dx
C0152599|ICD9CM|PT|011.66|Tuberculous pneumonia [any form], tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152599|ICD9CM|AB|011.66|TB pneumonia-oth test
C0152600|ICD9CM|HT|011.7|Tuberculous pneumothorax
C0152600|ICD9CM|AB|011.70|TB pneumothorax-unspec
C0152600|ICD9CM|PT|011.70|Tuberculous pneumothorax, unspecified
C0152601|ICD9CM|PT|011.71|Tuberculous pneumothorax, bacteriological or histological examination not done
C0152601|ICD9CM|AB|011.71|TB pneumothorax-no exam
C0152602|ICD9CM|PT|011.72|Tuberculous pneumothorax, bacteriological or histological examination unknown (at present)
C0152602|ICD9CM|AB|011.72|TB pneumothorx-exam unkn
C0152603|ICD9CM|PT|011.73|Tuberculous pneumothorax, tubercle bacilli found (in sputum) by microscopy
C0152603|ICD9CM|AB|011.73|TB pneumothorax-micro dx
C0152604|ICD9CM|PT|011.74|Tuberculous pneumothorax, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152604|ICD9CM|AB|011.74|TB pneumothorax-cult dx
C0152605|ICD9CM|PT|011.75|Tuberculous pneumothorax, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152605|ICD9CM|AB|011.75|TB pneumothorax-histo dx
C0152606|ICD9CM|PT|011.76|Tuberculous pneumothorax, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152606|ICD9CM|AB|011.76|TB pneumothorax-oth test
C0152607|ICD9CM|HT|011.8|Other specified pulmonary tuberculosis
C0152608|ICD9CM|PT|011.81|Other specified pulmonary tuberculosis, bacteriological or histological examination not done
C0152608|ICD9CM|AB|011.81|Pulmonary TB NEC-no exam
C0152609|ICD9CM|PT|011.82|Other specified pulmonary tuberculosis, bacteriological or histological examination unknown (at present)
C0152609|ICD9CM|AB|011.82|Pulmon TB NEC-exam unkn
C0152610|ICD9CM|PT|011.83|Other specified pulmonary tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152610|ICD9CM|AB|011.83|Pulmon TB NEC-micro dx
C0152611|ICD9CM|PT|011.84|Other specified pulmonary tuberculosis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152611|ICD9CM|AB|011.84|Pulmon TB NEC-cult dx
C0152612|ICD9CM|PT|011.85|Other specified pulmonary tuberculosis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152612|ICD9CM|AB|011.85|Pulmon TB NEC-histo dx
C0152613|ICD9CM|PT|011.86|Other specified pulmonary tuberculosis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152613|ICD9CM|AB|011.86|Pulmon TB NEC-oth test
C0152614|ICD9CM|PT|011.91|Pulmonary tuberculosis, unspecified, bacteriological or histological examination not done
C0152614|ICD9CM|AB|011.91|Pulmonary TB NOS-no exam
C0152615|ICD9CM|PT|011.92|Pulmonary tuberculosis, unspecified, bacteriological or histological examination unknown (at present)
C0152615|ICD9CM|AB|011.92|Pulmon TB NOS-exam unkn
C0152616|ICD9CM|PT|011.93|Pulmonary tuberculosis, unspecified, tubercle bacilli found (in sputum) by microscopy
C0152616|ICD9CM|AB|011.93|Pulmon TB NOS-micro dx
C0152617|ICD9CM|PT|011.94|Pulmonary tuberculosis, unspecified, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152617|ICD9CM|AB|011.94|Pulmon TB NOS-cult dx
C0152618|ICD9CM|PT|011.95|Pulmonary tuberculosis, unspecified, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152618|ICD9CM|AB|011.95|Pulmon TB NOS-histo dx
C0152619|ICD9CM|PT|011.96|Pulmonary tuberculosis, unspecified, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152619|ICD9CM|AB|011.96|Pulmon TB NOS-oth test
C0152620|ICD9CM|HT|012|Other respiratory tuberculosis
C0152621|ICD9CM|PT|012.01|Tuberculous pleurisy, bacteriological or histological examination not done
C0152621|ICD9CM|AB|012.01|TB pleurisy-no exam
C0152622|ICD9CM|PT|012.02|Tuberculous pleurisy, bacteriological or histological examination unknown (at present)
C0152622|ICD9CM|AB|012.02|TB pleurisy-exam unkn
C0152623|ICD9CM|PT|012.03|Tuberculous pleurisy, tubercle bacilli found (in sputum) by microscopy
C0152623|ICD9CM|AB|012.03|TB pleurisy-micro dx
C0152624|ICD9CM|PT|012.04|Tuberculous pleurisy, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152624|ICD9CM|AB|012.04|TB pleurisy-cult dx
C0152625|ICD9CM|PT|012.05|Tuberculous pleurisy, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152625|ICD9CM|AB|012.05|TB pleurisy-histolog dx
C0152626|ICD9CM|PT|012.06|Tuberculous pleurisy, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152626|ICD9CM|AB|012.06|TB pleurisy-oth test
C0152627|ICD9CM|HT|012.1|Tuberculosis of intrathoracic lymph nodes
C0152627|ICD9CM|AB|012.10|TB thoracic nodes-unspec
C0152627|ICD9CM|PT|012.10|Tuberculosis of intrathoracic lymph nodes, unspecified
C0152628|ICD9CM|PT|012.11|Tuberculosis of intrathoracic lymph nodes, bacteriological or histological examination not done
C0152628|ICD9CM|AB|012.11|TB thorax node-no exam
C0152629|ICD9CM|PT|012.12|Tuberculosis of intrathoracic lymph nodes, bacteriological or histological examination unknown (at present)
C0152629|ICD9CM|AB|012.12|TB thorax node-exam unkn
C0152630|ICD9CM|PT|012.13|Tuberculosis of intrathoracic lymph nodes, tubercle bacilli found (in sputum) by microscopy
C0152630|ICD9CM|AB|012.13|TB thorax node-micro dx
C0152631|ICD9CM|PT|012.14|Tuberculosis of intrathoracic lymph nodes, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152631|ICD9CM|AB|012.14|TB thorax node-cult dx
C0152632|ICD9CM|PT|012.15|Tuberculosis of intrathoracic lymph nodes, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152632|ICD9CM|AB|012.15|TB thorax node-histo dx
C0152633|ICD9CM|PT|012.16|Tuberculosis of intrathoracic lymph nodes, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152633|ICD9CM|AB|012.16|TB thorax node-oth test
C0152634|ICD9CM|HT|012.2|Isolated tracheal or bronchial tuberculosis
C0152634|ICD9CM|AB|012.20|Isol tracheal tb-unspec
C0152634|ICD9CM|PT|012.20|Isolated tracheal or bronchial tuberculosis, unspecified
C0152635|ICD9CM|PT|012.21|Isolated tracheal or bronchial tuberculosis, bacteriological or histological examination not done
C0152635|ICD9CM|AB|012.21|Isol tracheal tb-no exam
C0152636|ICD9CM|PT|012.22|Isolated tracheal or bronchial tuberculosis, bacteriological or histological examination unknown (at present)
C0152636|ICD9CM|AB|012.22|Isol trach tb-exam unkn
C0152637|ICD9CM|PT|012.23|Isolated tracheal or bronchial tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152637|ICD9CM|AB|012.23|Isolat trach tb-micro dx
C0152638|ICD9CM|PT|012.24|Isolated tracheal or bronchial tuberculosis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152638|ICD9CM|AB|012.24|Isol tracheal tb-cult dx
C0152639|ICD9CM|PT|012.25|Isolated tracheal or bronchial tuberculosis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152639|ICD9CM|AB|012.25|Isolat trach tb-histo dx
C0152640|ICD9CM|PT|012.26|Isolated tracheal or bronchial tuberculosis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152640|ICD9CM|AB|012.26|Isolat trach tb-oth test
C0152641|ICD9CM|PT|012.31|Tuberculous laryngitis, bacteriological or histological examination not done
C0152641|ICD9CM|AB|012.31|TB laryngitis-no exam
C0152642|ICD9CM|PT|012.32|Tuberculous laryngitis, bacteriological or histological examination unknown (at present)
C0152642|ICD9CM|AB|012.32|TB laryngitis-exam unkn
C0152643|ICD9CM|PT|012.33|Tuberculous laryngitis, tubercle bacilli found (in sputum) by microscopy
C0152643|ICD9CM|AB|012.33|TB laryngitis-micro dx
C0152644|ICD9CM|PT|012.34|Tuberculous laryngitis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152644|ICD9CM|AB|012.34|TB laryngitis-cult dx
C0152645|ICD9CM|PT|012.35|Tuberculous laryngitis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152645|ICD9CM|AB|012.35|TB laryngitis-histo dx
C0152646|ICD9CM|PT|012.36|Tuberculous laryngitis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152646|ICD9CM|AB|012.36|TB laryngitis-oth test
C0152647|ICD9CM|PT|012.80|Other specified respiratory tuberculosis, unspecified
C0152647|ICD9CM|HT|012.8|Other specified respiratory tuberculosis
C0152647|ICD9CM|AB|012.80|Resp TB NEC-unspec
C0152648|ICD9CM|PT|012.81|Other specified respiratory tuberculosis, bacteriological or histological examination not done
C0152648|ICD9CM|AB|012.81|Resp TB NEC-no exam
C0152649|ICD9CM|PT|012.82|Other specified respiratory tuberculosis, bacteriological or histological examination unknown (at present)
C0152649|ICD9CM|AB|012.82|Resp TB NEC-exam unkn
C0152650|ICD9CM|PT|012.83|Other specified respiratory tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152650|ICD9CM|AB|012.83|Resp TB NEC-micro dx
C0152651|ICD9CM|PT|012.84|Other specified respiratory tuberculosis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152651|ICD9CM|AB|012.84|Resp TB NEC-cult dx
C0152652|ICD9CM|PT|012.85|Other specified respiratory tuberculosis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152652|ICD9CM|AB|012.85|Resp TB NEC-histo dx
C0152653|ICD9CM|PT|012.86|Other specified respiratory tuberculosis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152653|ICD9CM|AB|012.86|Resp TB NEC-oth test
C0152654|ICD9CM|HT|013|Tuberculosis of meninges and central nervous system
C0152655|ICD9CM|PT|013.01|Tuberculous meningitis, bacteriological or histological examination not done
C0152655|ICD9CM|AB|013.01|TB meningitis-no exam
C0152656|ICD9CM|PT|013.02|Tuberculous meningitis, bacteriological or histological examination unknown (at present)
C0152656|ICD9CM|AB|013.02|TB meningitis-exam unkn
C0152657|ICD9CM|PT|013.03|Tuberculous meningitis, tubercle bacilli found (in sputum) by microscopy
C0152657|ICD9CM|AB|013.03|TB meningitis-micro dx
C0152658|ICD9CM|PT|013.04|Tuberculous meningitis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152658|ICD9CM|AB|013.04|TB meningitis-cult dx
C0152659|ICD9CM|PT|013.05|Tuberculous meningitis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152659|ICD9CM|AB|013.05|TB meningitis-histo dx
C0152660|ICD9CM|PT|013.06|Tuberculous meningitis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152660|ICD9CM|AB|013.06|TB meningitis-oth test
C0152661|ICD9CM|HT|013.1|Tuberculoma of meninges
C0152661|ICD9CM|AB|013.10|Tubrclma meninges-unspec
C0152661|ICD9CM|PT|013.10|Tuberculoma of meninges, unspecified
C0152662|ICD9CM|PT|013.11|Tuberculoma of meninges, bacteriological or histological examination not done
C0152662|ICD9CM|AB|013.11|Tubrclma mening-no exam
C0152663|ICD9CM|PT|013.12|Tuberculoma of meninges, bacteriological or histological examination unknown (at present)
C0152663|ICD9CM|AB|013.12|Tubrclma menin-exam unkn
C0152664|ICD9CM|PT|013.13|Tuberculoma of meninges, tubercle bacilli found (in sputum) by microscopy
C0152664|ICD9CM|AB|013.13|Tubrclma mening-micro dx
C0152665|ICD9CM|PT|013.14|Tuberculoma of meninges, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152665|ICD9CM|AB|013.14|Tubrclma mening-cult dx
C0152666|ICD9CM|PT|013.15|Tuberculoma of meninges, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152666|ICD9CM|AB|013.15|Tubrclma mening-histo dx
C0152667|ICD9CM|PT|013.16|Tuberculoma of meninges, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152667|ICD9CM|AB|013.16|Tubrclma mening-oth test
C0152669|ICD9CM|PT|013.21|Tuberculoma of brain, bacteriological or histological examination not done
C0152669|ICD9CM|AB|013.21|Tubrcloma brain-no exam
C0152670|ICD9CM|PT|013.22|Tuberculoma of brain, bacteriological or histological examination unknown (at present)
C0152670|ICD9CM|AB|013.22|Tubrclma brain-exam unkn
C0152671|ICD9CM|PT|013.23|Tuberculoma of brain, tubercle bacilli found (in sputum) by microscopy
C0152671|ICD9CM|AB|013.23|Tubrcloma brain-micro dx
C0152672|ICD9CM|PT|013.24|Tuberculoma of brain, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152672|ICD9CM|AB|013.24|Tubrcloma brain-cult dx
C0152673|ICD9CM|PT|013.25|Tuberculoma of brain, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152673|ICD9CM|AB|013.25|Tubrcloma brain-histo dx
C0152674|ICD9CM|PT|013.26|Tuberculoma of brain, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152674|ICD9CM|AB|013.26|Tubrcloma brain-oth test
C0152676|ICD9CM|PT|013.31|Tuberculous abscess of brain, bacteriological or histological examination not done
C0152676|ICD9CM|AB|013.31|TB brain abscess-no exam
C0152677|ICD9CM|PT|013.32|Tuberculous abscess of brain, bacteriological or histological examination unknown (at present)
C0152677|ICD9CM|AB|013.32|TB brain absc-exam unkn
C0152678|ICD9CM|PT|013.33|Tuberculous abscess of brain, tubercle bacilli found (in sputum) by microscopy
C0152678|ICD9CM|AB|013.33|TB brain absc-micro dx
C0152679|ICD9CM|PT|013.34|Tuberculous abscess of brain, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152679|ICD9CM|AB|013.34|TB brain abscess-cult dx
C0152680|ICD9CM|PT|013.35|Tuberculous abscess of brain, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152680|ICD9CM|AB|013.35|TB brain absc-histo dx
C0152681|ICD9CM|PT|013.36|Tuberculous abscess of brain, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152681|ICD9CM|AB|013.36|TB brain absc-oth test
C0152683|ICD9CM|PT|013.41|Tuberculoma of spinal cord, bacteriological or histological examination not done
C0152683|ICD9CM|AB|013.41|Tubrclma sp cord-no exam
C0152684|ICD9CM|PT|013.42|Tuberculoma of spinal cord, bacteriological or histological examination unknown (at present)
C0152684|ICD9CM|AB|013.42|Tubrclma sp cd-exam unkn
C0152685|ICD9CM|PT|013.43|Tuberculoma of spinal cord, tubercle bacilli found (in sputum) by microscopy
C0152685|ICD9CM|AB|013.43|Tubrclma sp crd-micro dx
C0152686|ICD9CM|PT|013.44|Tuberculoma of spinal cord, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152686|ICD9CM|AB|013.44|Tubrclma sp cord-cult dx
C0152687|ICD9CM|PT|013.45|Tuberculoma of spinal cord, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152687|ICD9CM|AB|013.45|Tubrclma sp crd-histo dx
C0152688|ICD9CM|PT|013.46|Tuberculoma of spinal cord, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152688|ICD9CM|AB|013.46|Tubrclma sp crd-oth test
C0152690|ICD9CM|PT|013.51|Tuberculous abscess of spinal cord, bacteriological or histological examination not done
C0152690|ICD9CM|AB|013.51|TB sp crd absc-no exam
C0152691|ICD9CM|PT|013.52|Tuberculous abscess of spinal cord, bacteriological or histological examination unknown (at present)
C0152691|ICD9CM|AB|013.52|TB sp crd absc-exam unkn
C0152692|ICD9CM|PT|013.53|Tuberculous abscess of spinal cord, tubercle bacilli found (in sputum) by microscopy
C0152692|ICD9CM|AB|013.53|TB sp crd absc-micro dx
C0152693|ICD9CM|PT|013.54|Tuberculous abscess of spinal cord, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152693|ICD9CM|AB|013.54|TB sp crd absc-cult dx
C0152694|ICD9CM|PT|013.55|Tuberculous abscess of spinal cord, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152694|ICD9CM|AB|013.55|TB sp crd absc-histo dx
C0152695|ICD9CM|PT|013.56|Tuberculous abscess of spinal cord, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152695|ICD9CM|AB|013.56|TB sp crd absc-oth test
C0152696|ICD9CM|PT|013.60|Tuberculous encephalitis or myelitis, unspecified
C0152696|ICD9CM|HT|013.6|Tuberculous encephalitis or myelitis
C0152696|ICD9CM|AB|013.60|TB encephalitis-unspec
C0152697|ICD9CM|PT|013.61|Tuberculous encephalitis or myelitis, bacteriological or histological examination not done
C0152697|ICD9CM|AB|013.61|TB encephalitis-no exam
C0152698|ICD9CM|PT|013.62|Tuberculous encephalitis or myelitis, bacteriological or histological examination unknown (at present)
C0152698|ICD9CM|AB|013.62|TB encephalit-exam unkn
C0152699|ICD9CM|PT|013.63|Tuberculous encephalitis or myelitis, tubercle bacilli found (in sputum) by microscopy
C0152699|ICD9CM|AB|013.63|TB encephalitis-micro dx
C0152700|ICD9CM|PT|013.64|Tuberculous encephalitis or myelitis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152700|ICD9CM|AB|013.64|TB encephalitis-cult dx
C0152701|ICD9CM|PT|013.65|Tuberculous encephalitis or myelitis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152701|ICD9CM|AB|013.65|TB encephalitis-histo dx
C0152702|ICD9CM|PT|013.66|Tuberculous encephalitis or myelitis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152702|ICD9CM|AB|013.66|TB encephalitis-oth test
C0152703|ICD9CM|HT|013.8|Other specified tuberculosis of central nervous system
C0152704|ICD9CM|PT|013.81|Other specified tuberculosis of central nervous system, bacteriological or histological examination not done
C0152704|ICD9CM|AB|013.81|Cns TB NEC-no exam
C0152705|ICD9CM|PT|013.82|Other specified tuberculosis of central nervous system, bacteriological or histological examination unknown (at present)
C0152705|ICD9CM|AB|013.82|Cns TB NEC-exam unkn
C0152706|ICD9CM|PT|013.83|Other specified tuberculosis of central nervous system, tubercle bacilli found (in sputum) by microscopy
C0152706|ICD9CM|AB|013.83|Cns TB NEC-micro dx
C0152707|ICD9CM|PT|013.84|Other specified tuberculosis of central nervous system, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152707|ICD9CM|AB|013.84|Cns TB NEC-cult dx
C0152708|ICD9CM|PT|013.85|Other specified tuberculosis of central nervous system, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152708|ICD9CM|AB|013.85|Cns TB NEC-histo dx
C0152709|ICD9CM|PT|013.86|Other specified tuberculosis of central nervous system, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152709|ICD9CM|AB|013.86|Cns TB NEC-oth test
C0152711|ICD9CM|PT|013.91|Unspecified tuberculosis of central nervous system, bacteriological or histological examination not done
C0152711|ICD9CM|AB|013.91|Cns TB NOS-no exam
C0152712|ICD9CM|PT|013.92|Unspecified tuberculosis of central nervous system, bacteriological or histological examination unknown (at present)
C0152712|ICD9CM|AB|013.92|Cns TB NOS-exam unkn
C0152713|ICD9CM|PT|013.93|Unspecified tuberculosis of central nervous system, tubercle bacilli found (in sputum) by microscopy
C0152713|ICD9CM|AB|013.93|Cns TB NOS-micro dx
C0152714|ICD9CM|PT|013.94|Unspecified tuberculosis of central nervous system, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152714|ICD9CM|AB|013.94|Cns TB NOS-cult dx
C0152715|ICD9CM|PT|013.95|Unspecified tuberculosis of central nervous system, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152715|ICD9CM|AB|013.95|Cns TB NOS-histo dx
C0152716|ICD9CM|PT|013.96|Unspecified tuberculosis of central nervous system, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152716|ICD9CM|AB|013.96|Cns TB NOS-oth test
C0152717|ICD9CM|HT|014|Tuberculosis of intestines, peritoneum, and mesenteric glands
C0152718|ICD9CM|PT|014.01|Tuberculous peritonitis, bacteriological or histological examination not done
C0152718|ICD9CM|AB|014.01|TB peritonitis-no exam
C0152719|ICD9CM|PT|014.02|Tuberculous peritonitis, bacteriological or histological examination unknown (at present)
C0152719|ICD9CM|AB|014.02|TB peritonitis-exam unkn
C0152720|ICD9CM|PT|014.03|Tuberculous peritonitis, tubercle bacilli found (in sputum) by microscopy
C0152720|ICD9CM|AB|014.03|TB peritonitis-micro dx
C0152721|ICD9CM|PT|014.04|Tuberculous peritonitis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152721|ICD9CM|AB|014.04|TB peritonitis-cult dx
C0152722|ICD9CM|PT|014.05|Tuberculous peritonitis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152722|ICD9CM|AB|014.05|TB peritonitis-histo dx
C0152723|ICD9CM|PT|014.06|Tuberculous peritonitis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152723|ICD9CM|AB|014.06|TB peritonitis-oth test
C0152724|ICD9CM|HT|014.8|Tuberculosis of intestines and mesenteric glands
C0152725|ICD9CM|PT|014.81|Other tuberculosis of intestines, peritoneum, and mesenteric glands, bacteriological or histological examination not done
C0152725|ICD9CM|AB|014.81|Intestin TB NEC-no exam
C0152726|ICD9CM|PT|014.82|Other tuberculosis of intestines, peritoneum, and mesenteric glands, bacteriological or histological examination unknown (at present)
C0152726|ICD9CM|AB|014.82|Intest TB NEC-exam unkn
C0152727|ICD9CM|PT|014.83|Other tuberculosis of intestines, peritoneum, and mesenteric glands, tubercle bacilli found (in sputum) by microscopy
C0152727|ICD9CM|AB|014.83|Intestin TB NEC-micro dx
C0152728|ICD9CM|PT|014.84|Other tuberculosis of intestines, peritoneum, and mesenteric glands, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152728|ICD9CM|AB|014.84|Intestin TB NEC-cult dx
C0152729|ICD9CM|PT|014.85|Other tuberculosis of intestines, peritoneum, and mesenteric glands, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152729|ICD9CM|AB|014.85|Intestin TB NEC-histo dx
C0152730|ICD9CM|PT|014.86|Other tuberculosis of intestines, peritoneum, and mesenteric glands, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152730|ICD9CM|AB|014.86|Intestin TB NEC-oth test
C0152731|ICD9CM|PT|015.01|Tuberculosis of vertebral column, bacteriological or histological examination not done
C0152731|ICD9CM|AB|015.01|TB of vertebra-no exam
C0152732|ICD9CM|PT|015.02|Tuberculosis of vertebral column, bacteriological or histological examination unknown (at present)
C0152732|ICD9CM|AB|015.02|TB of vertebra-exam unkn
C0152733|ICD9CM|PT|015.03|Tuberculosis of vertebral column, tubercle bacilli found (in sputum) by microscopy
C0152733|ICD9CM|AB|015.03|TB of vertebra-micro dx
C0152734|ICD9CM|PT|015.04|Tuberculosis of vertebral column, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152734|ICD9CM|AB|015.04|TB of vertebra-cult dx
C0152735|ICD9CM|PT|015.05|Tuberculosis of vertebral column, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152735|ICD9CM|AB|015.05|TB of vertebra-histo dx
C0152736|ICD9CM|PT|015.06|Tuberculosis of vertebral column, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152736|ICD9CM|AB|015.06|TB of vertebra-oth test
C0152737|ICD9CM|HT|015.1|Tuberculosis of hip
C0152738|ICD9CM|PT|015.11|Tuberculosis of hip, bacteriological or histological examination not done
C0152738|ICD9CM|AB|015.11|TB of hip-no exam
C0152739|ICD9CM|PT|015.12|Tuberculosis of hip, bacteriological or histological examination unknown (at present)
C0152739|ICD9CM|AB|015.12|TB of hip-exam unkn
C0152740|ICD9CM|PT|015.13|Tuberculosis of hip, tubercle bacilli found (in sputum) by microscopy
C0152740|ICD9CM|AB|015.13|TB of hip-micro dx
C0152741|ICD9CM|PT|015.14|Tuberculosis of hip, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152741|ICD9CM|AB|015.14|TB of hip-cult dx
C0152742|ICD9CM|PT|015.15|Tuberculosis of hip, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152742|ICD9CM|AB|015.15|TB of hip-histo dx
C0152743|ICD9CM|PT|015.16|Tuberculosis of hip, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152743|ICD9CM|AB|015.16|TB of hip-oth test
C0152744|ICD9CM|HT|015.2|Tuberculosis of knee
C0152745|ICD9CM|PT|015.21|Tuberculosis of knee, bacteriological or histological examination not done
C0152745|ICD9CM|AB|015.21|TB of knee-no exam
C0152746|ICD9CM|PT|015.22|Tuberculosis of knee, bacteriological or histological examination unknown (at present)
C0152746|ICD9CM|AB|015.22|TB of knee-exam unkn
C0152747|ICD9CM|PT|015.23|Tuberculosis of knee, tubercle bacilli found (in sputum) by microscopy
C0152747|ICD9CM|AB|015.23|TB of knee-micro dx
C0152748|ICD9CM|PT|015.24|Tuberculosis of knee, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152748|ICD9CM|AB|015.24|TB of knee-cult dx
C0152749|ICD9CM|PT|015.25|Tuberculosis of knee, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152749|ICD9CM|AB|015.25|TB of knee-histo dx
C0152750|ICD9CM|PT|015.26|Tuberculosis of knee, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152750|ICD9CM|AB|015.26|TB of knee-oth test
C0152752|ICD9CM|PT|015.51|Tuberculosis of limb bones, bacteriological or histological examination not done
C0152752|ICD9CM|AB|015.51|TB limb bones-no exam
C0152753|ICD9CM|PT|015.52|Tuberculosis of limb bones, bacteriological or histological examination unknown (at present)
C0152753|ICD9CM|AB|015.52|TB limb bones-exam unkn
C0152754|ICD9CM|PT|015.53|Tuberculosis of limb bones, tubercle bacilli found (in sputum) by microscopy
C0152754|ICD9CM|AB|015.53|TB limb bones-micro dx
C0152755|ICD9CM|PT|015.54|Tuberculosis of limb bones, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152755|ICD9CM|AB|015.54|TB limb bones-cult dx
C0152756|ICD9CM|PT|015.55|Tuberculosis of limb bones, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152756|ICD9CM|AB|015.55|TB limb bones-histo dx
C0152757|ICD9CM|PT|015.56|Tuberculosis of limb bones, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152757|ICD9CM|AB|015.56|TB limb bones-oth test
C0152759|ICD9CM|PT|015.61|Tuberculosis of mastoid, bacteriological or histological examination not done
C0152759|ICD9CM|AB|015.61|TB of mastoid-no exam
C0152760|ICD9CM|PT|015.62|Tuberculosis of mastoid, bacteriological or histological examination unknown (at present)
C0152760|ICD9CM|AB|015.62|TB of mastoid-exam unkn
C0152761|ICD9CM|PT|015.63|Tuberculosis of mastoid, tubercle bacilli found (in sputum) by microscopy
C0152761|ICD9CM|AB|015.63|TB of mastoid-micro dx
C0152762|ICD9CM|PT|015.64|Tuberculosis of mastoid, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152762|ICD9CM|AB|015.64|TB of mastoid-cult dx
C0152763|ICD9CM|PT|015.65|Tuberculosis of mastoid, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152763|ICD9CM|AB|015.65|TB of mastoid-histo dx
C0152764|ICD9CM|PT|015.66|Tuberculosis of mastoid, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152764|ICD9CM|AB|015.66|TB of mastoid-oth test
C0152765|ICD9CM|HT|015.7|Tuberculosis of other specified bone
C0152766|ICD9CM|PT|015.71|Tuberculosis of other specified bone, bacteriological or histological examination not done
C0152766|ICD9CM|AB|015.71|TB of bone NEC-no exam
C0152767|ICD9CM|PT|015.72|Tuberculosis of other specified bone, bacteriological or histological examination unknown (at present)
C0152767|ICD9CM|AB|015.72|TB of bone NEC-exam unkn
C0152768|ICD9CM|PT|015.73|Tuberculosis of other specified bone, tubercle bacilli found (in sputum) by microscopy
C0152768|ICD9CM|AB|015.73|TB of bone NEC-micro dx
C0152769|ICD9CM|PT|015.74|Tuberculosis of other specified bone, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152769|ICD9CM|AB|015.74|TB of bone NEC-cult dx
C0152770|ICD9CM|PT|015.75|Tuberculosis of other specified bone, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152770|ICD9CM|AB|015.75|TB of bone NEC-histo dx
C0152771|ICD9CM|PT|015.76|Tuberculosis of other specified bone, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152771|ICD9CM|AB|015.76|TB of bone NEC-oth test
C0152772|ICD9CM|HT|015.8|Tuberculosis of other specified joint
C0152773|ICD9CM|PT|015.81|Tuberculosis of other specified joint, bacteriological or histological examination not done
C0152773|ICD9CM|AB|015.81|TB of joint NEC-no exam
C0152774|ICD9CM|PT|015.82|Tuberculosis of other specified joint, bacteriological or histological examination unknown (at present)
C0152774|ICD9CM|AB|015.82|TB joint NEC-exam unkn
C0152775|ICD9CM|PT|015.83|Tuberculosis of other specified joint, tubercle bacilli found (in sputum) by microscopy
C0152775|ICD9CM|AB|015.83|TB of joint NEC-micro dx
C0152776|ICD9CM|PT|015.84|Tuberculosis of other specified joint, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152776|ICD9CM|AB|015.84|TB of joint NEC-cult dx
C0152777|ICD9CM|PT|015.85|Tuberculosis of other specified joint, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152777|ICD9CM|AB|015.85|TB of joint NEC-histo dx
C0152778|ICD9CM|PT|015.86|Tuberculosis of other specified joint, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152778|ICD9CM|AB|015.86|TB of joint NEC-oth test
C0152780|ICD9CM|PT|015.91|Tuberculosis of unspecified bones and joints, bacteriological or histological examination not done
C0152780|ICD9CM|AB|015.91|TB bone/jt NOS-no exam
C0152781|ICD9CM|PT|015.92|Tuberculosis of unspecified bones and joints, bacteriological or histological examination unknown (at present)
C0152781|ICD9CM|AB|015.92|TB bone/jt NOS-exam unkn
C0152782|ICD9CM|PT|015.93|Tuberculosis of unspecified bones and joints, tubercle bacilli found (in sputum) by microscopy
C0152782|ICD9CM|AB|015.93|TB bone/jt NOS-micro dx
C0152783|ICD9CM|PT|015.94|Tuberculosis of unspecified bones and joints, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152783|ICD9CM|AB|015.94|TB bone/jt NOS-cult dx
C0152784|ICD9CM|PT|015.95|Tuberculosis of unspecified bones and joints, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152784|ICD9CM|AB|015.95|TB bone/jt NOS-histo dx
C0152785|ICD9CM|PT|015.96|Tuberculosis of unspecified bones and joints, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152785|ICD9CM|AB|015.96|TB bone/jt NOS-oth test
C0152787|ICD9CM|PT|016.01|Tuberculosis of kidney, bacteriological or histological examination not done
C0152787|ICD9CM|AB|016.01|TB of kidney-no exam
C0152788|ICD9CM|PT|016.02|Tuberculosis of kidney, bacteriological or histological examination unknown (at present)
C0152788|ICD9CM|AB|016.02|TB of kidney-exam unkn
C0152789|ICD9CM|PT|016.03|Tuberculosis of kidney, tubercle bacilli found (in sputum) by microscopy
C0152789|ICD9CM|AB|016.03|TB of kidney-micro dx
C0152790|ICD9CM|PT|016.04|Tuberculosis of kidney, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152790|ICD9CM|AB|016.04|TB of kidney-cult dx
C0152791|ICD9CM|PT|016.05|Tuberculosis of kidney, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152791|ICD9CM|AB|016.05|TB of kidney-histo dx
C0152792|ICD9CM|PT|016.06|Tuberculosis of kidney, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152792|ICD9CM|AB|016.06|TB of kidney-oth test
C0152793|ICD9CM|HT|016.1|Tuberculosis of bladder
C0152793|ICD9CM|AB|016.10|TB of bladder-unspec
C0152793|ICD9CM|PT|016.10|Tuberculosis of bladder, unspecified
C0152794|ICD9CM|PT|016.11|Tuberculosis of bladder, bacteriological or histological examination not done
C0152794|ICD9CM|AB|016.11|TB of bladder-no exam
C0152795|ICD9CM|PT|016.12|Tuberculosis of bladder, bacteriological or histological examination unknown (at present)
C0152795|ICD9CM|AB|016.12|TB of bladder-exam unkn
C0152796|ICD9CM|PT|016.13|Tuberculosis of bladder, tubercle bacilli found (in sputum) by microscopy
C0152796|ICD9CM|AB|016.13|TB of bladder-micro dx
C0152797|ICD9CM|PT|016.14|Tuberculosis of bladder, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152797|ICD9CM|AB|016.14|TB of bladder-cult dx
C0152798|ICD9CM|PT|016.15|Tuberculosis of bladder, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152798|ICD9CM|AB|016.15|TB of bladder-histo dx
C0152799|ICD9CM|PT|016.16|Tuberculosis of bladder, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152799|ICD9CM|AB|016.16|TB of bladder-oth test
C0152800|ICD9CM|HT|016.2|Tuberculosis of ureter
C0152801|ICD9CM|PT|016.21|Tuberculosis of ureter, bacteriological or histological examination not done
C0152801|ICD9CM|AB|016.21|TB of ureter-no exam
C0152802|ICD9CM|PT|016.22|Tuberculosis of ureter, bacteriological or histological examination unknown (at present)
C0152802|ICD9CM|AB|016.22|TB of ureter-exam unkn
C0152803|ICD9CM|PT|016.23|Tuberculosis of ureter, tubercle bacilli found (in sputum) by microscopy
C0152803|ICD9CM|AB|016.23|TB of ureter-micro dx
C0152804|ICD9CM|PT|016.24|Tuberculosis of ureter, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152804|ICD9CM|AB|016.24|TB of ureter-cult dx
C0152805|ICD9CM|PT|016.25|Tuberculosis of ureter, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152805|ICD9CM|AB|016.25|TB of ureter-histo dx
C0152806|ICD9CM|PT|016.26|Tuberculosis of ureter, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152806|ICD9CM|AB|016.26|TB of ureter-oth test
C0152808|ICD9CM|PT|016.31|Tuberculosis of other urinary organs, bacteriological or histological examination not done
C0152808|ICD9CM|AB|016.31|TB urinary NEC-no exam
C0152809|ICD9CM|PT|016.32|Tuberculosis of other urinary organs, bacteriological or histological examination unknown (at present)
C0152809|ICD9CM|AB|016.32|TB urinary NEC-exam unkn
C0152810|ICD9CM|PT|016.33|Tuberculosis of other urinary organs, tubercle bacilli found (in sputum) by microscopy
C0152810|ICD9CM|AB|016.33|TB urinary NEC-micro dx
C0152811|ICD9CM|PT|016.34|Tuberculosis of other urinary organs, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152811|ICD9CM|AB|016.34|TB urinary NEC-cult dx
C0152812|ICD9CM|PT|016.35|Tuberculosis of other urinary organs, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152812|ICD9CM|AB|016.35|TB urinary NEC-histo dx
C0152813|ICD9CM|PT|016.36|Tuberculosis of other urinary organs, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152813|ICD9CM|AB|016.36|TB urinary NEC-oth test
C0152814|ICD9CM|HT|016.4|Tuberculosis of epididymis
C0152815|ICD9CM|PT|016.41|Tuberculosis of epididymis, bacteriological or histological examination not done
C0152815|ICD9CM|AB|016.41|TB epididymis-no exam
C0152816|ICD9CM|PT|016.42|Tuberculosis of epididymis, bacteriological or histological examination unknown (at present)
C0152816|ICD9CM|AB|016.42|TB epididymis-exam unkn
C0152817|ICD9CM|PT|016.43|Tuberculosis of epididymis, tubercle bacilli found (in sputum) by microscopy
C0152817|ICD9CM|AB|016.43|TB epididymis-micro dx
C0152818|ICD9CM|PT|016.44|Tuberculosis of epididymis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152818|ICD9CM|AB|016.44|TB epididymis-cult dx
C0152819|ICD9CM|PT|016.45|Tuberculosis of epididymis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152819|ICD9CM|AB|016.45|TB epididymis-histo dx
C0152820|ICD9CM|PT|016.46|Tuberculosis of epididymis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152820|ICD9CM|AB|016.46|TB epididymis-oth test
C0152821|ICD9CM|HT|016.5|Tuberculosis of other male genital organs
C0152821|ICD9CM|AB|016.50|TB male genit NEC-unspec
C0152821|ICD9CM|PT|016.50|Tuberculosis of other male genital organs, unspecified
C0152822|ICD9CM|PT|016.51|Tuberculosis of other male genital organs, bacteriological or histological examination not done
C0152822|ICD9CM|AB|016.51|TB male gen NEC-no exam
C0152823|ICD9CM|PT|016.52|Tuberculosis of other male genital organs, bacteriological or histological examination unknown (at present)
C0152823|ICD9CM|AB|016.52|TB male gen NEC-ex unkn
C0152824|ICD9CM|PT|016.53|Tuberculosis of other male genital organs, tubercle bacilli found (in sputum) by microscopy
C0152824|ICD9CM|AB|016.53|TB male gen NEC-micro dx
C0152825|ICD9CM|PT|016.54|Tuberculosis of other male genital organs, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152825|ICD9CM|AB|016.54|TB male gen NEC-cult dx
C0152826|ICD9CM|PT|016.55|Tuberculosis of other male genital organs, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152826|ICD9CM|AB|016.55|TB male gen NEC-histo dx
C0152827|ICD9CM|PT|016.56|Tuberculosis of other male genital organs, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152827|ICD9CM|AB|016.56|TB male gen NEC-oth test
C0152828|ICD9CM|HT|016.6|Tuberculous oophoritis and salpingitis
C0152829|ICD9CM|PT|016.61|Tuberculous oophoritis and salpingitis, bacteriological or histological examination not done
C0152829|ICD9CM|AB|016.61|TB ovary & tube-no exam
C0152830|ICD9CM|PT|016.62|Tuberculous oophoritis and salpingitis, bacteriological or histological examination unknown (at present)
C0152830|ICD9CM|AB|016.62|TB ovary/tube-exam unkn
C0152831|ICD9CM|PT|016.63|Tuberculous oophoritis and salpingitis, tubercle bacilli found (in sputum) by microscopy
C0152831|ICD9CM|AB|016.63|TB ovary & tube-micro dx
C0152832|ICD9CM|PT|016.64|Tuberculous oophoritis and salpingitis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152832|ICD9CM|AB|016.64|TB ovary & tube-cult dx
C0152833|ICD9CM|PT|016.65|Tuberculous oophoritis and salpingitis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152833|ICD9CM|AB|016.65|TB ovary & tube-histo dx
C0152834|ICD9CM|PT|016.66|Tuberculous oophoritis and salpingitis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152834|ICD9CM|AB|016.66|TB ovary & tube-oth test
C0152835|ICD9CM|HT|016.7|Tuberculosis of other female genital organs
C0152835|ICD9CM|AB|016.70|TB female gen NEC-unspec
C0152835|ICD9CM|PT|016.70|Tuberculosis of other female genital organs, unspecified
C0152836|ICD9CM|PT|016.71|Tuberculosis of other female genital organs, bacteriological or histological examination not done
C0152836|ICD9CM|AB|016.71|TB fem gen NEC-no exam
C0152837|ICD9CM|PT|016.72|Tuberculosis of other female genital organs, bacteriological or histological examination unknown (at present)
C0152837|ICD9CM|AB|016.72|TB fem gen NEC-exam unkn
C0152838|ICD9CM|PT|016.73|Tuberculosis of other female genital organs, tubercle bacilli found (in sputum) by microscopy
C0152838|ICD9CM|AB|016.73|TB fem gen NEC-micro dx
C0152839|ICD9CM|PT|016.74|Tuberculosis of other female genital organs, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152839|ICD9CM|AB|016.74|TB fem gen NEC-cult dx
C0152840|ICD9CM|PT|016.75|Tuberculosis of other female genital organs, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152840|ICD9CM|AB|016.75|TB fem gen NEC-histo dx
C0152841|ICD9CM|PT|016.76|Tuberculosis of other female genital organs, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152841|ICD9CM|AB|016.76|TB fem gen NEC-oth test
C0152843|ICD9CM|PT|016.91|Genitourinary tuberculosis, unspecified, bacteriological or histological examination not done
C0152843|ICD9CM|AB|016.91|Gu TB NOS-no exam
C0152844|ICD9CM|PT|016.92|Genitourinary tuberculosis, unspecified, bacteriological or histological examination unknown (at present)
C0152844|ICD9CM|AB|016.92|Gu TB NOS-exam unkn
C0152845|ICD9CM|PT|016.93|Genitourinary tuberculosis, unspecified, tubercle bacilli found (in sputum) by microscopy
C0152845|ICD9CM|AB|016.93|Gu TB NOS-micro dx
C0152846|ICD9CM|PT|016.94|Genitourinary tuberculosis, unspecified, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152846|ICD9CM|AB|016.94|Gu TB NOS-cult dx
C0152847|ICD9CM|PT|016.95|Genitourinary tuberculosis, unspecified, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152847|ICD9CM|AB|016.95|Gu TB NOS-histo dx
C0152848|ICD9CM|PT|016.96|Genitourinary tuberculosis, unspecified, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152848|ICD9CM|AB|016.96|Gu TB NOS-oth test
C0152849|ICD9CM|PT|017.01|Tuberculosis of skin and subcutaneous cellular tissue, bacteriological or histological examination not done
C0152849|ICD9CM|AB|017.01|TB skin/subcut-no exam
C0152850|ICD9CM|PT|017.02|Tuberculosis of skin and subcutaneous cellular tissue, bacteriological or histological examination unknown (at present)
C0152850|ICD9CM|AB|017.02|TB skin/subcut-exam unkn
C0152851|ICD9CM|PT|017.03|Tuberculosis of skin and subcutaneous cellular tissue, tubercle bacilli found (in sputum) by microscopy
C0152851|ICD9CM|AB|017.03|TB skin/subcut-micro dx
C0152852|ICD9CM|PT|017.04|Tuberculosis of skin and subcutaneous cellular tissue, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152852|ICD9CM|AB|017.04|TB skin/subcut-cult dx
C0152853|ICD9CM|PT|017.05|Tuberculosis of skin and subcutaneous cellular tissue, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152853|ICD9CM|AB|017.05|TB skin/subcut-histo dx
C0152854|ICD9CM|PT|017.06|Tuberculosis of skin and subcutaneous cellular tissue, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152854|ICD9CM|AB|017.06|TB skin/subcut-oth test
C0152855|ICD9CM|PT|017.11|Erythema nodosum with hypersensitivity reaction in tuberculosis, bacteriological or histological examination not done
C0152855|ICD9CM|AB|017.11|Erythem nodos tb-no exam
C0152856|ICD9CM|PT|017.12|Erythema nodosum with hypersensitivity reaction in tuberculosis, bacteriological or histological examination unknown (at present)
C0152856|ICD9CM|AB|017.12|Erythem nod tb-exam unkn
C0152857|ICD9CM|PT|017.13|Erythema nodosum with hypersensitivity reaction in tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152857|ICD9CM|AB|017.13|Erythem nod tb-micro dx
C0152858|ICD9CM|PT|017.14|Erythema nodosum with hypersensitivity reaction in tuberculosis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152858|ICD9CM|AB|017.14|Erythem nodos tb-cult dx
C0152859|ICD9CM|PT|017.15|Erythema nodosum with hypersensitivity reaction in tuberculosis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152859|ICD9CM|AB|017.15|Erythem nod tb-histo dx
C0152860|ICD9CM|PT|017.16|Erythema nodosum with hypersensitivity reaction in tuberculosis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152860|ICD9CM|AB|017.16|Erythem nod tb-oth test
C0152861|ICD9CM|HT|017.2|Tuberculosis of peripheral lymph nodes
C0152861|ICD9CM|AB|017.20|TB periph lymph-unspec
C0152861|ICD9CM|PT|017.20|Tuberculosis of peripheral lymph nodes, unspecified
C0152862|ICD9CM|PT|017.21|Tuberculosis of peripheral lymph nodes, bacteriological or histological examination not done
C0152862|ICD9CM|AB|017.21|TB periph lymph-no exam
C0152863|ICD9CM|PT|017.22|Tuberculosis of peripheral lymph nodes, bacteriological or histological examination unknown (at present)
C0152863|ICD9CM|AB|017.22|TB periph lymph-exam unk
C0152864|ICD9CM|PT|017.23|Tuberculosis of peripheral lymph nodes, tubercle bacilli found (in sputum) by microscopy
C0152864|ICD9CM|AB|017.23|TB periph lymph-micro dx
C0152865|ICD9CM|PT|017.24|Tuberculosis of peripheral lymph nodes, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152865|ICD9CM|AB|017.24|TB periph lymph-cult dx
C0152866|ICD9CM|PT|017.25|Tuberculosis of peripheral lymph nodes, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152866|ICD9CM|AB|017.25|TB periph lymph-histo dx
C0152867|ICD9CM|PT|017.26|Tuberculosis of peripheral lymph nodes, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152867|ICD9CM|AB|017.26|TB periph lymph-oth test
C0152868|ICD9CM|PT|017.31|Tuberculosis of eye, bacteriological or histological examination not done
C0152868|ICD9CM|AB|017.31|TB of eye-no exam
C0152869|ICD9CM|PT|017.32|Tuberculosis of eye, bacteriological or histological examination unknown (at present)
C0152869|ICD9CM|AB|017.32|TB of eye-exam unkn
C0152870|ICD9CM|PT|017.33|Tuberculosis of eye, tubercle bacilli found (in sputum) by microscopy
C0152870|ICD9CM|AB|017.33|TB of eye-micro dx
C0152871|ICD9CM|PT|017.34|Tuberculosis of eye, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152871|ICD9CM|AB|017.34|TB of eye-cult dx
C0152872|ICD9CM|PT|017.35|Tuberculosis of eye, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152872|ICD9CM|AB|017.35|TB of eye-histo dx
C0152873|ICD9CM|PT|017.36|Tuberculosis of eye, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152873|ICD9CM|AB|017.36|TB of eye-oth test
C0152874|ICD9CM|HT|017.4|Tuberculosis of ear
C0152875|ICD9CM|PT|017.41|Tuberculosis of ear, bacteriological or histological examination not done
C0152875|ICD9CM|AB|017.41|TB of ear-no exam
C0152876|ICD9CM|PT|017.42|Tuberculosis of ear, bacteriological or histological examination unknown (at present)
C0152876|ICD9CM|AB|017.42|TB of ear-exam unkn
C0152877|ICD9CM|PT|017.43|Tuberculosis of ear, tubercle bacilli found (in sputum) by microscopy
C0152877|ICD9CM|AB|017.43|TB of ear-micro dx
C0152878|ICD9CM|PT|017.44|Tuberculosis of ear, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152878|ICD9CM|AB|017.44|TB of ear-cult dx
C0152879|ICD9CM|PT|017.45|Tuberculosis of ear, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152879|ICD9CM|AB|017.45|TB of ear-histo dx
C0152880|ICD9CM|PT|017.46|Tuberculosis of ear, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152880|ICD9CM|AB|017.46|TB of ear-oth test
C0152881|ICD9CM|HT|017.5|Tuberculosis of thyroid gland
C0152882|ICD9CM|PT|017.50|Tuberculosis of thyroid gland, unspecified
C0152882|ICD9CM|AB|017.50|TB of thyroid-unspec
C0152883|ICD9CM|PT|017.51|Tuberculosis of thyroid gland, bacteriological or histological examination not done
C0152883|ICD9CM|AB|017.51|TB of thyroid-no exam
C0152884|ICD9CM|PT|017.52|Tuberculosis of thyroid gland, bacteriological or histological examination unknown (at present)
C0152884|ICD9CM|AB|017.52|TB of thyroid-exam unkn
C0152885|ICD9CM|PT|017.53|Tuberculosis of thyroid gland, tubercle bacilli found (in sputum) by microscopy
C0152885|ICD9CM|AB|017.53|TB of thyroid-micro dx
C0152886|ICD9CM|PT|017.54|Tuberculosis of thyroid gland, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152886|ICD9CM|AB|017.54|TB of thyroid-cult dx
C0152887|ICD9CM|PT|017.55|Tuberculosis of thyroid gland, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152887|ICD9CM|AB|017.55|TB of thyroid-histo dx
C0152888|ICD9CM|PT|017.56|Tuberculosis of thyroid gland, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152888|ICD9CM|AB|017.56|TB of thyroid-oth test
C0152889|ICD9CM|HT|017.6|Tuberculosis of adrenal glands
C0152889|ICD9CM|AB|017.60|TB of adrenal-unspec
C0152889|ICD9CM|PT|017.60|Tuberculosis of adrenal glands, unspecified
C0152890|ICD9CM|PT|017.61|Tuberculosis of adrenal glands, bacteriological or histological examination not done
C0152890|ICD9CM|AB|017.61|TB of adrenal-no exam
C0152891|ICD9CM|PT|017.62|Tuberculosis of adrenal glands, bacteriological or histological examination unknown (at present)
C0152891|ICD9CM|AB|017.62|TB of adrenal-exam unkn
C0152892|ICD9CM|PT|017.63|Tuberculosis of adrenal glands, tubercle bacilli found (in sputum) by microscopy
C0152892|ICD9CM|AB|017.63|TB of adrenal-micro dx
C0152893|ICD9CM|PT|017.64|Tuberculosis of adrenal glands, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152893|ICD9CM|AB|017.64|TB of adrenal-cult dx
C0152894|ICD9CM|PT|017.65|Tuberculosis of adrenal glands, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152894|ICD9CM|AB|017.65|TB of adrenal-histo dx
C0152895|ICD9CM|PT|017.66|Tuberculosis of adrenal glands, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152895|ICD9CM|AB|017.66|TB of adrenal-oth test
C0152896|ICD9CM|PT|017.71|Tuberculosis of spleen, bacteriological or histological examination not done
C0152896|ICD9CM|AB|017.71|TB of spleen-no exam
C0152897|ICD9CM|PT|017.72|Tuberculosis of spleen, bacteriological or histological examination unknown (at present)
C0152897|ICD9CM|AB|017.72|TB of spleen-exam unkn
C0152898|ICD9CM|PT|017.73|Tuberculosis of spleen, tubercle bacilli found (in sputum) by microscopy
C0152898|ICD9CM|AB|017.73|TB of spleen-micro dx
C0152899|ICD9CM|PT|017.74|Tuberculosis of spleen, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152899|ICD9CM|AB|017.74|TB of spleen-cult dx
C0152900|ICD9CM|PT|017.75|Tuberculosis of spleen, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152900|ICD9CM|AB|017.75|TB of spleen-histo dx
C0152901|ICD9CM|PT|017.76|Tuberculosis of spleen, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152901|ICD9CM|AB|017.76|TB of spleen-oth test
C0152902|ICD9CM|HT|017.8|Tuberculosis of esophagus
C0152903|ICD9CM|PT|017.81|Tuberculosis of esophagus, bacteriological or histological examination not done
C0152903|ICD9CM|AB|017.81|TB esophagus-no exam
C0152904|ICD9CM|PT|017.82|Tuberculosis of esophagus, bacteriological or histological examination unknown (at present)
C0152904|ICD9CM|AB|017.82|TB esophagus-exam unkn
C0152905|ICD9CM|PT|017.83|Tuberculosis of esophagus, tubercle bacilli found (in sputum) by microscopy
C0152905|ICD9CM|AB|017.83|TB esophagus-micro dx
C0152906|ICD9CM|PT|017.84|Tuberculosis of esophagus, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152906|ICD9CM|AB|017.84|TB esophagus-cult dx
C0152907|ICD9CM|PT|017.85|Tuberculosis of esophagus, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152907|ICD9CM|AB|017.85|TB esophagus-histo dx
C0152908|ICD9CM|PT|017.86|Tuberculosis of esophagus, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152908|ICD9CM|AB|017.86|TB esophagus-oth test
C0152909|ICD9CM|PT|017.91|Tuberculosis of other specified organs, bacteriological or histological examination not done
C0152909|ICD9CM|AB|017.91|TB of organ NEC-no exam
C0152910|ICD9CM|PT|017.92|Tuberculosis of other specified organs, bacteriological or histological examination unknown (at present)
C0152910|ICD9CM|AB|017.92|TB organ NEC-exam unkn
C0152911|ICD9CM|PT|017.93|Tuberculosis of other specified organs, tubercle bacilli found (in sputum) by microscopy
C0152911|ICD9CM|AB|017.93|TB of organ NEC-micro dx
C0152912|ICD9CM|PT|017.94|Tuberculosis of other specified organs, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152912|ICD9CM|AB|017.94|TB of organ NEC-cult dx
C0152913|ICD9CM|PT|017.95|Tuberculosis of other specified organs, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152913|ICD9CM|AB|017.95|TB of organ NEC-histo dx
C0152914|ICD9CM|PT|017.96|Tuberculosis of other specified organs, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152914|ICD9CM|AB|017.96|TB of organ NEC-oth test
C0152915|ICD9CM|HT|018.0|Acute miliary tuberculosis
C0152915|ICD9CM|PT|018.00|Acute miliary tuberculosis, unspecified
C0152915|ICD9CM|AB|018.00|Acute miliary tb-unspec
C0152916|ICD9CM|PT|018.01|Acute miliary tuberculosis, bacteriological or histological examination not done
C0152916|ICD9CM|AB|018.01|Acute miliary tb-no exam
C0152917|ICD9CM|PT|018.02|Acute miliary tuberculosis, bacteriological or histological examination unknown (at present)
C0152917|ICD9CM|AB|018.02|Ac miliary tb-exam unkn
C0152918|ICD9CM|PT|018.03|Acute miliary tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152918|ICD9CM|AB|018.03|Ac miliary tb-micro dx
C0152919|ICD9CM|PT|018.04|Acute miliary tuberculosis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152919|ICD9CM|AB|018.04|Acute miliary tb-cult dx
C0152920|ICD9CM|PT|018.05|Acute miliary tuberculosis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152920|ICD9CM|AB|018.05|Ac miliary tb-histo dx
C0152921|ICD9CM|PT|018.06|Acute miliary tuberculosis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152921|ICD9CM|AB|018.06|Ac miliary tb-oth test
C0152922|ICD9CM|PT|018.80|Other specified miliary tuberculosis, unspecified
C0152922|ICD9CM|HT|018.8|Other specified miliary tuberculosis
C0152922|ICD9CM|AB|018.80|Miliary TB NEC-unspec
C0152923|ICD9CM|PT|018.81|Other specified miliary tuberculosis, bacteriological or histological examination not done
C0152923|ICD9CM|AB|018.81|Miliary TB NEC-no exam
C0152924|ICD9CM|PT|018.82|Other specified miliary tuberculosis, bacteriological or histological examination unknown (at present)
C0152924|ICD9CM|AB|018.82|Miliary TB NEC-exam unkn
C0152925|ICD9CM|PT|018.83|Other specified miliary tuberculosis, tubercle bacilli found (in sputum) by microscopy
C0152925|ICD9CM|AB|018.83|Miliary TB NEC-micro dx
C0152926|ICD9CM|PT|018.84|Other specified miliary tuberculosis, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152926|ICD9CM|AB|018.84|Miliary TB NEC-cult dx
C0152927|ICD9CM|PT|018.85|Other specified miliary tuberculosis, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152927|ICD9CM|AB|018.85|Miliary TB NEC-histo dx
C0152928|ICD9CM|PT|018.86|Other specified miliary tuberculosis, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152928|ICD9CM|AB|018.86|Miliary TB NEC-oth test
C0152929|ICD9CM|PT|018.91|Miliary tuberculosis, unspecified, bacteriological or histological examination not done
C0152929|ICD9CM|AB|018.91|Miliary TB NOS-no exam
C0152930|ICD9CM|PT|018.92|Miliary tuberculosis, unspecified, bacteriological or histological examination unknown (at present)
C0152930|ICD9CM|AB|018.92|Miliary TB NOS-exam unkn
C0152931|ICD9CM|PT|018.93|Miliary tuberculosis, unspecified, tubercle bacilli found (in sputum) by microscopy
C0152931|ICD9CM|AB|018.93|Miliary TB NOS-micro dx
C0152932|ICD9CM|PT|018.94|Miliary tuberculosis, unspecified, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0152932|ICD9CM|AB|018.94|Miliary TB NOS-cult dx
C0152933|ICD9CM|PT|018.95|Miliary tuberculosis, unspecified, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0152933|ICD9CM|AB|018.95|Miliary TB NOS-histo dx
C0152934|ICD9CM|PT|018.96|Miliary tuberculosis, unspecified, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0152934|ICD9CM|AB|018.96|Miliary TB NOS-oth test
C0152935|ICD9CM|AB|020.1|Cellulocutaneous plague
C0152935|ICD9CM|PT|020.1|Cellulocutaneous plague
C0152936|ICD9CM|AB|020.2|Septicemic plague
C0152936|ICD9CM|PT|020.2|Septicemic plague
C0152937|ICD9CM|AB|020.3|Primary pneumonic plague
C0152937|ICD9CM|PT|020.3|Primary pneumonic plague
C0152938|ICD9CM|PT|020.4|Secondary pneumonic plague
C0152938|ICD9CM|AB|020.4|Secondary pneumon plague
C0152940|ICD9CM|PT|020.8|Other specified types of plague
C0152940|ICD9CM|AB|020.8|Other types of plague
C0152941|ICD9CM|PT|021.0|Ulceroglandular tularemia
C0152941|ICD9CM|AB|021.0|Ulceroglandul tularemia
C0152942|ICD9CM|AB|021.1|Enteric tularemia
C0152942|ICD9CM|PT|021.1|Enteric tularemia
C0152944|ICD9CM|AB|021.3|Oculoglandular tularemia
C0152944|ICD9CM|PT|021.3|Oculoglandular tularemia
C0152945|ICD9CM|AB|022.2|Gastrointestinal anthrax
C0152945|ICD9CM|PT|022.2|Gastrointestinal anthrax
C0152946|ICD9CM|AB|022.3|Anthrax septicemia
C0152946|ICD9CM|PT|022.3|Anthrax septicemia
C0152947|ICD9CM|PT|022.8|Other specified manifestations of anthrax
C0152947|ICD9CM|AB|022.8|Other anthrax manifest
C0152948|ICD9CM|HT|027|Other zoonotic bacterial diseases
C0152949|ICD9CM|PT|027.8|Other specified zoonotic bacterial diseases
C0152949|ICD9CM|AB|027.8|Zoonotic bact dis NEC
C0152950|ICD9CM|HT|031|Diseases due to other mycobacteria
C0152951|ICD9CM|PT|031.8|Other specified mycobacterial diseases
C0152951|ICD9CM|AB|031.8|Mycobacterial dis NEC
C0152952|ICD9CM|AB|032.82|Diphtheritic myocarditis
C0152952|ICD9CM|PT|032.82|Diphtheritic myocarditis
C0152953|ICD9CM|AB|032.83|Diphtheritic peritonitis
C0152953|ICD9CM|PT|032.83|Diphtheritic peritonitis
C0152954|ICD9CM|AB|032.84|Diphtheritic cystitis
C0152954|ICD9CM|PT|032.84|Diphtheritic cystitis
C0152957|ICD9CM|PT|036.1|Meningococcal encephalitis
C0152957|ICD9CM|AB|036.1|Meningococc encephalitis
C0152958|ICD9CM|HT|036.4|Meningococcal carditis
C0152958|ICD9CM|PT|036.40|Meningococcal carditis, unspecified
C0152958|ICD9CM|AB|036.40|Meningococc carditis NOS
C0152959|ICD9CM|PT|036.41|Meningococcal pericarditis
C0152959|ICD9CM|AB|036.41|Meningococc pericarditis
C0152960|ICD9CM|PT|036.42|Meningococcal endocarditis
C0152960|ICD9CM|AB|036.42|Meningococc endocarditis
C0152961|ICD9CM|PT|036.43|Meningococcal myocarditis
C0152961|ICD9CM|AB|036.43|Meningococc myocarditis
C0152962|ICD9CM|PT|036.81|Meningococcal optic neuritis
C0152962|ICD9CM|AB|036.81|Meningococc optic neurit
C0152964|ICD9CM|AB|038.0|Streptococcal septicemia
C0152964|ICD9CM|PT|038.0|Streptococcal septicemia
C0152965|ICD9CM|HT|038.1|Staphylococcal septicemia
C0152965|ICD9CM|PT|038.10|Staphylococcal septicemia, unspecified
C0152965|ICD9CM|AB|038.10|Staphylcocc septicem NOS
C0152966|ICD9CM|AB|038.2|Pneumococcal septicemia
C0152966|ICD9CM|PT|038.2|Pneumococcal septicemia [Streptococcus pneumoniae septicemia]
C0152967|ICD9CM|PT|038.3|Septicemia due to anaerobes
C0152967|ICD9CM|AB|038.3|Anaerobic septicemia
C0152972|ICD9CM|PT|038.43|Septicemia due to pseudomonas
C0152972|ICD9CM|AB|038.43|Pseudomonas septicemia
C0152973|ICD9CM|PT|038.44|Septicemia due to serratia
C0152973|ICD9CM|AB|038.44|Serratia septicemia
C0152977|ICD9CM|PT|040.89|Other specified bacterial diseases
C0152977|ICD9CM|HT|040.8|Other specified bacterial disease
C0152977|ICD9CM|AB|040.89|Bacterial diseases NEC
C0152989|ICD9CM|PT|045.00|Acute paralytic poliomyelitis specified as bulbar, poliovirus, unspecified type
C0152989|ICD9CM|AB|045.00|Ac bulbar polio-type NOS
C0152990|ICD9CM|PT|045.01|Acute paralytic poliomyelitis specified as bulbar, poliovirus type I
C0152990|ICD9CM|AB|045.01|Ac bulbar polio-type 1
C0152991|ICD9CM|PT|045.02|Acute paralytic poliomyelitis specified as bulbar, poliovirus type II
C0152991|ICD9CM|AB|045.02|Ac bulbar polio-type 2
C0152992|ICD9CM|PT|045.03|Acute paralytic poliomyelitis specified as bulbar, poliovirus type III
C0152992|ICD9CM|AB|045.03|Ac bulbar polio-type 3
C0152993|ICD9CM|HT|045.1|Acute poliomyelitis with other paralysis
C0152994|ICD9CM|PT|045.10|Acute poliomyelitis with other paralysis, poliovirus, unspecified type
C0152994|ICD9CM|AB|045.10|Paral polio NEC-type NOS
C0152995|ICD9CM|PT|045.11|Acute poliomyelitis with other paralysis, poliovirus type I
C0152995|ICD9CM|AB|045.11|Paral polio NEC-type 1
C0152996|ICD9CM|PT|045.12|Acute poliomyelitis with other paralysis, poliovirus type II
C0152996|ICD9CM|AB|045.12|Paral polio NEC-type 2
C0152997|ICD9CM|PT|045.13|Acute poliomyelitis with other paralysis, poliovirus type III
C0152997|ICD9CM|AB|045.13|Paral polio NEC-type 3
C0152998|ICD9CM|HT|045.2|Acute nonparalytic poliomyelitis
C0152998|ICD9CM|PT|045.20|Acute nonparalytic poliomyelitis, poliovirus, unspecified type
C0152998|ICD9CM|AB|045.20|Nonparaly polio-type NOS
C0153004|ICD9CM|PT|045.91|Acute poliomyelitis, unspecified, poliovirus type I
C0153004|ICD9CM|AB|045.91|Ac polio NOS-type 1
C0153005|ICD9CM|PT|045.92|Acute poliomyelitis, unspecified, poliovirus type II
C0153005|ICD9CM|AB|045.92|Ac polio NOS-type 2
C0153006|ICD9CM|PT|045.93|Acute poliomyelitis, unspecified, poliovirus type III
C0153006|ICD9CM|AB|045.93|Ac polio NOS-type 3
C0153007|ICD9CM|PT|046.8|Other specified slow virus infection of central nervous system
C0153007|ICD9CM|AB|046.8|Cns slow virus infec NEC
C0153008|ICD9CM|PT|046.9|Unspecified slow virus infection of central nervous system
C0153008|ICD9CM|AB|046.9|Cns slow virus infec NOS
C0153012|ICD9CM|PT|048|Other enterovirus diseases of central nervous system
C0153012|ICD9CM|AB|048|Oth enteroviral cns dis
C0153013|ICD9CM|HT|049|Other non-arthropod-borne viral diseases of central nervous system
C0153014|ICD9CM|PT|049.0|Lymphocytic choriomeningitis
C0153014|ICD9CM|AB|049.0|Lymphocytic choriomening
C0153015|ICD9CM|AB|049.1|Adenoviral meningitis
C0153015|ICD9CM|PT|049.1|Meningitis due to adenovirus
C0153016|ICD9CM|HT|051|Cowpox and paravaccinia
C0153017|ICD9CM|PT|052.0|Postvaricella encephalitis
C0153017|ICD9CM|AB|052.0|Postvaricella encephalit
C0153018|ICD9CM|PT|052.1|Varicella (hemorrhagic) pneumonitis
C0153018|ICD9CM|AB|052.1|Varicella pneumonitis
C0153019|ICD9CM|PT|052.7|Chickenpox with other specified complications
C0153019|ICD9CM|AB|052.7|Varicella complicat NEC
C0153022|ICD9CM|HT|053.1|Herpes zoster with other nervous system complications
C0153022|ICD9CM|PT|053.19|Herpes zoster with other nervous system complications
C0153022|ICD9CM|AB|053.19|H zoster nerv syst NEC
C0153024|ICD9CM|PT|053.12|Postherpetic trigeminal neuralgia
C0153024|ICD9CM|AB|053.12|Postherpes trigem neural
C0153025|ICD9CM|PT|053.13|Postherpetic polyneuropathy
C0153025|ICD9CM|AB|053.13|Postherpes polyneuropath
C0153027|ICD9CM|PT|053.21|Herpes zoster keratoconjunctivitis
C0153027|ICD9CM|AB|053.21|H zoster keratoconjunct
C0153028|ICD9CM|PT|053.22|Herpes zoster iridocyclitis
C0153028|ICD9CM|AB|053.22|H zoster iridocyclitis
C0153030|ICD9CM|HT|053.7|Herpes zoster with other specified complications
C0153030|ICD9CM|PT|053.79|Herpes zoster with other specified complications
C0153030|ICD9CM|AB|053.79|H zoster complicated NEC
C0153031|ICD9CM|PT|053.71|Otitis externa due to herpes zoster
C0153031|ICD9CM|AB|053.71|H zoster otitis externa
C0153033|ICD9CM|PT|054.12|Herpetic ulceration of vulva
C0153033|ICD9CM|AB|054.12|Herpetic ulcer of vulva
C0153034|ICD9CM|PT|054.13|Herpetic infection of penis
C0153034|ICD9CM|AB|054.13|Herpetic infect of penis
C0153036|ICD9CM|HT|054.4|Herpes simplex with ophthalmic complications
C0153036|ICD9CM|PT|054.40|Herpes simplex with unspecified ophthalmic complication
C0153036|ICD9CM|AB|054.40|Herpes simplex eye NOS
C0153037|ICD9CM|PT|054.41|Herpes simplex dermatitis of eyelid
C0153037|ICD9CM|AB|054.41|Herpes simplex of eyelid
C0153038|ICD9CM|PT|054.43|Herpes simplex disciform keratitis
C0153038|ICD9CM|AB|054.43|H simplex keratitis
C0153039|ICD9CM|PT|054.44|Herpes simplex iridocyclitis
C0153039|ICD9CM|AB|054.44|H simplex iridocyclitis
C0153040|ICD9CM|PT|054.49|Herpes simplex with other ophthalmic complications
C0153040|ICD9CM|AB|054.49|Herpes simplex eye NEC
C0153041|ICD9CM|AB|054.5|Herpetic septicemia
C0153041|ICD9CM|PT|054.5|Herpetic septicemia
C0153042|ICD9CM|AB|054.6|Herpetic whitlow
C0153042|ICD9CM|PT|054.6|Herpetic whitlow
C0153043|ICD9CM|HT|054.7|Herpes simplex with other specified complications
C0153043|ICD9CM|PT|054.79|Herpes simplex with other specified complications
C0153043|ICD9CM|AB|054.79|H simplex complicat NEC
C0153045|ICD9CM|PT|054.72|Herpes simplex meningitis
C0153045|ICD9CM|AB|054.72|H simplex meningitis
C0153046|ICD9CM|PT|054.73|Herpes simplex otitis externa
C0153046|ICD9CM|AB|054.73|H simplex otitis externa
C0153047|ICD9CM|PT|054.8|Herpes simplex with unspecified complication
C0153047|ICD9CM|AB|054.8|H simplex complicat NOS
C0153048|ICD9CM|AB|055.0|Postmeasles encephalitis
C0153048|ICD9CM|PT|055.0|Postmeasles encephalitis
C0153050|ICD9CM|AB|055.2|Postmeasles otitis media
C0153050|ICD9CM|PT|055.2|Postmeasles otitis media
C0153051|ICD9CM|HT|055.7|Measles with other specified complications
C0153051|ICD9CM|PT|055.79|Measles with other specified complications
C0153051|ICD9CM|AB|055.79|Measles complication NEC
C0153052|ICD9CM|PT|055.71|Measles keratoconjunctivitis
C0153052|ICD9CM|AB|055.71|Measles keratitis
C0153053|ICD9CM|AB|055.8|Measles complication NOS
C0153053|ICD9CM|PT|055.8|Measles with unspecified complication
C0153057|ICD9CM|PT|056.09|Rubella with other neurological complications
C0153057|ICD9CM|AB|056.09|Rubella nerve compl NEC
C0153058|ICD9CM|HT|056.7|Rubella with other specified complications
C0153058|ICD9CM|PT|056.79|Rubella with other specified complications
C0153058|ICD9CM|AB|056.79|Rubella complication NEC
C0153060|ICD9CM|AB|056.8|Rubella complication NOS
C0153060|ICD9CM|PT|056.8|Rubella with unspecified complications
C0153061|ICD9CM|HT|057|Other viral exanthemata
C0153062|ICD9CM|AB|057.9|Viral exanthemata NOS
C0153062|ICD9CM|PT|057.9|Viral exanthem, unspecified
C0153064|ICD9CM|PT|062.1|Western equine encephalitis
C0153064|ICD9CM|AB|062.1|West equine encephalitis
C0153065|ICD9CM|PT|062.2|Eastern equine encephalitis
C0153065|ICD9CM|AB|062.2|East equine encephalitis
C0153066|ICD9CM|AB|062.4|Australian encephalitis
C0153066|ICD9CM|PT|062.4|Australian encephalitis
C0153069|ICD9CM|PT|064|Viral encephalitis transmitted by other and unspecified arthropods
C0153069|ICD9CM|AB|064|Vir enceph arthropod NEC
C0153070|ICD9CM|PT|065.3|Other tick-borne hemorrhagic fever
C0153070|ICD9CM|AB|065.3|Tick-borne hem fever NEC
C0153071|ICD9CM|PT|065.4|Mosquito-borne hemorrhagic fever
C0153071|ICD9CM|AB|065.4|Mosquito-borne hem fever
C0153072|ICD9CM|PT|065.8|Other specified arthropod-borne hemorrhagic fever
C0153072|ICD9CM|AB|065.8|Arthropod hem fever NEC
C0153073|ICD9CM|HT|066|Other arthropod-borne viral diseases
C0153074|ICD9CM|PT|066.8|Other specified arthropod-borne viral diseases
C0153074|ICD9CM|AB|066.8|Arthropod virus NEC
C0153075|ICD9CM|PT|070.0|Viral hepatitis A with hepatic coma
C0153075|ICD9CM|AB|070.0|Hepatitis A with coma
C0153076|ICD9CM|HT|070.2|Viral hepatitis B with hepatic coma
C0153081|ICD9CM|HT|070.4|Other specified viral hepatitis with hepatic coma
C0153081|ICD9CM|PT|070.49|Other specified viral hepatitis with hepatic coma
C0153081|ICD9CM|AB|070.49|Oth vrl hepat w hpt coma
C0153083|ICD9CM|PT|070.42|Hepatitis delta without mention of active hepatitis B disease with hepatic coma
C0153083|ICD9CM|AB|070.42|Hpt dlt wo b w hpt coma
C0153084|ICD9CM|PT|070.43|Hepatitis E with hepatic coma
C0153084|ICD9CM|AB|070.43|Hpt E w hepat Coma
C0153085|ICD9CM|HT|070.5|Other specified viral hepatitis without mention of hepatic coma
C0153085|ICD9CM|PT|070.59|Other specified viral hepatitis without mention of hepatic coma
C0153085|ICD9CM|AB|070.59|Oth vrl hpat wo hpt coma
C0153088|ICD9CM|PT|070.53|Hepatitis E without mention of hepatic coma
C0153088|ICD9CM|AB|070.53|Hpt E wo hepat Coma
C0153089|ICD9CM|PT|070.6|Unspecified viral hepatitis with hepatic coma
C0153089|ICD9CM|AB|070.6|Viral hepat NOS w coma
C0153091|ICD9CM|AB|072.0|Mumps orchitis
C0153091|ICD9CM|PT|072.0|Mumps orchitis
C0153092|ICD9CM|AB|072.1|Mumps meningitis
C0153092|ICD9CM|PT|072.1|Mumps meningitis
C0153093|ICD9CM|AB|072.2|Mumps encephalitis
C0153093|ICD9CM|PT|072.2|Mumps encephalitis
C0153094|ICD9CM|AB|072.3|Mumps pancreatitis
C0153094|ICD9CM|PT|072.3|Mumps pancreatitis
C0153095|ICD9CM|PT|072.79|Other mumps with other specified complications
C0153095|ICD9CM|HT|072.7|Mumps with other specified complications
C0153095|ICD9CM|AB|072.79|Mumps complication NEC
C0153096|ICD9CM|AB|072.71|Mumps hepatitis
C0153096|ICD9CM|PT|072.71|Mumps hepatitis
C0153097|ICD9CM|AB|072.72|Mumps polyneuropathy
C0153097|ICD9CM|PT|072.72|Mumps polyneuropathy
C0153098|ICD9CM|AB|072.8|Mumps complication NOS
C0153098|ICD9CM|PT|072.8|Mumps with unspecified complication
C0153099|ICD9CM|PT|073.0|Ornithosis with pneumonia
C0153099|ICD9CM|AB|073.0|Ornithosis pneumonia
C0153100|ICD9CM|PT|073.7|Ornithosis with other specified complications
C0153100|ICD9CM|AB|073.7|Ornithosis complicat NEC
C0153101|ICD9CM|PT|073.8|Ornithosis with unspecified complication
C0153101|ICD9CM|AB|073.8|Ornithosis complicat NOS
C0153103|ICD9CM|HT|074.2|Coxsackie carditis
C0153103|ICD9CM|AB|074.20|Coxsackie carditis NOS
C0153103|ICD9CM|PT|074.20|Coxsackie carditis, unspecified
C0153104|ICD9CM|AB|074.21|Coxsackie pericarditis
C0153104|ICD9CM|PT|074.21|Coxsackie pericarditis
C0153105|ICD9CM|AB|074.22|Coxsackie endocarditis
C0153105|ICD9CM|PT|074.22|Coxsackie endocarditis
C0153106|ICD9CM|AB|074.23|Coxsackie myocarditis
C0153106|ICD9CM|PT|074.23|Coxsackie myocarditis
C0153107|ICD9CM|AB|076.0|Trachoma, initial stage
C0153107|ICD9CM|PT|076.0|Trachoma, initial stage
C0153108|ICD9CM|AB|076.1|Trachoma, active stage
C0153108|ICD9CM|PT|076.1|Trachoma, active stage
C0153109|ICD9CM|HT|077|Other diseases of conjunctiva due to viruses and Chlamydiae
C0153110|ICD9CM|PT|077.3|Other adenoviral conjunctivitis
C0153110|ICD9CM|AB|077.3|Adenoviral conjunct NEC
C0153111|ICD9CM|HT|078|Other diseases due to viruses and Chlamydiae
C0153111|ICD9CM|HT|070-079.99|OTHER DISEASES DUE TO VIRUSES AND CHLAMYDIAE
C0153112|ICD9CM|PT|078.7|Arenaviral hemorrhagic fever
C0153112|ICD9CM|AB|078.7|Arenaviral hem fever
C0153114|ICD9CM|AB|079.99|Viral infection NOS
C0153114|ICD9CM|PT|079.99|Unspecified viral infection
C0153115|ICD9CM|PT|079.3|Rhinovirus infection in conditions classified elsewhere and of unspecified site
C0153115|ICD9CM|AB|079.3|Rhinovirus infect NOS
C0153116|ICD9CM|HT|081|Other typhus
C0153117|ICD9CM|HT|082|Tick-borne rickettsioses
C0153117|ICD9CM|PT|082.9|Tick-borne rickettsiosis, unspecified
C0153117|ICD9CM|AB|082.9|Tick-borne ricketts NOS
C0153118|ICD9CM|PT|082.8|Other specified tick-borne rickettsioses
C0153118|ICD9CM|AB|082.8|Tick-borne ricketts NEC
C0153119|ICD9CM|HT|083|Other rickettsioses
C0153120|ICD9CM|PT|083.8|Other specified rickettsioses
C0153120|ICD9CM|AB|083.8|Rickettsioses NEC
C0153121|ICD9CM|AB|084.5|Mixed malaria
C0153121|ICD9CM|PT|084.5|Mixed malaria
C0153122|ICD9CM|AB|084.7|Induced malaria
C0153122|ICD9CM|PT|084.7|Induced malaria
C0153123|ICD9CM|PT|084.9|Other pernicious complications of malaria
C0153123|ICD9CM|AB|084.9|Malaria complicated NEC
C0153125|ICD9CM|PT|086.1|Chagas' disease with other organ involvement
C0153125|ICD9CM|AB|086.1|Chagas dis of oth organ
C0153126|ICD9CM|HT|088|Other arthropod-borne diseases
C0153129|ICD9CM|PT|090.1|Early congenital syphilis, latent
C0153129|ICD9CM|AB|090.1|Early congen syph latent
C0153132|ICD9CM|HT|090.4|Juvenile neurosyphilis
C0153132|ICD9CM|PT|090.40|Juvenile neurosyphilis, unspecified
C0153132|ICD9CM|AB|090.40|Juvenile neurosyph NOS
C0153133|ICD9CM|PT|090.41|Congenital syphilitic encephalitis
C0153133|ICD9CM|AB|090.41|Congen syph encephalitis
C0153134|ICD9CM|PT|090.42|Congenital syphilitic meningitis
C0153134|ICD9CM|AB|090.42|Congen syph meningitis
C0153135|ICD9CM|PT|090.49|Other juvenile neurosyphilis
C0153135|ICD9CM|AB|090.49|Juvenile neurosyph NEC
C0153136|ICD9CM|PT|090.5|Other late congenital syphilis, symptomatic
C0153136|ICD9CM|AB|090.5|Late congen syph symptom
C0153139|ICD9CM|HT|091|Early syphilis, symptomatic
C0153140|ICD9CM|AB|091.1|Primary anal syphilis
C0153140|ICD9CM|PT|091.1|Primary anal syphilis
C0153141|ICD9CM|PT|091.2|Other primary syphilis
C0153141|ICD9CM|AB|091.2|Primary syphilis NEC
C0153145|ICD9CM|PT|091.51|Syphilitic chorioretinitis (secondary)
C0153145|ICD9CM|AB|091.51|Syphilit chorioretinitis
C0153146|ICD9CM|PT|091.52|Syphilitic iridocyclitis (secondary)
C0153146|ICD9CM|AB|091.52|Syphilitic iridocyclitis
C0153148|ICD9CM|PT|091.61|Secondary syphilitic periostitis
C0153148|ICD9CM|AB|091.61|Syphilitic periostitis
C0153149|ICD9CM|PT|091.62|Secondary syphilitic hepatitis
C0153149|ICD9CM|AB|091.62|Syphilitic hepatitis
C0153150|ICD9CM|PT|091.69|Secondary syphilis of other viscera
C0153150|ICD9CM|AB|091.69|Second syph viscera NEC
C0153151|ICD9CM|PT|091.7|Secondary syphilis, relapse
C0153151|ICD9CM|AB|091.7|Second syphilis relapse
C0153156|ICD9CM|PT|092.0|Early syphilis, latent, serological relapse after treatment
C0153156|ICD9CM|AB|092.0|Early syph latent relaps
C0153158|ICD9CM|HT|093.2|Syphilitic endocarditis
C0153160|ICD9CM|PT|093.21|Syphilitic endocarditis of mitral valve
C0153160|ICD9CM|AB|093.21|Syphilitic mitral valve
C0153161|ICD9CM|PT|093.22|Syphilitic endocarditis of aortic valve
C0153161|ICD9CM|AB|093.22|Syphilitic aortic valve
C0153162|ICD9CM|PT|093.23|Syphilitic endocarditis of tricuspid valve
C0153162|ICD9CM|AB|093.23|Syphil tricuspid valve
C0153163|ICD9CM|PT|093.24|Syphilitic endocarditis of pulmonary valve
C0153163|ICD9CM|AB|093.24|Syphil pulmonary valve
C0153164|ICD9CM|AB|093.81|Syphilitic pericarditis
C0153164|ICD9CM|PT|093.81|Syphilitic pericarditis
C0153165|ICD9CM|AB|093.82|Syphilitic myocarditis
C0153165|ICD9CM|PT|093.82|Syphilitic myocarditis
C0153166|ICD9CM|AB|094.2|Syphilitic meningitis
C0153166|ICD9CM|PT|094.2|Syphilitic meningitis
C0153167|ICD9CM|PT|094.3|Asymptomatic neurosyphilis
C0153167|ICD9CM|AB|094.3|Asymptomat neurosyphilis
C0153168|ICD9CM|AB|094.81|Syphilitic encephalitis
C0153168|ICD9CM|PT|094.81|Syphilitic encephalitis
C0153169|ICD9CM|AB|094.82|Syphilitic parkinsonism
C0153169|ICD9CM|PT|094.82|Syphilitic parkinsonism
C0153170|ICD9CM|PT|094.83|Syphilitic disseminated retinochoroiditis
C0153170|ICD9CM|AB|094.83|Syph dissem retinitis
C0153171|ICD9CM|AB|094.84|Syphilitic optic atrophy
C0153171|ICD9CM|PT|094.84|Syphilitic optic atrophy
C0153172|ICD9CM|PT|094.85|Syphilitic retrobulbar neuritis
C0153172|ICD9CM|AB|094.85|Syph retrobulb neuritis
C0153173|ICD9CM|PT|094.86|Syphilitic acoustic neuritis
C0153173|ICD9CM|AB|094.86|Syphil acoustic neuritis
C0153174|ICD9CM|PT|094.87|Syphilitic ruptured cerebral aneurysm
C0153174|ICD9CM|AB|094.87|Syph rupt cereb aneurysm
C0153176|ICD9CM|AB|095.0|Syphilitic episcleritis
C0153176|ICD9CM|PT|095.0|Syphilitic episcleritis
C0153177|ICD9CM|AB|095.1|Syphilis of lung
C0153177|ICD9CM|PT|095.1|Syphilis of lung
C0153178|ICD9CM|AB|095.2|Syphilitic peritonitis
C0153178|ICD9CM|PT|095.2|Syphilitic peritonitis
C0153179|ICD9CM|AB|095.3|Syphilis of liver
C0153179|ICD9CM|PT|095.3|Syphilis of liver
C0153180|ICD9CM|AB|095.4|Syphilis of kidney
C0153180|ICD9CM|PT|095.4|Syphilis of kidney
C0153181|ICD9CM|AB|095.5|Syphilis of bone
C0153181|ICD9CM|PT|095.5|Syphilis of bone
C0153182|ICD9CM|AB|095.6|Syphilis of muscle
C0153182|ICD9CM|PT|095.6|Syphilis of muscle
C0153183|ICD9CM|PT|095.7|Syphilis of synovium, tendon, and bursa
C0153183|ICD9CM|AB|095.7|Syphilis of tendon/bursa
C0153185|ICD9CM|PT|095.9|Late symptomatic syphilis, unspecified
C0153185|ICD9CM|AB|095.9|Late sympt syphilis NOS
C0153188|ICD9CM|AB|097.0|Late syphilis NOS
C0153188|ICD9CM|PT|097.0|Late syphilis, unspecified
C0153191|ICD9CM|PT|098.11|Gonococcal cystitis (acute)
C0153191|ICD9CM|AB|098.11|Gc cystitis (acute)
C0153192|ICD9CM|PT|098.12|Gonococcal prostatitis (acute)
C0153192|ICD9CM|AB|098.12|Gc prostatitis (acute)
C0153193|ICD9CM|PT|098.13|Gonococcal epididymo-orchitis (acute)
C0153193|ICD9CM|AB|098.13|Gc orchitis (acute)
C0153194|ICD9CM|PT|098.14|Gonococcal seminal vesiculitis (acute)
C0153194|ICD9CM|AB|098.14|Gc sem vesiculit (acute)
C0153195|ICD9CM|PT|098.15|Gonococcal cervicitis (acute)
C0153195|ICD9CM|AB|098.15|Gc cervicitis (acute)
C0153196|ICD9CM|PT|098.16|Gonococcal endometritis (acute)
C0153196|ICD9CM|AB|098.16|Gc endometritis (acute)
C0153198|ICD9CM|PT|098.19|Other gonococcal infection (acute) of upper genitourinary tract
C0153198|ICD9CM|AB|098.19|Gc (acute) upper gu NEC
C0153199|ICD9CM|PT|098.2|Gonococcal infection, chronic, of lower genitourinary tract
C0153199|ICD9CM|AB|098.2|Chr gc infect lower gu
C0153202|ICD9CM|PT|098.31|Gonococcal cystitis, chronic
C0153202|ICD9CM|AB|098.31|Gc cystitis, chronic
C0153203|ICD9CM|PT|098.32|Gonococcal prostatitis, chronic
C0153203|ICD9CM|AB|098.32|Gc prostatitis, chronic
C0153204|ICD9CM|PT|098.33|Gonococcal epididymo-orchitis, chronic
C0153204|ICD9CM|AB|098.33|Gc orchitis, chronic
C0153205|ICD9CM|PT|098.34|Gonococcal seminal vesiculitis, chronic
C0153205|ICD9CM|AB|098.34|Gc sem vesiculitis, chr
C0153206|ICD9CM|PT|098.35|Gonococcal cervicitis, chronic
C0153206|ICD9CM|AB|098.35|Gc cervicitis, chronic
C0153207|ICD9CM|PT|098.36|Gonococcal endometritis, chronic
C0153207|ICD9CM|AB|098.36|Gc endometritis, chronic
C0153208|ICD9CM|PT|098.37|Gonococcal salpingitis (chronic)
C0153208|ICD9CM|AB|098.37|Gc salpingitis (chronic)
C0153209|ICD9CM|PT|098.39|Other chronic gonococcal infection of upper genitourinary tract
C0153209|ICD9CM|AB|098.39|Chr gc upper gu NEC
C0153210|ICD9CM|HT|098.4|Gonococcal infection of eye
C0153212|ICD9CM|AB|098.41|Gonococcal iridocyclitis
C0153212|ICD9CM|PT|098.41|Gonococcal iridocyclitis
C0153213|ICD9CM|AB|098.42|Gonococcal endophthalmia
C0153213|ICD9CM|PT|098.42|Gonococcal endophthalmia
C0153214|ICD9CM|AB|098.43|Gonococcal keratitis
C0153214|ICD9CM|PT|098.43|Gonococcal keratitis
C0153215|ICD9CM|PT|098.49|Other gonococcal infection of eye
C0153215|ICD9CM|AB|098.49|Gonococcal eye NEC
C0153216|ICD9CM|HT|098.5|Gonococcal infection of joint
C0153216|ICD9CM|AB|098.50|Gonococcal arthritis
C0153216|ICD9CM|PT|098.50|Gonococcal arthritis
C0153218|ICD9CM|AB|098.52|Gonococcal bursitis
C0153218|ICD9CM|PT|098.52|Gonococcal bursitis
C0153219|ICD9CM|AB|098.53|Gonococcal spondylitis
C0153219|ICD9CM|PT|098.53|Gonococcal spondylitis
C0153220|ICD9CM|PT|098.59|Other gonococcal infection of joint
C0153220|ICD9CM|AB|098.59|Gc infect joint NEC
C0153222|ICD9CM|PT|098.7|Gonococcal infection of anus and rectum
C0153222|ICD9CM|AB|098.7|Gc infect anus & rectum
C0153223|ICD9CM|HT|098.8|Gonococcal infection of other specified sites
C0153223|ICD9CM|PT|098.89|Gonococcal infection of other specified sites
C0153223|ICD9CM|AB|098.89|Gonococcal inf site NEC
C0153225|ICD9CM|AB|098.82|Gonococcal meningitis
C0153225|ICD9CM|PT|098.82|Gonococcal meningitis
C0153226|ICD9CM|AB|098.83|Gonococcal pericarditis
C0153226|ICD9CM|PT|098.83|Gonococcal pericarditis
C0153227|ICD9CM|AB|098.84|Gonococcal endocarditis
C0153227|ICD9CM|PT|098.84|Gonococcal endocarditis
C0153228|ICD9CM|PT|098.85|Other gonococcal heart disease
C0153228|ICD9CM|AB|098.85|Gonococcal heart dis NEC
C0153229|ICD9CM|HT|099|Other venereal diseases
C0153231|ICD9CM|HT|100.8|Other specified leptospiral infections
C0153231|ICD9CM|PT|100.89|Other specified leptospiral infections
C0153231|ICD9CM|AB|100.89|Leptospiral infect NEC
C0153232|ICD9CM|AB|100.81|Leptospiral meningitis
C0153232|ICD9CM|PT|100.81|Leptospiral meningitis (aseptic)
C0153234|ICD9CM|PT|102.1|Multiple papillomata due to yaws and wet crab yaws
C0153234|ICD9CM|AB|102.1|Multiple papillomata
C0153235|ICD9CM|PT|102.2|Other early skin lesions of yaws
C0153235|ICD9CM|AB|102.2|Early skin yaws NEC
C0153239|ICD9CM|PT|102.7|Other manifestations of yaws
C0153239|ICD9CM|AB|102.7|Yaws manifestations NEC
C0153240|ICD9CM|AB|102.8|Latent yaws
C0153240|ICD9CM|PT|102.8|Latent yaws
C0153241|ICD9CM|PT|103.0|Primary lesions of pinta
C0153241|ICD9CM|AB|103.0|Pinta primary lesions
C0153242|ICD9CM|PT|103.1|Intermediate lesions of pinta
C0153242|ICD9CM|AB|103.1|Pinta intermed lesions
C0153243|ICD9CM|PT|103.2|Late lesions of pinta
C0153243|ICD9CM|AB|103.2|Pinta late lesions
C0153244|ICD9CM|PT|103.3|Mixed lesions of pinta
C0153244|ICD9CM|AB|103.3|Pinta mixed lesions
C0153245|ICD9CM|HT|104|Other spirochetal infection
C0153246|ICD9CM|AB|110.2|Dermatophytosis of hand
C0153246|ICD9CM|PT|110.2|Dermatophytosis of hand
C0153248|ICD9CM|PT|110.8|Dermatophytosis of other specified sites
C0153248|ICD9CM|AB|110.8|Dermatophytosis site NEC
C0153249|ICD9CM|AB|111.3|Black piedra
C0153249|ICD9CM|PT|111.3|Black piedra
C0153250|ICD9CM|PT|112.2|Candidiasis of other urogenital sites
C0153250|ICD9CM|AB|112.2|Candidias urogenital NEC
C0153251|ICD9CM|AB|112.4|Candidiasis of lung
C0153251|ICD9CM|PT|112.4|Candidiasis of lung
C0153252|ICD9CM|AB|112.5|Disseminated candidiasis
C0153252|ICD9CM|PT|112.5|Disseminated candidiasis
C0153253|ICD9CM|HT|112.8|Candidiasis of other specified sites
C0153254|ICD9CM|AB|112.81|Candidal endocarditis
C0153254|ICD9CM|PT|112.81|Candidal endocarditis
C0153255|ICD9CM|AB|112.82|Candidal otitis externa
C0153255|ICD9CM|PT|112.82|Candidal otitis externa
C0153256|ICD9CM|AB|112.83|Candidal meningitis
C0153256|ICD9CM|PT|112.83|Candidal meningitis
C0153257|ICD9CM|PT|114.0|Primary coccidioidomycosis (pulmonary)
C0153257|ICD9CM|AB|114.0|Primary coccidioidomycos
C0153259|ICD9CM|AB|114.2|Coccidioidal meningitis
C0153259|ICD9CM|PT|114.2|Coccidioidal meningitis
C0153261|ICD9CM|HT|115.0|Infection by Histoplasma capsulatum
C0153262|ICD9CM|PT|115.00|Infection by Histoplasma capsulatum, without mention of manifestation
C0153262|ICD9CM|AB|115.00|Histoplasma capsulat NOS
C0153263|ICD9CM|PT|115.01|Infection by Histoplasma capsulatum, meningitis
C0153263|ICD9CM|AB|115.01|Histoplasm capsul mening
C0153264|ICD9CM|PT|115.02|Infection by Histoplasma capsulatum, retinitis
C0153264|ICD9CM|AB|115.02|Histoplasm capsul retina
C0153265|ICD9CM|PT|115.03|Infection by Histoplasma capsulatum, pericarditis
C0153265|ICD9CM|AB|115.03|Histoplasm caps pericard
C0153266|ICD9CM|PT|115.04|Infection by Histoplasma capsulatum, endocarditis
C0153266|ICD9CM|PT|115.94|Histoplasmosis, unspecified, endocarditis
C0153266|ICD9CM|AB|115.04|Histoplasm caps endocard
C0153266|ICD9CM|AB|115.94|Histoplasmosis endocard
C0153268|ICD9CM|PT|115.09|Infection by Histoplasma capsulatum, other
C0153268|ICD9CM|AB|115.09|Histoplasma capsulat NEC
C0153270|ICD9CM|PT|115.10|Infection by Histoplasma duboisii, without mention of manifestation
C0153270|ICD9CM|AB|115.10|Histoplasma duboisii NOS
C0153271|ICD9CM|PT|115.11|Infection by Histoplasma duboisii, meningitis
C0153271|ICD9CM|AB|115.11|Histoplasm dubois mening
C0153272|ICD9CM|PT|115.12|Infection by Histoplasma duboisii, retinitis
C0153272|ICD9CM|AB|115.12|Histoplasm dubois retina
C0153273|ICD9CM|PT|115.13|Infection by Histoplasma duboisii, pericarditis
C0153273|ICD9CM|AB|115.13|Histoplasm dub pericard
C0153274|ICD9CM|PT|115.14|Infection by Histoplasma duboisii, endocarditis
C0153274|ICD9CM|AB|115.14|Histoplasm dub endocard
C0153275|ICD9CM|PT|115.15|Infection by Histoplasma duboisii, pneumonia
C0153275|ICD9CM|AB|115.15|Histoplasm dub pneumonia
C0153276|ICD9CM|PT|115.19|Infection by Histoplasma duboisii, other
C0153276|ICD9CM|AB|115.19|Histoplasma duboisii NEC
C0153277|ICD9CM|PT|115.91|Histoplasmosis, unspecified, meningitis
C0153277|ICD9CM|AB|115.91|Histoplasmosis meningit
C0153278|ICD9CM|AB|115.92|Histoplasmosis retinitis
C0153278|ICD9CM|PT|115.92|Histoplasmosis, unspecified, retinitis
C0153279|ICD9CM|PT|115.93|Histoplasmosis, unspecified, pericarditis
C0153279|ICD9CM|AB|115.93|Histoplasmosis pericard
C0153281|ICD9CM|AB|115.95|Histoplasmosis pneumonia
C0153281|ICD9CM|PT|115.95|Histoplasmosis, unspecified, pneumonia
C0153285|ICD9CM|AB|117.6|Allescheriosis
C0153285|ICD9CM|PT|117.6|Allescheriosis [Petriellidosis]
C0153288|ICD9CM|HT|121|Other trematode infections
C0153289|ICD9CM|PT|122.0|Echinococcus granulosus infection of liver
C0153289|ICD9CM|AB|122.0|Echinococc granul liver
C0153290|ICD9CM|PT|122.1|Echinococcus granulosus infection of lung
C0153290|ICD9CM|AB|122.1|Echinococc granul lung
C0153291|ICD9CM|PT|122.2|Echinococcus granulosus infection of thyroid
C0153291|ICD9CM|AB|122.2|Echinococc gran thyroid
C0153292|ICD9CM|PT|122.3|Echinococcus granulosus infection, other
C0153292|ICD9CM|AB|122.3|Echinococc granul NEC
C0153293|ICD9CM|PT|122.5|Echinococcus multilocularis infection of liver
C0153293|ICD9CM|AB|122.5|Echinococ multiloc liver
C0153296|ICD9CM|HT|123|Other cestode infection
C0153298|ICD9CM|HT|125|Filarial infection and dracontiasis
C0153299|ICD9CM|AB|126.2|Ancylostoma braziliense
C0153299|ICD9CM|PT|126.2|Ancylostomiasis due to ancylostoma braziliense
C0153302|ICD9CM|HT|127|Other intestinal helminthiases
C0153303|ICD9CM|PT|127.8|Mixed intestinal helminthiasis
C0153303|ICD9CM|AB|127.8|Mixed intestine helminth
C0153307|ICD9CM|PT|130.1|Conjunctivitis due to toxoplasmosis
C0153307|ICD9CM|AB|130.1|Toxoplasm conjunctivitis
C0153308|ICD9CM|PT|130.2|Chorioretinitis due to toxoplasmosis
C0153308|ICD9CM|AB|130.2|Toxoplasm chorioretinit
C0153312|ICD9CM|PT|130.7|Toxoplasmosis of other specified sites
C0153312|ICD9CM|AB|130.7|Toxoplasmosis site NEC
C0153314|ICD9CM|AB|131.02|Trichomonal urethritis
C0153314|ICD9CM|PT|131.02|Trichomonal urethritis
C0153315|ICD9CM|AB|131.03|Trichomonal prostatitis
C0153315|ICD9CM|PT|131.03|Trichomonal prostatitis
C0153316|ICD9CM|PT|131.09|Other urogenital trichomoniasis
C0153316|ICD9CM|AB|131.09|Urogenital trichomon NEC
C0153317|ICD9CM|HT|132|Pediculosis and phthirus infestation
C0153322|ICD9CM|HT|134|Other infestation
C0153323|ICD9CM|PT|134.1|Other arthropod infestation
C0153323|ICD9CM|AB|134.1|Arthropod infest NEC
C0153324|ICD9CM|PT|134.8|Other specified infestations
C0153324|ICD9CM|AB|134.8|Infestation NEC
C0153325|ICD9CM|HT|136|Other and unspecified infectious and parasitic diseases
C0153325|ICD9CM|HT|130-136.99|OTHER INFECTIOUS AND PARASITIC DISEASES
C0153326|ICD9CM|HT|136.2|Specific infections by free-living amebae
C0153327|ICD9CM|AB|136.4|Psorospermiasis
C0153327|ICD9CM|PT|136.4|Psorospermiasis
C0153328|ICD9CM|PT|136.8|Other specified infectious and parasitic diseases
C0153328|ICD9CM|AB|136.8|Infect/parasite dis NEC
C0153329|ICD9CM|HT|137|Late effects of tuberculosis
C0153331|ICD9CM|PT|137.1|Late effects of central nervous system tuberculosis
C0153331|ICD9CM|AB|137.1|Late effect cns TB
C0153333|ICD9CM|PT|137.3|Late effects of tuberculosis of bones and joints
C0153333|ICD9CM|AB|137.3|Late eff bone & joint TB
C0153334|ICD9CM|PT|137.4|Late effects of tuberculosis of other specified organs
C0153334|ICD9CM|AB|137.4|Late effect TB NEC
C0153336|ICD9CM|HT|139|Late effects of other infectious and parasitic diseases
C0153336|ICD9CM|PT|139.8|Late effects of other and unspecified infectious and parasitic diseases
C0153336|ICD9CM|AB|139.8|Late eff infect dis NEC
C0153337|ICD9CM|PT|139.0|Late effects of viral encephalitis
C0153337|ICD9CM|AB|139.0|Late eff viral encephal
C0153338|ICD9CM|PT|139.1|Late effects of trachoma
C0153338|ICD9CM|AB|139.1|Late effect of trachoma
C0153340|ICD9CM|HT|140|Malignant neoplasm of lip
C0153346|ICD9CM|PT|140.6|Malignant neoplasm of commissure of lip
C0153346|ICD9CM|AB|140.6|Mal neo lip, commissure
C0153347|ICD9CM|PT|140.8|Malignant neoplasm of other sites of lip
C0153347|ICD9CM|AB|140.8|Mal neo lip NEC
C0153349|ICD9CM|HT|141|Malignant neoplasm of tongue
C0153349|ICD9CM|PT|141.9|Malignant neoplasm of tongue, unspecified
C0153349|ICD9CM|AB|141.9|Malig neo tongue NOS
C0153350|ICD9CM|PT|141.0|Malignant neoplasm of base of tongue
C0153350|ICD9CM|AB|141.0|Mal neo tongue base
C0153351|ICD9CM|PT|141.1|Malignant neoplasm of dorsal surface of tongue
C0153351|ICD9CM|AB|141.1|Mal neo dorsal tongue
C0153354|ICD9CM|PT|141.4|Malignant neoplasm of anterior two-thirds of tongue, part unspecified
C0153354|ICD9CM|AB|141.4|Mal neo ant 2/3 tongue
C0153356|ICD9CM|PT|141.6|Malignant neoplasm of lingual tonsil
C0153356|ICD9CM|AB|141.6|Mal neo lingual tonsil
C0153357|ICD9CM|PT|141.8|Malignant neoplasm of other sites of tongue
C0153357|ICD9CM|AB|141.8|Malig neo tongue NEC
C0153360|ICD9CM|PT|142.1|Malignant neoplasm of submandibular gland
C0153360|ICD9CM|AB|142.1|Malig neo submandibular
C0153361|ICD9CM|PT|142.2|Malignant neoplasm of sublingual gland
C0153361|ICD9CM|AB|142.2|Malig neo sublingual
C0153362|ICD9CM|PT|142.8|Malignant neoplasm of other major salivary glands
C0153362|ICD9CM|AB|142.8|Mal neo maj salivary NEC
C0153364|ICD9CM|HT|143|Malignant neoplasm of gum
C0153364|ICD9CM|PT|143.9|Malignant neoplasm of gum, unspecified
C0153364|ICD9CM|AB|143.9|Malig neo gum NOS
C0153365|ICD9CM|PT|143.0|Malignant neoplasm of upper gum
C0153365|ICD9CM|AB|143.0|Malig neo upper gum
C0153367|ICD9CM|PT|143.8|Malignant neoplasm of other sites of gum
C0153367|ICD9CM|AB|143.8|Malig neo gum NEC
C0153368|ICD9CM|HT|144|Malignant neoplasm of floor of mouth
C0153368|ICD9CM|PT|144.9|Malignant neoplasm of floor of mouth, part unspecified
C0153368|ICD9CM|AB|144.9|Mal neo mouth floor NOS
C0153369|ICD9CM|PT|144.0|Malignant neoplasm of anterior portion of floor of mouth
C0153369|ICD9CM|AB|144.0|Mal neo ant floor mouth
C0153371|ICD9CM|PT|144.8|Malignant neoplasm of other sites of floor of mouth
C0153371|ICD9CM|AB|144.8|Mal neo mouth floor NEC
C0153372|ICD9CM|HT|145|Malignant neoplasm of other and unspecified parts of mouth
C0153373|ICD9CM|PT|145.0|Malignant neoplasm of cheek mucosa
C0153373|ICD9CM|AB|145.0|Mal neo cheek mucosa
C0153374|ICD9CM|PT|145.1|Malignant neoplasm of vestibule of mouth
C0153374|ICD9CM|AB|145.1|Mal neo mouth vestibule
C0153375|ICD9CM|PT|145.2|Malignant neoplasm of hard palate
C0153375|ICD9CM|AB|145.2|Malig neo hard palate
C0153376|ICD9CM|PT|145.3|Malignant neoplasm of soft palate
C0153376|ICD9CM|AB|145.3|Malig neo soft palate
C0153377|ICD9CM|PT|145.4|Malignant neoplasm of uvula
C0153377|ICD9CM|AB|145.4|Malignant neoplasm uvula
C0153378|ICD9CM|PT|145.5|Malignant neoplasm of palate, unspecified
C0153378|ICD9CM|AB|145.5|Malignant neo palate NOS
C0153379|ICD9CM|PT|145.6|Malignant neoplasm of retromolar area
C0153379|ICD9CM|AB|145.6|Malig neo retromolar
C0153380|ICD9CM|PT|145.8|Malignant neoplasm of other specified parts of mouth
C0153380|ICD9CM|AB|145.8|Malig neoplasm mouth NEC
C0153381|ICD9CM|PT|145.9|Malignant neoplasm of mouth, unspecified
C0153381|ICD9CM|AB|145.9|Malig neoplasm mouth NOS
C0153382|ICD9CM|HT|146|Malignant neoplasm of oropharynx
C0153382|ICD9CM|PT|146.9|Malignant neoplasm of oropharynx, unspecified site
C0153382|ICD9CM|AB|146.9|Malig neo oropharynx NOS
C0153384|ICD9CM|PT|146.1|Malignant neoplasm of tonsillar fossa
C0153384|ICD9CM|AB|146.1|Mal neo tonsillar fossa
C0153385|ICD9CM|PT|146.2|Malignant neoplasm of tonsillar pillars (anterior) (posterior)
C0153385|ICD9CM|AB|146.2|Mal neo tonsil pillars
C0153386|ICD9CM|PT|146.3|Malignant neoplasm of vallecula epiglottica
C0153386|ICD9CM|AB|146.3|Malign neopl vallecula
C0153388|ICD9CM|PT|146.5|Malignant neoplasm of junctional region of oropharynx
C0153388|ICD9CM|AB|146.5|Mal neo epiglottis junct
C0153389|ICD9CM|PT|146.6|Malignant neoplasm of lateral wall of oropharynx
C0153389|ICD9CM|AB|146.6|Mal neo lat oropharynx
C0153390|ICD9CM|PT|146.7|Malignant neoplasm of posterior wall of oropharynx
C0153390|ICD9CM|AB|146.7|Mal neo post oropharynx
C0153391|ICD9CM|PT|146.8|Malignant neoplasm of other specified sites of oropharynx
C0153391|ICD9CM|AB|146.8|Mal neo oropharynx NEC
C0153392|ICD9CM|HT|147|Malignant neoplasm of nasopharynx
C0153392|ICD9CM|PT|147.9|Malignant neoplasm of nasopharynx, unspecified site
C0153392|ICD9CM|AB|147.9|Mal neo nasopharynx NOS
C0153393|ICD9CM|PT|147.0|Malignant neoplasm of superior wall of nasopharynx
C0153393|ICD9CM|AB|147.0|Mal neo super nasopharyn
C0153394|ICD9CM|PT|147.1|Malignant neoplasm of posterior wall of nasopharynx
C0153394|ICD9CM|AB|147.1|Mal neo post nasopharynx
C0153395|ICD9CM|PT|147.2|Malignant neoplasm of lateral wall of nasopharynx
C0153395|ICD9CM|AB|147.2|Mal neo lat nasopharynx
C0153396|ICD9CM|PT|147.3|Malignant neoplasm of anterior wall of nasopharynx
C0153396|ICD9CM|AB|147.3|Mal neo ant nasopharynx
C0153397|ICD9CM|PT|147.8|Malignant neoplasm of other specified sites of nasopharynx
C0153397|ICD9CM|AB|147.8|Mal neo nasopharynx NEC
C0153398|ICD9CM|HT|148|Malignant neoplasm of hypopharynx
C0153398|ICD9CM|PT|148.9|Malignant neoplasm of hypopharynx, unspecified site
C0153398|ICD9CM|AB|148.9|Mal neo hypopharynx NOS
C0153400|ICD9CM|PT|148.1|Malignant neoplasm of pyriform sinus
C0153400|ICD9CM|AB|148.1|Mal neo pyriform sinus
C0153401|ICD9CM|PT|148.2|Malignant neoplasm of aryepiglottic fold, hypopharyngeal aspect
C0153401|ICD9CM|AB|148.2|Mal neo aryepiglott fold
C0153403|ICD9CM|PT|148.8|Malignant neoplasm of other specified sites of hypopharynx
C0153403|ICD9CM|AB|148.8|Mal neo hypopharynx NEC
C0153404|ICD9CM|HT|149|Malignant neoplasm of other and ill-defined sites within the lip, oral cavity, and pharynx
C0153405|ICD9CM|PT|149.0|Malignant neoplasm of pharynx, unspecified
C0153405|ICD9CM|AB|149.0|Mal neo pharynx NOS
C0153406|ICD9CM|PT|149.1|Malignant neoplasm of waldeyer's ring
C0153406|ICD9CM|AB|149.1|Mal neo waldeyer's ring
C0153407|ICD9CM|PT|149.8|Malignant neoplasm of other sites within the lip and oral cavity
C0153407|ICD9CM|AB|149.8|Mal neo oral/pharynx NEC
C0153408|ICD9CM|PT|149.9|Malignant neoplasm of ill-defined sites within the lip and oral cavity
C0153408|ICD9CM|AB|149.9|Mal neo orophryn ill-def
C0153411|ICD9CM|PT|150.1|Malignant neoplasm of thoracic esophagus
C0153411|ICD9CM|AB|150.1|Mal neo thoracic esophag
C0153413|ICD9CM|PT|150.3|Malignant neoplasm of upper third of esophagus
C0153413|ICD9CM|AB|150.3|Mal neo upper 3rd esoph
C0153414|ICD9CM|PT|150.4|Malignant neoplasm of middle third of esophagus
C0153414|ICD9CM|AB|150.4|Mal neo middle 3rd esoph
C0153415|ICD9CM|PT|150.5|Malignant neoplasm of lower third of esophagus
C0153415|ICD9CM|AB|150.5|Mal neo lower 3rd esoph
C0153416|ICD9CM|PT|150.8|Malignant neoplasm of other specified part of esophagus
C0153416|ICD9CM|AB|150.8|Mal neo esophagus NEC
C0153417|ICD9CM|PT|151.0|Malignant neoplasm of cardia
C0153417|ICD9CM|AB|151.0|Mal neo stomach cardia
C0153418|ICD9CM|PT|151.1|Malignant neoplasm of pylorus
C0153418|ICD9CM|AB|151.1|Malignant neo pylorus
C0153419|ICD9CM|PT|151.2|Malignant neoplasm of pyloric antrum
C0153419|ICD9CM|AB|151.2|Mal neo pyloric antrum
C0153420|ICD9CM|PT|151.3|Malignant neoplasm of fundus of stomach
C0153420|ICD9CM|AB|151.3|Mal neo stomach fundus
C0153421|ICD9CM|PT|151.4|Malignant neoplasm of body of stomach
C0153421|ICD9CM|AB|151.4|Mal neo stomach body
C0153422|ICD9CM|PT|151.5|Malignant neoplasm of lesser curvature of stomach, unspecified
C0153422|ICD9CM|AB|151.5|Mal neo stom lesser curv
C0153423|ICD9CM|PT|151.6|Malignant neoplasm of greater curvature of stomach, unspecified
C0153423|ICD9CM|AB|151.6|Mal neo stom great curv
C0153424|ICD9CM|PT|151.8|Malignant neoplasm of other specified sites of stomach
C0153424|ICD9CM|AB|151.8|Malig neopl stomach NEC
C0153425|ICD9CM|PT|152.9|Malignant neoplasm of small intestine, unspecified site
C0153425|ICD9CM|AB|152.9|Mal neo small bowel NOS
C0153426|ICD9CM|PT|152.0|Malignant neoplasm of duodenum
C0153426|ICD9CM|AB|152.0|Malignant neopl duodenum
C0153427|ICD9CM|PT|152.1|Malignant neoplasm of jejunum
C0153427|ICD9CM|AB|152.1|Malignant neopl jejunum
C0153428|ICD9CM|PT|152.2|Malignant neoplasm of ileum
C0153428|ICD9CM|AB|152.2|Malignant neoplasm ileum
C0153429|ICD9CM|PT|152.3|Malignant neoplasm of Meckel's diverticulum
C0153429|ICD9CM|AB|152.3|Mal neo meckel's divert
C0153430|ICD9CM|PT|152.8|Malignant neoplasm of other specified sites of small intestine
C0153430|ICD9CM|AB|152.8|Mal neo small bowel NEC
C0153433|ICD9CM|PT|153.0|Malignant neoplasm of hepatic flexure
C0153433|ICD9CM|AB|153.0|Mal neo hepatic flexure
C0153434|ICD9CM|PT|153.1|Malignant neoplasm of transverse colon
C0153434|ICD9CM|AB|153.1|Mal neo transverse colon
C0153435|ICD9CM|PT|153.2|Malignant neoplasm of descending colon
C0153435|ICD9CM|AB|153.2|Mal neo descend colon
C0153436|ICD9CM|PT|153.3|Malignant neoplasm of sigmoid colon
C0153436|ICD9CM|AB|153.3|Mal neo sigmoid colon
C0153437|ICD9CM|PT|153.4|Malignant neoplasm of cecum
C0153437|ICD9CM|AB|153.4|Malignant neoplasm cecum
C0153439|ICD9CM|PT|153.6|Malignant neoplasm of ascending colon
C0153439|ICD9CM|AB|153.6|Malig neo ascend colon
C0153440|ICD9CM|PT|153.7|Malignant neoplasm of splenic flexure
C0153440|ICD9CM|AB|153.7|Mal neo splenic flexure
C0153441|ICD9CM|PT|153.8|Malignant neoplasm of other specified sites of large intestine
C0153441|ICD9CM|AB|153.8|Malignant neo colon NEC
C0153442|ICD9CM|HT|154|Malignant neoplasm of rectum, rectosigmoid junction, and anus
C0153443|ICD9CM|PT|154.0|Malignant neoplasm of rectosigmoid junction
C0153443|ICD9CM|AB|154.0|Mal neo rectosigmoid jct
C0153445|ICD9CM|PT|154.2|Malignant neoplasm of anal canal
C0153445|ICD9CM|AB|154.2|Malig neopl anal canal
C0153446|ICD9CM|PT|154.3|Malignant neoplasm of anus, unspecified site
C0153446|ICD9CM|AB|154.3|Malignant neo anus NOS
C0153447|ICD9CM|PT|154.8|Malignant neoplasm of other sites of rectum, rectosigmoid junction, and anus
C0153447|ICD9CM|AB|154.8|Mal neo rectum/anus NEC
C0153448|ICD9CM|HT|155|Malignant neoplasm of liver and intrahepatic bile ducts
C0153452|ICD9CM|PT|156.0|Malignant neoplasm of gallbladder
C0153452|ICD9CM|AB|156.0|Malig neo gallbladder
C0153453|ICD9CM|PT|156.1|Malignant neoplasm of extrahepatic bile ducts
C0153453|ICD9CM|AB|156.1|Mal neo extrahepat ducts
C0153454|ICD9CM|PT|156.2|Malignant neoplasm of ampulla of vater
C0153454|ICD9CM|AB|156.2|Mal neo ampulla of vater
C0153455|ICD9CM|PT|156.8|Malignant neoplasm of other specified sites of gallbladder and extrahepatic bile ducts
C0153455|ICD9CM|AB|156.8|Malig neo biliary NEC
C0153458|ICD9CM|PT|157.0|Malignant neoplasm of head of pancreas
C0153458|ICD9CM|AB|157.0|Mal neo pancreas head
C0153459|ICD9CM|PT|157.1|Malignant neoplasm of body of pancreas
C0153459|ICD9CM|AB|157.1|Mal neo pancreas body
C0153460|ICD9CM|PT|157.2|Malignant neoplasm of tail of pancreas
C0153460|ICD9CM|AB|157.2|Mal neo pancreas tail
C0153461|ICD9CM|PT|157.3|Malignant neoplasm of pancreatic duct
C0153461|ICD9CM|AB|157.3|Mal neo pancreatic duct
C0153463|ICD9CM|PT|157.8|Malignant neoplasm of other specified sites of pancreas
C0153463|ICD9CM|AB|157.8|Malig neo pancreas NEC
C0153464|ICD9CM|HT|158|Malignant neoplasm of retroperitoneum and peritoneum
C0153465|ICD9CM|PT|158.0|Malignant neoplasm of retroperitoneum
C0153465|ICD9CM|AB|158.0|Mal neo retroperitoneum
C0153466|ICD9CM|PT|158.8|Malignant neoplasm of specified parts of peritoneum
C0153466|ICD9CM|AB|158.8|Mal neo peritoneum NEC
C0153467|ICD9CM|PT|158.9|Malignant neoplasm of peritoneum, unspecified
C0153467|ICD9CM|AB|158.9|Mal neo peritoneum NOS
C0153468|ICD9CM|HT|159|Malignant neoplasm of other and ill-defined sites within the digestive organs and peritoneum
C0153471|ICD9CM|PT|159.8|Malignant neoplasm of other sites of digestive system and intra-abdominal organs
C0153471|ICD9CM|AB|159.8|Mal neo gi/intra-abd NEC
C0153472|ICD9CM|PT|159.9|Malignant neoplasm of ill-defined sites within the digestive organs and peritoneum
C0153472|ICD9CM|AB|159.9|Mal neo GI tract ill-def
C0153473|ICD9CM|HT|160|Malignant neoplasm of nasal cavities, middle ear, and accessory sinuses
C0153474|ICD9CM|PT|160.9|Malignant neoplasm of accessory sinus, unspecified
C0153474|ICD9CM|AB|160.9|Mal neo access sinus NOS
C0153475|ICD9CM|PT|160.1|Malignant neoplasm of auditory tube, middle ear, and mastoid air cells
C0153475|ICD9CM|AB|160.1|Malig neo middle ear
C0153476|ICD9CM|PT|160.2|Malignant neoplasm of maxillary sinus
C0153476|ICD9CM|AB|160.2|Mal neo maxillary sinus
C0153477|ICD9CM|PT|160.3|Malignant neoplasm of ethmoidal sinus
C0153477|ICD9CM|AB|160.3|Mal neo ethmoidal sinus
C0153478|ICD9CM|PT|160.4|Malignant neoplasm of frontal sinus
C0153478|ICD9CM|AB|160.4|Malig neo frontal sinus
C0153479|ICD9CM|PT|160.5|Malignant neoplasm of sphenoidal sinus
C0153479|ICD9CM|AB|160.5|Mal neo sphenoid sinus
C0153480|ICD9CM|PT|160.8|Malignant neoplasm of other accessory sinuses
C0153480|ICD9CM|AB|160.8|Mal neo access sinus NEC
C0153483|ICD9CM|PT|161.0|Malignant neoplasm of glottis
C0153483|ICD9CM|AB|161.0|Malignant neo glottis
C0153484|ICD9CM|PT|161.1|Malignant neoplasm of supraglottis
C0153484|ICD9CM|AB|161.1|Malig neo supraglottis
C0153485|ICD9CM|PT|161.2|Malignant neoplasm of subglottis
C0153485|ICD9CM|AB|161.2|Malig neo subglottis
C0153486|ICD9CM|PT|161.3|Malignant neoplasm of laryngeal cartilages
C0153486|ICD9CM|AB|161.3|Mal neo cartilage larynx
C0153487|ICD9CM|PT|161.8|Malignant neoplasm of other specified sites of larynx
C0153487|ICD9CM|AB|161.8|Malignant neo larynx NEC
C0153488|ICD9CM|HT|162|Malignant neoplasm of trachea, bronchus, and lung
C0153489|ICD9CM|PT|162.0|Malignant neoplasm of trachea
C0153489|ICD9CM|AB|162.0|Malignant neo trachea
C0153490|ICD9CM|PT|162.2|Malignant neoplasm of main bronchus
C0153490|ICD9CM|AB|162.2|Malig neo main bronchus
C0153491|ICD9CM|PT|162.4|Malignant neoplasm of middle lobe, bronchus or lung
C0153491|ICD9CM|AB|162.4|Mal neo middle lobe lung
C0153492|ICD9CM|PT|162.5|Malignant neoplasm of lower lobe, bronchus or lung
C0153492|ICD9CM|AB|162.5|Mal neo lower lobe lung
C0153493|ICD9CM|PT|162.8|Malignant neoplasm of other parts of bronchus or lung
C0153493|ICD9CM|AB|162.8|Mal neo bronch/lung NEC
C0153494|ICD9CM|HT|163|Malignant neoplasm of pleura
C0153494|ICD9CM|PT|163.9|Malignant neoplasm of pleura, unspecified
C0153494|ICD9CM|AB|163.9|Malig neopl pleura NOS
C0153497|ICD9CM|PT|163.8|Malignant neoplasm of other specified sites of pleura
C0153497|ICD9CM|AB|163.8|Malig neopl pleura NEC
C0153498|ICD9CM|HT|164|Malignant neoplasm of thymus, heart, and mediastinum
C0153500|ICD9CM|PT|164.1|Malignant neoplasm of heart
C0153500|ICD9CM|AB|164.1|Malignant neopl heart
C0153501|ICD9CM|PT|164.2|Malignant neoplasm of anterior mediastinum
C0153501|ICD9CM|AB|164.2|Mal neo ant mediastinum
C0153502|ICD9CM|PT|164.3|Malignant neoplasm of posterior mediastinum
C0153502|ICD9CM|AB|164.3|Mal neo post mediastinum
C0153503|ICD9CM|PT|164.8|Malignant neoplasm of other parts of mediastinum
C0153503|ICD9CM|AB|164.8|Mal neo mediastinum NEC
C0153504|ICD9CM|PT|164.9|Malignant neoplasm of mediastinum, part unspecified
C0153504|ICD9CM|AB|164.9|Mal neo mediastinum NOS
C0153506|ICD9CM|PT|165.0|Malignant neoplasm of upper respiratory tract, part unspecified
C0153506|ICD9CM|AB|165.0|Mal neo upper resp NOS
C0153507|ICD9CM|PT|165.8|Malignant neoplasm of other sites within the respiratory system and intrathoracic organs
C0153507|ICD9CM|AB|165.8|Mal neo thorax/resp NEC
C0153508|ICD9CM|PT|165.9|Malignant neoplasm of ill-defined sites within the respiratory system
C0153508|ICD9CM|AB|165.9|Mal neo resp system NOS
C0153509|ICD9CM|HT|170|Malignant neoplasm of bone and articular cartilage
C0153509|ICD9CM|PT|170.9|Malignant neoplasm of bone and articular cartilage, site unspecified
C0153509|ICD9CM|AB|170.9|Malig neopl bone NOS
C0153510|ICD9CM|PT|170.0|Malignant neoplasm of bones of skull and face, except mandible
C0153510|ICD9CM|AB|170.0|Mal neo skull/face bone
C0153511|ICD9CM|PT|170.1|Malignant neoplasm of mandible
C0153511|ICD9CM|AB|170.1|Malignant neo mandible
C0153512|ICD9CM|PT|170.2|Malignant neoplasm of vertebral column, excluding sacrum and coccyx
C0153512|ICD9CM|AB|170.2|Malig neo vertebrae
C0153513|ICD9CM|PT|170.3|Malignant neoplasm of ribs, sternum, and clavicle
C0153513|ICD9CM|AB|170.3|Mal neo ribs/stern/clav
C0153514|ICD9CM|PT|170.4|Malignant neoplasm of scapula and long bones of upper limb
C0153514|ICD9CM|AB|170.4|Mal neo long bones arm
C0153515|ICD9CM|PT|170.5|Malignant neoplasm of short bones of upper limb
C0153515|ICD9CM|AB|170.5|Mal neo bones wrist/hand
C0153516|ICD9CM|PT|170.6|Malignant neoplasm of pelvic bones, sacrum, and coccyx
C0153516|ICD9CM|AB|170.6|Mal neo pelvic girdle
C0153517|ICD9CM|PT|170.7|Malignant neoplasm of long bones of lower limb
C0153517|ICD9CM|AB|170.7|Mal neo long bones leg
C0153518|ICD9CM|PT|170.8|Malignant neoplasm of short bones of lower limb
C0153518|ICD9CM|AB|170.8|Mal neo bones ankle/foot
C0153519|ICD9CM|PT|171.9|Malignant neoplasm of connective and other soft tissue, site unspecified
C0153519|ICD9CM|HT|171|Malignant neoplasm of connective and other soft tissue
C0153519|ICD9CM|AB|171.9|Mal neo soft tissue NOS
C0153520|ICD9CM|PT|171.0|Malignant neoplasm of connective and other soft tissue of head, face, and neck
C0153520|ICD9CM|AB|171.0|Mal neo soft tissue head
C0153521|ICD9CM|PT|171.2|Malignant neoplasm of connective and other soft tissue of upper limb, including shoulder
C0153521|ICD9CM|AB|171.2|Mal neo soft tissue arm
C0153522|ICD9CM|PT|171.3|Malignant neoplasm of connective and other soft tissue of lower limb, including hip
C0153522|ICD9CM|AB|171.3|Mal neo soft tissue leg
C0153523|ICD9CM|PT|171.4|Malignant neoplasm of connective and other soft tissue of thorax
C0153523|ICD9CM|AB|171.4|Mal neo soft tis thorax
C0153524|ICD9CM|PT|171.5|Malignant neoplasm of connective and other soft tissue of abdomen
C0153524|ICD9CM|AB|171.5|Mal neo soft tis abdomen
C0153525|ICD9CM|PT|171.6|Malignant neoplasm of connective and other soft tissue of pelvis
C0153525|ICD9CM|AB|171.6|Mal neo soft tis pelvis
C0153527|ICD9CM|PT|171.8|Malignant neoplasm of other specified sites of connective and other soft tissue
C0153527|ICD9CM|AB|171.8|Mal neo soft tissue NEC
C0153529|ICD9CM|PT|172.0|Malignant melanoma of skin of lip
C0153529|ICD9CM|AB|172.0|Malig melanoma lip
C0153532|ICD9CM|PT|172.3|Malignant melanoma of skin of other and unspecified parts of face
C0153532|ICD9CM|AB|172.3|Mal melanom face NEC/NOS
C0153537|ICD9CM|PT|172.8|Malignant melanoma of other specified sites of skin
C0153537|ICD9CM|AB|172.8|Malig melanoma skin NEC
C0153539|ICD9CM|HT|173.0|Other malignant neoplasm of skin of lip
C0153549|ICD9CM|PT|174.1|Malignant neoplasm of central portion of female breast
C0153549|ICD9CM|AB|174.1|Mal neo breast-central
C0153550|ICD9CM|PT|174.2|Malignant neoplasm of upper-inner quadrant of female breast
C0153550|ICD9CM|AB|174.2|Mal neo breast up-inner
C0153551|ICD9CM|PT|174.3|Malignant neoplasm of lower-inner quadrant of female breast
C0153551|ICD9CM|AB|174.3|Mal neo breast low-inner
C0153552|ICD9CM|PT|174.4|Malignant neoplasm of upper-outer quadrant of female breast
C0153552|ICD9CM|AB|174.4|Mal neo breast up-outer
C0153553|ICD9CM|PT|174.5|Malignant neoplasm of lower-outer quadrant of female breast
C0153553|ICD9CM|AB|174.5|Mal neo breast low-outer
C0153554|ICD9CM|PT|174.6|Malignant neoplasm of axillary tail of female breast
C0153554|ICD9CM|AB|174.6|Mal neo breast-axillary
C0153555|ICD9CM|PT|174.8|Malignant neoplasm of other specified sites of female breast
C0153555|ICD9CM|AB|174.8|Malign neopl breast NEC
C0153558|ICD9CM|PT|175.0|Malignant neoplasm of nipple and areola of male breast
C0153558|ICD9CM|AB|175.0|Mal neo male nipple
C0153559|ICD9CM|PT|175.9|Malignant neoplasm of other and unspecified sites of male breast
C0153559|ICD9CM|AB|175.9|Mal neo male breast NEC
C0153560|ICD9CM|PT|176.0|Kaposi's sarcoma, skin
C0153560|ICD9CM|AB|176.0|Skin - kaposi's sarcoma
C0153561|ICD9CM|PT|176.1|Kaposi's sarcoma, soft tissue
C0153561|ICD9CM|AB|176.1|Sft tisue - kpsi's srcma
C0153562|ICD9CM|PT|176.2|Kaposi's sarcoma, palate
C0153562|ICD9CM|AB|176.2|Palate - kpsi's sarcoma
C0153563|ICD9CM|PT|176.3|Kaposi's sarcoma, gastrointestinal sites
C0153563|ICD9CM|AB|176.3|GI sites - kpsi's srcoma
C0153564|ICD9CM|PT|176.4|Kaposi's sarcoma, lung
C0153564|ICD9CM|AB|176.4|Lung - kaposi's sarcoma
C0153565|ICD9CM|PT|176.5|Kaposi's sarcoma, lymph nodes
C0153565|ICD9CM|AB|176.5|Lym nds - kpsi's sarcoma
C0153566|ICD9CM|PT|176.8|Kaposi's sarcoma, other specified sites
C0153566|ICD9CM|AB|176.8|Spf sts - kpsi's sarcoma
C0153567|ICD9CM|PT|179|Malignant neoplasm of uterus, part unspecified
C0153567|ICD9CM|AB|179|Malig neopl uterus NOS
C0153569|ICD9CM|PT|180.0|Malignant neoplasm of endocervix
C0153569|ICD9CM|AB|180.0|Malig neo endocervix
C0153570|ICD9CM|PT|180.1|Malignant neoplasm of exocervix
C0153570|ICD9CM|AB|180.1|Malig neo exocervix
C0153571|ICD9CM|PT|180.8|Malignant neoplasm of other specified sites of cervix
C0153571|ICD9CM|AB|180.8|Malig neo cervix NEC
C0153572|ICD9CM|PT|181|Malignant neoplasm of placenta
C0153572|ICD9CM|AB|181|Malignant neopl placenta
C0153574|ICD9CM|HT|182|Malignant neoplasm of body of uterus
C0153575|ICD9CM|PT|182.1|Malignant neoplasm of isthmus
C0153575|ICD9CM|AB|182.1|Mal neo uterine isthmus
C0153576|ICD9CM|PT|182.8|Malignant neoplasm of other specified sites of body of uterus
C0153576|ICD9CM|AB|182.8|Mal neo body uterus NEC
C0153577|ICD9CM|HT|183|Malignant neoplasm of ovary and other uterine adnexa
C0153579|ICD9CM|PT|183.2|Malignant neoplasm of fallopian tube
C0153579|ICD9CM|AB|183.2|Mal neo fallopian tube
C0153581|ICD9CM|PT|183.4|Malignant neoplasm of parametrium
C0153581|ICD9CM|AB|183.4|Malig neo parametrium
C0153583|ICD9CM|PT|183.8|Malignant neoplasm of other specified sites of uterine adnexa
C0153583|ICD9CM|AB|183.8|Mal neo adnexa NEC
C0153584|ICD9CM|PT|183.9|Malignant neoplasm of uterine adnexa, unspecified site
C0153584|ICD9CM|AB|183.9|Mal neo adnexa NOS
C0153585|ICD9CM|HT|184|Malignant neoplasm of other and unspecified female genital organs
C0153589|ICD9CM|PT|184.3|Malignant neoplasm of clitoris
C0153589|ICD9CM|AB|184.3|Malign neopl clitoris
C0153591|ICD9CM|PT|184.8|Malignant neoplasm of other specified sites of female genital organs
C0153591|ICD9CM|AB|184.8|Mal neo female genit NEC
C0153592|ICD9CM|PT|184.9|Malignant neoplasm of female genital organ, site unspecified
C0153592|ICD9CM|AB|184.9|Mal neo female genit NOS
C0153594|ICD9CM|HT|186|Malignant neoplasm of testis
C0153595|ICD9CM|PT|186.0|Malignant neoplasm of undescended testis
C0153595|ICD9CM|AB|186.0|Mal neo undescend testis
C0153596|ICD9CM|PT|186.9|Malignant neoplasm of other and unspecified testis
C0153596|ICD9CM|AB|186.9|Malig neo testis NEC
C0153597|ICD9CM|HT|187|Malignant neoplasm of penis and other male genital organs
C0153598|ICD9CM|PT|187.1|Malignant neoplasm of prepuce
C0153598|ICD9CM|AB|187.1|Malign neopl prepuce
C0153599|ICD9CM|PT|187.2|Malignant neoplasm of glans penis
C0153599|ICD9CM|AB|187.2|Malig neo glans penis
C0153600|ICD9CM|PT|187.3|Malignant neoplasm of body of penis
C0153600|ICD9CM|AB|187.3|Malig neo penis body
C0153601|ICD9CM|PT|187.4|Malignant neoplasm of penis, part unspecified
C0153601|ICD9CM|AB|187.4|Malig neo penis NOS
C0153602|ICD9CM|PT|187.5|Malignant neoplasm of epididymis
C0153602|ICD9CM|AB|187.5|Malig neo epididymis
C0153603|ICD9CM|PT|187.6|Malignant neoplasm of spermatic cord
C0153603|ICD9CM|AB|187.6|Mal neo spermatic cord
C0153604|ICD9CM|PT|187.7|Malignant neoplasm of scrotum
C0153604|ICD9CM|AB|187.7|Malign neopl scrotum
C0153605|ICD9CM|PT|187.8|Malignant neoplasm of other specified sites of male genital organs
C0153605|ICD9CM|AB|187.8|Mal neo male genital NEC
C0153606|ICD9CM|PT|187.9|Malignant neoplasm of male genital organ, site unspecified
C0153606|ICD9CM|AB|187.9|Mal neo male genital NOS
C0153611|ICD9CM|PT|188.3|Malignant neoplasm of anterior wall of urinary bladder
C0153611|ICD9CM|AB|188.3|Mal neo bladder-anterior
C0153612|ICD9CM|PT|188.4|Malignant neoplasm of posterior wall of urinary bladder
C0153612|ICD9CM|AB|188.4|Mal neo bladder-post
C0153613|ICD9CM|PT|188.5|Malignant neoplasm of bladder neck
C0153613|ICD9CM|AB|188.5|Mal neo bladder neck
C0153614|ICD9CM|PT|188.6|Malignant neoplasm of ureteric orifice
C0153614|ICD9CM|AB|188.6|Mal neo ureteric orifice
C0153615|ICD9CM|PT|188.7|Malignant neoplasm of urachus
C0153615|ICD9CM|AB|188.7|Malig neo urachus
C0153616|ICD9CM|PT|188.8|Malignant neoplasm of other specified sites of bladder
C0153616|ICD9CM|AB|188.8|Malig neo bladder NEC
C0153617|ICD9CM|HT|189|Malignant neoplasm of kidney and other and unspecified urinary organs
C0153618|ICD9CM|PT|189.1|Malignant neoplasm of renal pelvis
C0153618|ICD9CM|AB|189.1|Malig neo renal pelvis
C0153619|ICD9CM|PT|189.2|Malignant neoplasm of ureter
C0153619|ICD9CM|AB|189.2|Malign neopl ureter
C0153620|ICD9CM|PT|189.3|Malignant neoplasm of urethra
C0153620|ICD9CM|AB|189.3|Malign neopl urethra
C0153621|ICD9CM|PT|189.4|Malignant neoplasm of paraurethral glands
C0153621|ICD9CM|AB|189.4|Mal neo paraurethral
C0153622|ICD9CM|PT|189.8|Malignant neoplasm of other specified sites of urinary organs
C0153622|ICD9CM|AB|189.8|Mal neo urinary NEC
C0153625|ICD9CM|PT|190.0|Malignant neoplasm of eyeball, except conjunctiva, cornea, retina, and choroid
C0153625|ICD9CM|AB|190.0|Malign neopl eyeball
C0153626|ICD9CM|PT|190.1|Malignant neoplasm of orbit
C0153626|ICD9CM|AB|190.1|Malign neopl orbit
C0153627|ICD9CM|PT|190.2|Malignant neoplasm of lacrimal gland
C0153627|ICD9CM|AB|190.2|Mal neo lacrimal gland
C0153628|ICD9CM|PT|190.3|Malignant neoplasm of conjunctiva
C0153628|ICD9CM|AB|190.3|Mal neo conjunctiva
C0153629|ICD9CM|PT|190.4|Malignant neoplasm of cornea
C0153629|ICD9CM|AB|190.4|Malign neopl cornea
C0153630|ICD9CM|PT|190.6|Malignant neoplasm of choroid
C0153630|ICD9CM|AB|190.6|Malign neopl choroid
C0153631|ICD9CM|PT|190.7|Malignant neoplasm of lacrimal duct
C0153631|ICD9CM|AB|190.7|Mal neo lacrimal duct
C0153632|ICD9CM|PT|190.8|Malignant neoplasm of other specified sites of eye
C0153632|ICD9CM|AB|190.8|Malign neopl eye NEC
C0153633|ICD9CM|HT|191|Malignant neoplasm of brain
C0153633|ICD9CM|PT|191.9|Malignant neoplasm of brain, unspecified
C0153633|ICD9CM|AB|191.9|Malig neo brain NOS
C0153634|ICD9CM|PT|191.0|Malignant neoplasm of cerebrum, except lobes and ventricles
C0153634|ICD9CM|AB|191.0|Malign neopl cerebrum
C0153635|ICD9CM|PT|191.1|Malignant neoplasm of frontal lobe
C0153635|ICD9CM|AB|191.1|Malig neo frontal lobe
C0153636|ICD9CM|PT|191.2|Malignant neoplasm of temporal lobe
C0153636|ICD9CM|AB|191.2|Mal neo temporal lobe
C0153637|ICD9CM|PT|191.3|Malignant neoplasm of parietal lobe
C0153637|ICD9CM|AB|191.3|Mal neo parietal lobe
C0153638|ICD9CM|PT|191.4|Malignant neoplasm of occipital lobe
C0153638|ICD9CM|AB|191.4|Mal neo occipital lobe
C0153640|ICD9CM|PT|191.6|Malignant neoplasm of cerebellum nos
C0153640|ICD9CM|AB|191.6|Mal neo cerebellum NOS
C0153641|ICD9CM|PT|191.7|Malignant neoplasm of brain stem
C0153641|ICD9CM|AB|191.7|Mal neo brain stem
C0153642|ICD9CM|PT|191.8|Malignant neoplasm of other parts of brain
C0153642|ICD9CM|AB|191.8|Malig neo brain NEC
C0153643|ICD9CM|PT|192.9|Malignant neoplasm of nervous system, part unspecified
C0153643|ICD9CM|HT|192|Malignant neoplasm of other and unspecified parts of nervous system
C0153643|ICD9CM|AB|192.9|Mal neo nervous syst NOS
C0153644|ICD9CM|PT|192.0|Malignant neoplasm of cranial nerves
C0153644|ICD9CM|AB|192.0|Mal neo cranial nerves
C0153645|ICD9CM|PT|192.1|Malignant neoplasm of cerebral meninges
C0153645|ICD9CM|AB|192.1|Mal neo cerebral mening
C0153646|ICD9CM|PT|192.2|Malignant neoplasm of spinal cord
C0153646|ICD9CM|AB|192.2|Mal neo spinal cord
C0153647|ICD9CM|PT|192.3|Malignant neoplasm of spinal meninges
C0153647|ICD9CM|AB|192.3|Mal neo spinal meninges
C0153648|ICD9CM|PT|192.8|Malignant neoplasm of other specified sites of nervous system
C0153648|ICD9CM|AB|192.8|Mal neo nervous syst NEC
C0153651|ICD9CM|HT|194|Malignant neoplasm of other endocrine glands and related structures
C0153651|ICD9CM|PT|194.8|Malignant neoplasm of other endocrine glands and related structures
C0153651|ICD9CM|AB|194.8|Mal neo endocrine NEC
C0153653|ICD9CM|PT|194.1|Malignant neoplasm of parathyroid gland
C0153653|ICD9CM|AB|194.1|Malig neo parathyroid
C0153654|ICD9CM|PT|194.3|Malignant neoplasm of pituitary gland and craniopharyngeal duct
C0153654|ICD9CM|AB|194.3|Malig neo pituitary
C0153655|ICD9CM|PT|194.4|Malignant neoplasm of pineal gland
C0153655|ICD9CM|AB|194.4|Malign neo pineal gland
C0153656|ICD9CM|PT|194.5|Malignant neoplasm of carotid body
C0153656|ICD9CM|AB|194.5|Mal neo carotid body
C0153658|ICD9CM|PT|194.9|Malignant neoplasm of endocrine gland, site unspecified
C0153658|ICD9CM|AB|194.9|Mal neo endocrine NOS
C0153659|ICD9CM|HT|195|Malignant neoplasm of other and ill-defined sites
C0153660|ICD9CM|PT|195.0|Malignant neoplasm of head, face, and neck
C0153660|ICD9CM|AB|195.0|Mal neo head/face/neck
C0153661|ICD9CM|PT|195.1|Malignant neoplasm of thorax
C0153661|ICD9CM|AB|195.1|Malign neopl thorax
C0153662|ICD9CM|PT|195.2|Malignant neoplasm of abdomen
C0153662|ICD9CM|AB|195.2|Malig neo abdomen
C0153663|ICD9CM|PT|195.3|Malignant neoplasm of pelvis
C0153663|ICD9CM|AB|195.3|Malign neopl pelvis
C0153664|ICD9CM|PT|195.4|Malignant neoplasm of upper limb
C0153664|ICD9CM|AB|195.4|Malign neopl arm
C0153665|ICD9CM|PT|195.5|Malignant neoplasm of lower limb
C0153665|ICD9CM|AB|195.5|Malign neopl leg
C0153666|ICD9CM|PT|195.8|Malignant neoplasm of other specified sites
C0153666|ICD9CM|AB|195.8|Malig neo site NEC
C0153668|ICD9CM|PT|196.0|Secondary and unspecified malignant neoplasm of lymph nodes of head, face, and neck
C0153668|ICD9CM|AB|196.0|Mal neo lymph-head/neck
C0153671|ICD9CM|PT|196.3|Secondary and unspecified malignant neoplasm of lymph nodes of axilla and upper limb
C0153671|ICD9CM|AB|196.3|Mal neo lymph-axilla/arm
C0153675|ICD9CM|HT|197|Secondary malignant neoplasm of respiratory and digestive systems
C0153676|ICD9CM|PT|197.0|Secondary malignant neoplasm of lung
C0153676|ICD9CM|AB|197.0|Secondary malig neo lung
C0153677|ICD9CM|PT|197.1|Secondary malignant neoplasm of mediastinum
C0153677|ICD9CM|AB|197.1|Sec mal neo mediastinum
C0153678|ICD9CM|PT|197.2|Secondary malignant neoplasm of pleura
C0153678|ICD9CM|AB|197.2|Second malig neo pleura
C0153681|ICD9CM|PT|197.5|Secondary malignant neoplasm of large intestine and rectum
C0153681|ICD9CM|AB|197.5|Sec malig neo lg bowel
C0153683|ICD9CM|PT|197.8|Secondary malignant neoplasm of other digestive organs and spleen
C0153683|ICD9CM|AB|197.8|Sec mal neo GI NEC
C0153684|ICD9CM|HT|198|Secondary malignant neoplasm of other specified sites
C0153684|ICD9CM|HT|198.8|Secondary malignant neoplasm of other specified sites
C0153684|ICD9CM|PT|198.89|Secondary malignant neoplasm of other specified sites
C0153684|ICD9CM|AB|198.89|Secondary malig neo NEC
C0153685|ICD9CM|PT|198.0|Secondary malignant neoplasm of kidney
C0153685|ICD9CM|AB|198.0|Second malig neo kidney
C0153687|ICD9CM|PT|198.2|Secondary malignant neoplasm of skin
C0153687|ICD9CM|AB|198.2|Secondary malig neo skin
C0153688|ICD9CM|PT|198.3|Secondary malignant neoplasm of brain and spinal cord
C0153688|ICD9CM|AB|198.3|Sec mal neo brain/spine
C0153689|ICD9CM|PT|198.4|Secondary malignant neoplasm of other parts of nervous system
C0153689|ICD9CM|AB|198.4|Sec malig neo nerve NEC
C0153690|ICD9CM|PT|198.5|Secondary malignant neoplasm of bone and bone marrow
C0153690|ICD9CM|AB|198.5|Secondary malig neo bone
C0153691|ICD9CM|PT|198.7|Secondary malignant neoplasm of adrenal gland
C0153691|ICD9CM|AB|198.7|Second malig neo adrenal
C0153693|ICD9CM|PT|198.82|Secondary malignant neoplasm of genital organs
C0153693|ICD9CM|AB|198.82|Second malig neo genital
C0153696|ICD9CM|PT|200.01|Reticulosarcoma, lymph nodes of head, face, and neck
C0153696|ICD9CM|AB|200.01|Reticulosarcoma head
C0153697|ICD9CM|PT|200.02|Reticulosarcoma, intrathoracic lymph nodes
C0153697|ICD9CM|AB|200.02|Reticulosarcoma thorax
C0153698|ICD9CM|PT|200.03|Reticulosarcoma, intra-abdominal lymph nodes
C0153698|ICD9CM|AB|200.03|Reticulosarcoma abdom
C0153699|ICD9CM|PT|200.04|Reticulosarcoma, lymph nodes of axilla and upper limb
C0153699|ICD9CM|AB|200.04|Reticulosarcoma axilla
C0153700|ICD9CM|PT|200.05|Reticulosarcoma, lymph nodes of inguinal region and lower limb
C0153700|ICD9CM|AB|200.05|Reticulosarcoma inguin
C0153701|ICD9CM|PT|200.06|Reticulosarcoma, intrapelvic lymph nodes
C0153701|ICD9CM|AB|200.06|Reticulosarcoma pelvic
C0153702|ICD9CM|AB|200.07|Reticulosarcoma spleen
C0153702|ICD9CM|PT|200.07|Reticulosarcoma, spleen
C0153703|ICD9CM|PT|200.08|Reticulosarcoma, lymph nodes of multiple sites
C0153703|ICD9CM|AB|200.08|Reticulosarcoma mult
C0153704|ICD9CM|PT|200.11|Lymphosarcoma, lymph nodes of head, face, and neck
C0153704|ICD9CM|AB|200.11|Lymphosarcoma head
C0153705|ICD9CM|PT|200.12|Lymphosarcoma, intrathoracic lymph nodes
C0153705|ICD9CM|AB|200.12|Lymphosarcoma thorax
C0153706|ICD9CM|PT|200.13|Lymphosarcoma, intra-abdominal lymph nodes
C0153706|ICD9CM|AB|200.13|Lymphosarcoma abdom
C0153707|ICD9CM|PT|200.14|Lymphosarcoma, lymph nodes of axilla and upper limb
C0153707|ICD9CM|AB|200.14|Lymphosarcoma axilla
C0153708|ICD9CM|PT|200.15|Lymphosarcoma, lymph nodes of inguinal region and lower limb
C0153708|ICD9CM|AB|200.15|Lymphosarcoma inguin
C0153709|ICD9CM|PT|200.16|Lymphosarcoma, intrapelvic lymph nodes
C0153709|ICD9CM|AB|200.16|Lymphosarcoma pelvic
C0153710|ICD9CM|AB|200.17|Lymphosarcoma spleen
C0153710|ICD9CM|PT|200.17|Lymphosarcoma, spleen
C0153711|ICD9CM|PT|200.18|Lymphosarcoma, lymph nodes of multiple sites
C0153711|ICD9CM|AB|200.18|Lymphosarcoma mult
C0153712|ICD9CM|PT|200.21|Burkitt's tumor or lymphoma, lymph nodes of head, face, and neck
C0153712|ICD9CM|AB|200.21|Burkitt's tumor head
C0153713|ICD9CM|PT|200.22|Burkitt's tumor or lymphoma, intrathoracic lymph nodes
C0153713|ICD9CM|AB|200.22|Burkitt's tumor thorax
C0153714|ICD9CM|PT|200.23|Burkitt's tumor or lymphoma, intra-abdominal lymph nodes
C0153714|ICD9CM|AB|200.23|Burkitt's tumor abdom
C0153715|ICD9CM|PT|200.24|Burkitt's tumor or lymphoma, lymph nodes of axilla and upper limb
C0153715|ICD9CM|AB|200.24|Burkitt's tumor axilla
C0153716|ICD9CM|PT|200.25|Burkitt's tumor or lymphoma, lymph nodes of inguinal region and lower limb
C0153716|ICD9CM|AB|200.25|Burkitt's tumor inguin
C0153717|ICD9CM|PT|200.26|Burkitt's tumor or lymphoma, intrapelvic lymph nodes
C0153717|ICD9CM|AB|200.26|Burkitt's tumor pelvic
C0153719|ICD9CM|PT|200.28|Burkitt's tumor or lymphoma, lymph nodes of multiple sites
C0153719|ICD9CM|AB|200.28|Burkitt's tumor mult
C0153720|ICD9CM|PT|200.81|Other named variants of lymphosarcoma and reticulosarcoma, lymph nodes of head, face, and neck
C0153720|ICD9CM|AB|200.81|Mixed lymphosarc head
C0153721|ICD9CM|PT|200.82|Other named variants of lymphosarcoma and reticulosarcoma,intrathoracic lymph nodes
C0153721|ICD9CM|AB|200.82|Mixed lymphosarc thorax
C0153722|ICD9CM|PT|200.83|Other named variants of lymphosarcoma and reticulosarcoma, intra-abdominal lymph nodes
C0153722|ICD9CM|AB|200.83|Mixed lymphosarc abdom
C0153723|ICD9CM|PT|200.84|Other named variants of lymphosarcoma and reticulosarcoma, lymph nodes of axilla and upper limb
C0153723|ICD9CM|AB|200.84|Mixed lymphosarc axilla
C0153724|ICD9CM|PT|200.85|Other named variants of lymphosarcoma and reticulosarcoma, lymph nodes of inguinal region and lower limb
C0153724|ICD9CM|AB|200.85|Mixed lymphosarc inguin
C0153725|ICD9CM|PT|200.86|Other named variants of lymphosarcoma and reticulosarcoma, intrapelvic lymph nodes
C0153725|ICD9CM|AB|200.86|Mixed lymphosarc pelvic
C0153726|ICD9CM|PT|200.87|Other named variants of lymphosarcoma and reticulosarcoma, spleen
C0153726|ICD9CM|AB|200.87|Mixed lymphosarc spleen
C0153727|ICD9CM|PT|200.88|Other named variants of lymphosarcoma and reticulosarcoma, lymph nodes of multiple sites
C0153727|ICD9CM|AB|200.88|Mixed lymphosarc mult
C0153728|ICD9CM|PT|201.01|Hodgkin's paragranuloma, lymph nodes of head, face, and neck
C0153728|ICD9CM|AB|201.01|Hodgkins paragran head
C0153729|ICD9CM|PT|201.02|Hodgkin's paragranuloma, intrathoracic lymph nodes
C0153729|ICD9CM|AB|201.02|Hodgkins paragran thorax
C0153730|ICD9CM|PT|201.03|Hodgkin's paragranuloma, intra-abdominal lymph nodes
C0153730|ICD9CM|AB|201.03|Hodgkins paragran abdom
C0153731|ICD9CM|PT|201.04|Hodgkin's paragranuloma, lymph nodes of axilla and upper limb
C0153731|ICD9CM|AB|201.04|Hodgkins paragran axilla
C0153732|ICD9CM|PT|201.05|Hodgkin's paragranuloma, lymph nodes of inguinal region and lower limb
C0153732|ICD9CM|AB|201.05|Hodgkins paragran inguin
C0153733|ICD9CM|PT|201.06|Hodgkin's paragranuloma, intrapelvic lymph nodes
C0153733|ICD9CM|AB|201.06|Hodgkins paragran pelvic
C0153734|ICD9CM|PT|201.07|Hodgkin's paragranuloma, spleen
C0153734|ICD9CM|AB|201.07|Hodgkins paragran spleen
C0153736|ICD9CM|PT|201.11|Hodgkin's granuloma, lymph nodes of head, face, and neck
C0153736|ICD9CM|AB|201.11|Hodgkins granulom head
C0153737|ICD9CM|PT|201.12|Hodgkin's granuloma, intrathoracic lymph nodes
C0153737|ICD9CM|AB|201.12|Hodgkins granulom thorax
C0153738|ICD9CM|PT|201.13|Hodgkin's granuloma, intra-abdominal lymph nodes
C0153738|ICD9CM|AB|201.13|Hodgkins granulom abdom
C0153739|ICD9CM|PT|201.14|Hodgkin's granuloma, lymph nodes of axilla and upper limb
C0153739|ICD9CM|AB|201.14|Hodgkins granulom axilla
C0153740|ICD9CM|PT|201.15|Hodgkin's granuloma, lymph nodes of inguinal region and lower limb
C0153740|ICD9CM|AB|201.15|Hodgkins granulom inguin
C0153741|ICD9CM|PT|201.16|Hodgkin's granuloma, intrapelvic lymph nodes
C0153741|ICD9CM|AB|201.16|Hodgkins granulom pelvic
C0153742|ICD9CM|PT|201.18|Hodgkin's granuloma, lymph nodes of multiple sites
C0153742|ICD9CM|AB|201.18|Hodgkins granulom mult
C0153744|ICD9CM|PT|201.21|Hodgkin's sarcoma, lymph nodes of head, face, and neck
C0153744|ICD9CM|AB|201.21|Hodgkins sarcoma head
C0153745|ICD9CM|PT|201.22|Hodgkin's sarcoma, intrathoracic lymph nodes
C0153745|ICD9CM|AB|201.22|Hodgkins sarcoma thorax
C0153746|ICD9CM|PT|201.23|Hodgkin's sarcoma, intra-abdominal lymph nodes
C0153746|ICD9CM|AB|201.23|Hodgkins sarcoma abdom
C0153747|ICD9CM|PT|201.24|Hodgkin's sarcoma, lymph nodes of axilla and upper limb
C0153747|ICD9CM|AB|201.24|Hodgkins sarcoma axilla
C0153748|ICD9CM|PT|201.25|Hodgkin's sarcoma, lymph nodes of inguinal region and lower limb
C0153748|ICD9CM|AB|201.25|Hodgkins sarcoma inguin
C0153749|ICD9CM|PT|201.26|Hodgkin's sarcoma, intrapelvic lymph nodes
C0153749|ICD9CM|AB|201.26|Hodgkins sarcoma pelvic
C0153750|ICD9CM|AB|201.27|Hodgkins sarcoma spleen
C0153750|ICD9CM|PT|201.27|Hodgkin's sarcoma, spleen
C0153751|ICD9CM|PT|201.28|Hodgkin's sarcoma, lymph nodes of multiple sites
C0153751|ICD9CM|AB|201.28|Hodgkins sarcoma mult
C0153752|ICD9CM|PT|201.41|Hodgkin's disease, lymphocytic-histiocytic predominance, lymph nodes of head, face, and neck
C0153752|ICD9CM|AB|201.41|Hodg lymph-histio head
C0153753|ICD9CM|PT|201.42|Hodgkin's disease, lymphocytic-histiocytic predominance, intrathoracic lymph nodes
C0153753|ICD9CM|AB|201.42|Hodg lymph-histio thorax
C0153754|ICD9CM|PT|201.43|Hodgkin's disease, lymphocytic-histiocytic predominance, intra-abdominal lymph nodes
C0153754|ICD9CM|AB|201.43|Hodg lymph-histio abdom
C0153755|ICD9CM|PT|201.44|Hodgkin's disease, lymphocytic-histiocytic predominance, lymph nodes of axilla and upper limb
C0153755|ICD9CM|AB|201.44|Hodg lymph-histio axilla
C0153756|ICD9CM|PT|201.45|Hodgkin's disease, lymphocytic-histiocytic predominance, lymph nodes of inguinal region and lower limb
C0153756|ICD9CM|AB|201.45|Hodg lymph-histio inguin
C0153757|ICD9CM|PT|201.46|Hodgkin's disease, lymphocytic-histiocytic predominance, intrapelvic lymph nodes
C0153757|ICD9CM|AB|201.46|Hodg lymph-histio pelvic
C0153758|ICD9CM|PT|201.47|Hodgkin's disease, lymphocytic-histiocytic predominance, spleen
C0153758|ICD9CM|AB|201.47|Hodg lymph-histio spleen
C0153759|ICD9CM|PT|201.48|Hodgkin's disease, lymphocytic-histiocytic predominance, lymph nodes of multiple sites
C0153759|ICD9CM|AB|201.48|Hodg lymph-histio mult
C0153760|ICD9CM|PT|201.51|Hodgkin's disease, nodular sclerosis, lymph nodes of head, face, and neck
C0153760|ICD9CM|AB|201.51|Hodg nodul sclero head
C0153761|ICD9CM|PT|201.52|Hodgkin's disease, nodular sclerosis, intrathoracic lymph nodes
C0153761|ICD9CM|AB|201.52|Hodg nodul sclero thorax
C0153762|ICD9CM|PT|201.53|Hodgkin's disease, nodular sclerosis, intra-abdominal lymph nodes
C0153762|ICD9CM|AB|201.53|Hodg nodul sclero abdom
C0153763|ICD9CM|PT|201.54|Hodgkin's disease, nodular sclerosis, lymph nodes of axilla and upper limb
C0153763|ICD9CM|AB|201.54|Hodg nodul sclero axilla
C0153764|ICD9CM|PT|201.55|Hodgkin's disease, nodular sclerosis, lymph nodes of inguinal region and lower limb
C0153764|ICD9CM|AB|201.55|Hodg nodul sclero inguin
C0153765|ICD9CM|PT|201.56|Hodgkin's disease, nodular sclerosis, intrapelvic lymph nodes
C0153765|ICD9CM|AB|201.56|Hodg nodul sclero pelvic
C0153766|ICD9CM|PT|201.57|Hodgkin's disease, nodular sclerosis, spleen
C0153766|ICD9CM|AB|201.57|Hodg nodul sclero spleen
C0153767|ICD9CM|PT|201.58|Hodgkin's disease, nodular sclerosis, lymph nodes of multiple sites
C0153767|ICD9CM|AB|201.58|Hodg nodul sclero mult
C0153768|ICD9CM|PT|201.61|Hodgkin's disease, mixed cellularity, lymph nodes of head, face, and neck
C0153768|ICD9CM|AB|201.61|Hodgkins mix cell head
C0153769|ICD9CM|PT|201.62|Hodgkin's disease, mixed cellularity, intrathoracic lymph nodes
C0153769|ICD9CM|AB|201.62|Hodgkins mix cell thorax
C0153770|ICD9CM|PT|201.63|Hodgkin's disease, mixed cellularity, intra-abdominal lymph nodes
C0153770|ICD9CM|AB|201.63|Hodgkins mix cell abdom
C0153771|ICD9CM|PT|201.64|Hodgkin's disease, mixed cellularity, lymph nodes of axilla and upper limb
C0153771|ICD9CM|AB|201.64|Hodgkins mix cell axilla
C0153772|ICD9CM|PT|201.65|Hodgkin's disease, mixed cellularity, lymph nodes of inguinal region and lower limb
C0153772|ICD9CM|AB|201.65|Hodgkins mix cell inguin
C0153773|ICD9CM|PT|201.66|Hodgkin's disease, mixed cellularity, intrapelvic lymph nodes
C0153773|ICD9CM|AB|201.66|Hodgkins mix cell pelvic
C0153774|ICD9CM|PT|201.67|Hodgkin's disease, mixed cellularity, spleen
C0153774|ICD9CM|AB|201.67|Hodgkins mix cell spleen
C0153775|ICD9CM|PT|201.68|Hodgkin's disease, mixed cellularity, lymph nodes of multiple sites
C0153775|ICD9CM|AB|201.68|Hodgkins mix cell mult
C0153776|ICD9CM|PT|201.71|Hodgkin's disease, lymphocytic depletion, lymph nodes of head, face, and neck
C0153776|ICD9CM|AB|201.71|Hodg lymph deplet head
C0153777|ICD9CM|PT|201.72|Hodgkin's disease, lymphocytic depletion, intrathoracic lymph nodes
C0153777|ICD9CM|AB|201.72|Hodg lymph deplet thorax
C0153778|ICD9CM|PT|201.73|Hodgkin's disease, lymphocytic depletion, intra-abdominal lymph nodes
C0153778|ICD9CM|AB|201.73|Hodg lymph deplet abdom
C0153779|ICD9CM|PT|201.74|Hodgkin's disease, lymphocytic depletion, lymph nodes of axilla and upper limb
C0153779|ICD9CM|AB|201.74|Hodg lymph deplet axilla
C0153780|ICD9CM|PT|201.75|Hodgkin's disease, lymphocytic depletion, lymph nodes of inguinal region and lower limb
C0153780|ICD9CM|AB|201.75|Hodg lymph deplet inguin
C0153781|ICD9CM|PT|201.76|Hodgkin's disease, lymphocytic depletion, intrapelvic lymph nodes
C0153781|ICD9CM|AB|201.76|Hodg lymph deplet pelvic
C0153782|ICD9CM|PT|201.77|Hodgkin's disease, lymphocytic depletion, spleen
C0153782|ICD9CM|AB|201.77|Hodg lymph deplet spleen
C0153783|ICD9CM|PT|201.78|Hodgkin's disease, lymphocytic depletion, lymph nodes of multiple sites
C0153783|ICD9CM|AB|201.78|Hodg lymph deplet mult
C0153785|ICD9CM|PT|201.91|Hodgkin's disease, unspecified type, lymph nodes of head, face, and neck
C0153785|ICD9CM|AB|201.91|Hodgkins dis NOS head
C0153786|ICD9CM|PT|201.92|Hodgkin's disease, unspecified type, intrathoracic lymph nodes
C0153786|ICD9CM|AB|201.92|Hodgkins dis NOS thorax
C0153788|ICD9CM|PT|201.94|Hodgkin's disease, unspecified type, lymph nodes of axilla and upper limb
C0153788|ICD9CM|AB|201.94|Hodgkins dis NOS axilla
C0153789|ICD9CM|PT|201.95|Hodgkin's disease, unspecified type, lymph nodes of inguinal region and lower limb
C0153789|ICD9CM|AB|201.95|Hodgkins dis NOS inguin
C0153790|ICD9CM|PT|201.96|Hodgkin's disease, unspecified type, intrapelvic lymph nodes
C0153790|ICD9CM|AB|201.96|Hodgkins dis NOS pelvic
C0153791|ICD9CM|AB|201.97|Hodgkins dis NOS spleen
C0153791|ICD9CM|PT|201.97|Hodgkin's disease, unspecified type, spleen
C0153792|ICD9CM|PT|201.98|Hodgkin's disease, unspecified type, lymph nodes of multiple sites
C0153792|ICD9CM|AB|201.98|Hodgkins dis NOS mult
C0153793|ICD9CM|HT|202|Other malignant neoplasms of lymphoid and histiocytic tissue
C0153794|ICD9CM|PT|202.01|Nodular lymphoma, lymph nodes of head, face, and neck
C0153794|ICD9CM|AB|202.01|Nodular lymphoma head
C0153795|ICD9CM|PT|202.02|Nodular lymphoma, intrathoracic lymph nodes
C0153795|ICD9CM|AB|202.02|Nodular lymphoma thorax
C0153796|ICD9CM|PT|202.03|Nodular lymphoma, intra-abdominal lymph nodes
C0153796|ICD9CM|AB|202.03|Nodular lymphoma abdom
C0153797|ICD9CM|PT|202.04|Nodular lymphoma, lymph nodes of axilla and upper limb
C0153797|ICD9CM|AB|202.04|Nodular lymphoma axilla
C0153798|ICD9CM|PT|202.05|Nodular lymphoma, lymph nodes of inguinal region and lower limb
C0153798|ICD9CM|AB|202.05|Nodular lymphoma inguin
C0153799|ICD9CM|PT|202.06|Nodular lymphoma, intrapelvic lymph nodes
C0153799|ICD9CM|AB|202.06|Nodular lymphoma pelvic
C0153800|ICD9CM|AB|202.07|Nodular lymphoma spleen
C0153800|ICD9CM|PT|202.07|Nodular lymphoma, spleen
C0153801|ICD9CM|PT|202.08|Nodular lymphoma, lymph nodes of multiple sites
C0153801|ICD9CM|AB|202.08|Nodular lymphoma mult
C0153802|ICD9CM|PT|202.11|Mycosis fungoides, lymph nodes of head, face, and neck
C0153802|ICD9CM|AB|202.11|Mycosis fungoides head
C0153803|ICD9CM|PT|202.12|Mycosis fungoides, intrathoracic lymph nodes
C0153803|ICD9CM|AB|202.12|Mycosis fungoides thorax
C0153804|ICD9CM|PT|202.13|Mycosis fungoides, intra-abdominal lymph nodes
C0153804|ICD9CM|AB|202.13|Mycosis fungoides abdom
C0153805|ICD9CM|PT|202.14|Mycosis fungoides, lymph nodes of axilla and upper limb
C0153805|ICD9CM|AB|202.14|Mycosis fungoides axilla
C0153806|ICD9CM|PT|202.15|Mycosis fungoides, lymph nodes of inguinal region and lower limb
C0153806|ICD9CM|AB|202.15|Mycosis fungoides inguin
C0153807|ICD9CM|PT|202.16|Mycosis fungoides, intrapelvic lymph nodes
C0153807|ICD9CM|AB|202.16|Mycosis fungoides pelvic
C0153808|ICD9CM|AB|202.17|Mycosis fungoides spleen
C0153808|ICD9CM|PT|202.17|Mycosis fungoides, spleen
C0153809|ICD9CM|PT|202.18|Mycosis fungoides, lymph nodes of multiple sites
C0153809|ICD9CM|AB|202.18|Mycosis fungoides mult
C0153810|ICD9CM|PT|202.21|Sezary's disease, lymph nodes of head, face, and neck
C0153810|ICD9CM|AB|202.21|Sezary's disease head
C0153811|ICD9CM|PT|202.22|Sezary's disease, intrathoracic lymph nodes
C0153811|ICD9CM|AB|202.22|Sezary's disease thorax
C0153812|ICD9CM|PT|202.23|Sezary's disease, intra-abdominal lymph nodes
C0153812|ICD9CM|AB|202.23|Sezary's disease abdom
C0153813|ICD9CM|PT|202.24|Sezary's disease, lymph nodes of axilla and upper limb
C0153813|ICD9CM|AB|202.24|Sezary's disease axilla
C0153814|ICD9CM|PT|202.25|Sezary's disease, lymph nodes of inguinal region and lower limb
C0153814|ICD9CM|AB|202.25|Sezary's disease inguin
C0153815|ICD9CM|PT|202.26|Sezary's disease, intrapelvic lymph nodes
C0153815|ICD9CM|AB|202.26|Sezary's disease pelvic
C0153816|ICD9CM|AB|202.27|Sezary's disease spleen
C0153816|ICD9CM|PT|202.27|Sezary's disease, spleen
C0153817|ICD9CM|PT|202.28|Sezary's disease, lymph nodes of multiple sites
C0153817|ICD9CM|AB|202.28|Sezary's disease mult
C0153826|ICD9CM|PT|202.41|Leukemic reticuloendotheliosis, lymph nodes of head, face, and neck
C0153826|ICD9CM|AB|202.41|Hairy-cell leukem head
C0153827|ICD9CM|PT|202.42|Leukemic reticuloendotheliosis, intrathoracic lymph nodes
C0153827|ICD9CM|AB|202.42|Hairy-cell leukem thorax
C0153828|ICD9CM|PT|202.43|Leukemic reticuloendotheliosis, intra-abdominal lymph nodes
C0153828|ICD9CM|AB|202.43|Hairy-cell leukem abdom
C0153829|ICD9CM|PT|202.44|Leukemic reticuloendotheliosis, lymph nodes of axilla and upper arm
C0153829|ICD9CM|AB|202.44|Hairy-cell leukem axilla
C0153830|ICD9CM|PT|202.45|Leukemic reticuloendotheliosis, lymph nodes of inguinal region and lower limb
C0153830|ICD9CM|AB|202.45|Hairy-cell leukem inguin
C0153831|ICD9CM|PT|202.46|Leukemic reticuloendotheliosis, intrapelvic lymph nodes
C0153831|ICD9CM|AB|202.46|Hairy-cell leukem pelvic
C0153832|ICD9CM|PT|202.47|Leukemic reticuloendotheliosis, spleen
C0153832|ICD9CM|AB|202.47|Hairy-cell leukem spleen
C0153833|ICD9CM|PT|202.48|Leukemic reticuloendotheliosis, lymph nodes of multiple sites
C0153833|ICD9CM|AB|202.48|Hairy-cell leukem mult
C0153843|ICD9CM|PT|202.62|Malignant mast cell tumors, intrathoracic lymph nodes
C0153843|ICD9CM|AB|202.62|Mal mastocytosis thorax
C0153844|ICD9CM|PT|202.63|Malignant mast cell tumors, intra-abdominal lymph nodes
C0153844|ICD9CM|AB|202.63|Mal mastocytosis abdom
C0153845|ICD9CM|PT|202.64|Malignant mast cell tumors, lymph nodes of axilla and upper limb
C0153845|ICD9CM|AB|202.64|Mal mastocytosis axilla
C0153846|ICD9CM|PT|202.65|Malignant mast cell tumors, lymph nodes of inguinal region and lower limb
C0153846|ICD9CM|AB|202.65|Mal mastocytosis inguin
C0153847|ICD9CM|PT|202.66|Malignant mast cell tumors, intrapelvic lymph nodes
C0153847|ICD9CM|AB|202.66|Mal mastocytosis pelvic
C0153848|ICD9CM|PT|202.67|Malignant mast cell tumors, spleen
C0153848|ICD9CM|AB|202.67|Mal mastocytosis spleen
C0153849|ICD9CM|PT|202.68|Malignant mast cell tumors, lymph nodes of multiple sites
C0153849|ICD9CM|AB|202.68|Mal mastocytosis mult
C0153850|ICD9CM|PT|202.81|Other malignant lymphomas, lymph nodes of head, face, and neck
C0153850|ICD9CM|AB|202.81|Lymphomas NEC head
C0153851|ICD9CM|PT|202.82|Other malignant lymphomas, intrathoracic lymph nodes
C0153851|ICD9CM|AB|202.82|Lymphomas NEC thorax
C0153852|ICD9CM|PT|202.83|Other malignant lymphomas, intra-abdominal lymph nodes
C0153852|ICD9CM|AB|202.83|Lymphomas NEC abdom
C0153853|ICD9CM|PT|202.84|Other malignant lymphomas, lymph nodes of axilla and upper limb
C0153853|ICD9CM|AB|202.84|Lymphomas NEC axilla
C0153854|ICD9CM|PT|202.85|Other malignant lymphomas, lymph nodes of inguinal region and lower limb
C0153854|ICD9CM|AB|202.85|Lymphomas NEC inguin
C0153855|ICD9CM|PT|202.86|Other malignant lymphomas, intrapelvic lymph nodes
C0153855|ICD9CM|AB|202.86|Lymphomas NEC pelvic
C0153856|ICD9CM|PT|202.87|Other malignant lymphomas, spleen
C0153856|ICD9CM|AB|202.87|Lymphomas NEC spleen
C0153858|ICD9CM|HT|202.9|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue
C0153859|ICD9CM|PT|202.91|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue, lymph nodes of head, face, and neck
C0153859|ICD9CM|AB|202.91|Lymphoid mal NEC head
C0153860|ICD9CM|PT|202.92|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue, intrathoracic lymph nodes
C0153860|ICD9CM|AB|202.92|Lymphoid mal NEC thorax
C0153861|ICD9CM|PT|202.93|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue, intra-abdominal lymph nodes
C0153861|ICD9CM|AB|202.93|Lymphoid mal NEC abdom
C0153862|ICD9CM|PT|202.94|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue, lymph nodes of axilla and upper limb
C0153862|ICD9CM|AB|202.94|Lymphoid mal NEC axilla
C0153863|ICD9CM|PT|202.95|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue, lymph nodes of inguinal region and lower limb
C0153863|ICD9CM|AB|202.95|Lymphoid mal NEC inguin
C0153864|ICD9CM|PT|202.96|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue, intrapelvic lymph nodes
C0153864|ICD9CM|AB|202.96|Lymphoid mal NEC pelvic
C0153865|ICD9CM|PT|202.97|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue, spleen
C0153865|ICD9CM|AB|202.97|Lymphoid mal NEC spleen
C0153866|ICD9CM|PT|202.98|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue, lymph nodes of multiple sites
C0153866|ICD9CM|AB|202.98|Lymphoid mal NEC mult
C0153867|ICD9CM|HT|203|Multiple myeloma and immunoproliferative neoplasms
C0153869|ICD9CM|PT|203.01|Multiple myeloma, in remission
C0153869|ICD9CM|AB|203.01|Mult myelm w remission
C0153871|ICD9CM|PT|203.11|Plasma cell leukemia, in remission
C0153871|ICD9CM|AB|203.11|Plsm cell leuk w rmson
C0153872|ICD9CM|HT|203.8|Other immunoproliferative neoplasms
C0153874|ICD9CM|PT|203.81|Other immunoproliferative neoplasms, in remission
C0153874|ICD9CM|AB|203.81|Oth imnprfl npl w rmsn
C0153876|ICD9CM|PT|204.01|Acute lymphoid leukemia, in remission
C0153876|ICD9CM|AB|204.01|Act lym leuk w rmsion
C0153878|ICD9CM|PT|204.11|Chronic lymphoid leukemia, in remission
C0153878|ICD9CM|AB|204.11|Chr lym leuk w rmsion
C0153880|ICD9CM|PT|204.21|Subacute lymphoid leukemia, in remission
C0153880|ICD9CM|AB|204.21|Sbac lym leuk w rmsion
C0153882|ICD9CM|PT|204.81|Other lymphoid leukemia, in remission
C0153882|ICD9CM|AB|204.81|Oth lym leuk w rmsion
C0153886|ICD9CM|PT|205.01|Acute myeloid leukemia, in remission
C0153886|ICD9CM|AB|205.01|Act myl leuk w rmsion
C0153888|ICD9CM|PT|205.11|Chronic myeloid leukemia, in remission
C0153888|ICD9CM|AB|205.11|Chr myl leuk w rmsion
C0153890|ICD9CM|PT|205.21|Subacute myeloid leukemia,in remission
C0153890|ICD9CM|AB|205.21|Sbac myl leuk w rmsion
C0153892|ICD9CM|PT|205.31|Myeloid sarcoma, in remission
C0153892|ICD9CM|AB|205.31|Myl srcoma w rmsion
C0153894|ICD9CM|PT|205.81|Other myeloid leukemia, in remission
C0153894|ICD9CM|AB|205.81|Oth myl leuk w rmsion
C0153898|ICD9CM|PT|206.01|Acute monocytic leukemia,in remission
C0153898|ICD9CM|AB|206.01|Act mono leuk w rmsion
C0153900|ICD9CM|PT|206.11|Chronic monocytic leukemia, in remission
C0153900|ICD9CM|AB|206.11|Chr mono leuk w rmsion
C0153902|ICD9CM|PT|206.21|Subacute monocytic leukemia, in remission
C0153902|ICD9CM|AB|206.21|Sbac mono leuk w rmsion
C0153903|ICD9CM|HT|206.8|Other monocytic leukemia
C0153905|ICD9CM|PT|206.81|Other monocytic leukemia, in remission
C0153905|ICD9CM|AB|206.81|Oth mono leuk w rmsion
C0153910|ICD9CM|PT|207.01|Acute erythremia and erythroleukemia, in remission
C0153910|ICD9CM|AB|207.01|Act erth/erylk w rmson
C0153912|ICD9CM|PT|207.11|Chronic erythremia, in remission
C0153912|ICD9CM|AB|207.11|Chr erythrm w remision
C0153914|ICD9CM|PT|207.21|Megakaryocytic leukemia, in remission
C0153914|ICD9CM|AB|207.21|Mgkrycyt leuk w rmsion
C0153916|ICD9CM|PT|207.81|Other specified leukemia, in remission
C0153916|ICD9CM|AB|207.81|Oth spf leuk w remsion
C0153924|ICD9CM|HT|208.2|Leukemia of unspecified cell type, subacute
C0153928|ICD9CM|PT|208.81|Other leukemia of unspecified cell type, in remission
C0153928|ICD9CM|AB|208.81|Oth leuk uns cl w rmson
C0153931|ICD9CM|HT|210|Benign neoplasm of lip, oral cavity, and pharynx
C0153932|ICD9CM|PT|210.0|Benign neoplasm of lip
C0153932|ICD9CM|AB|210.0|Benign neoplasm lip
C0153933|ICD9CM|PT|210.1|Benign neoplasm of tongue
C0153933|ICD9CM|AB|210.1|Benign neoplasm tongue
C0153934|ICD9CM|PT|210.3|Benign neoplasm of floor of mouth
C0153934|ICD9CM|AB|210.3|Benign neo mouth floor
C0153935|ICD9CM|PT|210.4|Benign neoplasm of other and unspecified parts of mouth
C0153935|ICD9CM|AB|210.4|Benign neo mouth NEC/NOS
C0153936|ICD9CM|PT|210.5|Benign neoplasm of tonsil
C0153936|ICD9CM|AB|210.5|Benign neoplasm tonsil
C0153937|ICD9CM|PT|210.6|Benign neoplasm of other parts of oropharynx
C0153937|ICD9CM|AB|210.6|Benign neo oropharyn NEC
C0153938|ICD9CM|PT|210.7|Benign neoplasm of nasopharynx
C0153938|ICD9CM|AB|210.7|Benign neo nasopharynx
C0153939|ICD9CM|PT|210.8|Benign neoplasm of hypopharynx
C0153939|ICD9CM|AB|210.8|Benign neo hypopharynx
C0153940|ICD9CM|PT|210.9|Benign neoplasm of pharynx, unspecified
C0153940|ICD9CM|AB|210.9|Benign neo pharynx NOS
C0153942|ICD9CM|PT|211.0|Benign neoplasm of esophagus
C0153942|ICD9CM|AB|211.0|Benign neo esophagus
C0153943|ICD9CM|PT|211.1|Benign neoplasm of stomach
C0153943|ICD9CM|AB|211.1|Benign neoplasm stomach
C0153944|ICD9CM|PT|211.2|Benign neoplasm of duodenum, jejunum, and ileum
C0153944|ICD9CM|AB|211.2|Benign neoplasm sm bowel
C0153945|ICD9CM|PT|211.4|Benign neoplasm of rectum and anal canal
C0153945|ICD9CM|AB|211.4|Benign neopl rectum/anus
C0153951|ICD9CM|PT|212.0|Benign neoplasm of nasal cavities, middle ear, and accessory sinuses
C0153951|ICD9CM|AB|212.0|Ben neo nasal cav/sinus
C0153952|ICD9CM|PT|212.1|Benign neoplasm of larynx
C0153952|ICD9CM|AB|212.1|Benign neo larynx
C0153953|ICD9CM|PT|212.2|Benign neoplasm of trachea
C0153953|ICD9CM|AB|212.2|Benign neo trachea
C0153954|ICD9CM|PT|212.3|Benign neoplasm of bronchus and lung
C0153954|ICD9CM|AB|212.3|Benign neo bronchus/lung
C0153955|ICD9CM|PT|212.4|Benign neoplasm of pleura
C0153955|ICD9CM|AB|212.4|Benign neoplasm pleura
C0153956|ICD9CM|PT|212.5|Benign neoplasm of mediastinum
C0153956|ICD9CM|AB|212.5|Benign neo mediastinum
C0153957|ICD9CM|PT|212.7|Benign neoplasm of heart
C0153957|ICD9CM|AB|212.7|Benign neoplasm heart
C0153958|ICD9CM|PT|212.8|Benign neoplasm of other specified sites of respiratory and intrathoracic organs
C0153958|ICD9CM|AB|212.8|Benign neo resp sys NEC
C0153959|ICD9CM|HT|213|Benign neoplasm of bone and articular cartilage
C0153959|ICD9CM|PT|213.9|Benign neoplasm of bone and articular cartilage, site unspecified
C0153959|ICD9CM|AB|213.9|Benign neo bone NOS
C0153960|ICD9CM|PT|213.0|Benign neoplasm of bones of skull and face
C0153960|ICD9CM|AB|213.0|Ben neo skull/face bone
C0153962|ICD9CM|PT|213.3|Benign neoplasm of ribs, sternum, and clavicle
C0153962|ICD9CM|AB|213.3|Ben neo ribs/stern/clav
C0153963|ICD9CM|PT|213.4|Benign neoplasm of scapula and long bones of upper limb
C0153963|ICD9CM|AB|213.4|Ben neo long bones arm
C0153964|ICD9CM|PT|213.5|Benign neoplasm of short bones of upper limb
C0153964|ICD9CM|AB|213.5|Ben neo bones wrist/hand
C0153965|ICD9CM|PT|213.6|Benign neoplasm of pelvic bones, sacrum, and coccyx
C0153965|ICD9CM|AB|213.6|Benign neo pelvic girdle
C0153966|ICD9CM|PT|213.7|Benign neoplasm of long bones of lower limb
C0153966|ICD9CM|AB|213.7|Ben neo long bones leg
C0153967|ICD9CM|PT|213.8|Benign neoplasm of short bones of lower limb
C0153967|ICD9CM|AB|213.8|Ben neo bones ankle/foot
C0153968|ICD9CM|PT|214.0|Lipoma of skin and subcutaneous tissue of face
C0153968|ICD9CM|AB|214.0|Lipoma skin face
C0153969|ICD9CM|PT|214.1|Lipoma of other skin and subcutaneous tissue
C0153969|ICD9CM|AB|214.1|Lipoma skin NEC
C0153970|ICD9CM|PT|214.2|Lipoma of intrathoracic organs
C0153970|ICD9CM|AB|214.2|Lipoma intrathoracic
C0153971|ICD9CM|PT|214.3|Lipoma of intra-abdominal organs
C0153971|ICD9CM|AB|214.3|Lipoma intra-abdominal
C0153972|ICD9CM|PT|214.4|Lipoma of spermatic cord
C0153972|ICD9CM|AB|214.4|Lipoma spermatic cord
C0153974|ICD9CM|PT|215.0|Other benign neoplasm of connective and other soft tissue of head, face, and neck
C0153974|ICD9CM|AB|215.0|Ben neo soft tissue head
C0153975|ICD9CM|PT|215.2|Other benign neoplasm of connective and other soft tissue of upper limb, including shoulder
C0153975|ICD9CM|AB|215.2|Ben neo soft tissue arm
C0153976|ICD9CM|PT|215.3|Other benign neoplasm of connective and other soft tissue of lower limb, including hip
C0153976|ICD9CM|AB|215.3|Ben neo soft tissue leg
C0153977|ICD9CM|PT|215.4|Other benign neoplasm of connective and other soft tissue of thorax
C0153977|ICD9CM|AB|215.4|Ben neo soft tis thorax
C0153978|ICD9CM|PT|215.5|Other benign neoplasm of connective and other soft tissue of abdomen
C0153978|ICD9CM|AB|215.5|Ben neo soft tis abdomen
C0153979|ICD9CM|PT|215.6|Other benign neoplasm of connective and other soft tissue of pelvis
C0153979|ICD9CM|AB|215.6|Ben neo soft tis pelvis
C0153981|ICD9CM|PT|215.8|Other benign neoplasm of connective and other soft tissue of other specified sites
C0153981|ICD9CM|AB|215.8|Ben neo soft tissue NEC
C0153982|ICD9CM|PT|216.0|Benign neoplasm of skin of lip
C0153982|ICD9CM|AB|216.0|Benign neo skin lip
C0153983|ICD9CM|PT|216.1|Benign neoplasm of eyelid, including canthus
C0153983|ICD9CM|AB|216.1|Benign neo skin eyelid
C0153984|ICD9CM|PT|216.2|Benign neoplasm of ear and external auditory canal
C0153984|ICD9CM|AB|216.2|Benign neo skin ear
C0153985|ICD9CM|PT|216.3|Benign neoplasm of skin of other and unspecified parts of face
C0153985|ICD9CM|AB|216.3|Benign neo skin face NEC
C0153986|ICD9CM|PT|216.4|Benign neoplasm of scalp and skin of neck
C0153986|ICD9CM|AB|216.4|Ben neo scalp/skin neck
C0153987|ICD9CM|PT|216.5|Benign neoplasm of skin of trunk, except scrotum
C0153987|ICD9CM|AB|216.5|Benign neo skin trunk
C0153988|ICD9CM|PT|216.6|Benign neoplasm of skin of upper limb, including shoulder
C0153988|ICD9CM|AB|216.6|Benign neo skin arm
C0153989|ICD9CM|PT|216.7|Benign neoplasm of skin of lower limb, including hip
C0153989|ICD9CM|AB|216.7|Benign neo skin leg
C0153990|ICD9CM|PT|216.8|Benign neoplasm of other specified sites of skin
C0153990|ICD9CM|AB|216.8|Benign neoplasm skin NEC
C0153993|ICD9CM|PT|218.0|Submucous leiomyoma of uterus
C0153993|ICD9CM|AB|218.0|Submucous leiomyoma
C0153994|ICD9CM|PT|218.1|Intramural leiomyoma of uterus
C0153994|ICD9CM|AB|218.1|Intramural leiomyoma
C0153995|ICD9CM|PT|218.2|Subserous leiomyoma of uterus
C0153995|ICD9CM|AB|218.2|Subserous leiomyoma
C0153996|ICD9CM|HT|219|Other benign neoplasm of uterus
C0153997|ICD9CM|PT|219.0|Benign neoplasm of cervix uteri
C0153997|ICD9CM|AB|219.0|Benign neo cervix uteri
C0153998|ICD9CM|PT|219.1|Benign neoplasm of corpus uteri
C0153998|ICD9CM|AB|219.1|Benign neo corpus uteri
C0153999|ICD9CM|PT|219.9|Benign neoplasm of uterus, part unspecified
C0153999|ICD9CM|AB|219.9|Benign neo uterus NOS
C0154000|ICD9CM|HT|221|Benign neoplasm of other female genital organs
C0154002|ICD9CM|AB|221.1|Benign neoplasm vagina
C0154002|ICD9CM|PT|221.1|Benign neoplasm of vagina
C0154003|ICD9CM|PT|221.2|Benign neoplasm of vulva
C0154003|ICD9CM|AB|221.2|Benign neoplasm vulva
C0154004|ICD9CM|PT|221.8|Benign neoplasm of other specified sites of female genital organs
C0154004|ICD9CM|AB|221.8|Ben neo fem genital NEC
C0154005|ICD9CM|PT|221.9|Benign neoplasm of female genital organ, site unspecified
C0154005|ICD9CM|AB|221.9|Ben neo fem genital NOS
C0154007|ICD9CM|PT|222.0|Benign neoplasm of testis
C0154007|ICD9CM|AB|222.0|Benign neoplasm testis
C0154009|ICD9CM|PT|222.2|Benign neoplasm of prostate
C0154009|ICD9CM|AB|222.2|Benign neoplasm prostate
C0154010|ICD9CM|PT|222.3|Benign neoplasm of epididymis
C0154010|ICD9CM|AB|222.3|Benign neo epididymis
C0154011|ICD9CM|PT|222.4|Benign neoplasm of scrotum
C0154011|ICD9CM|AB|222.4|Benign neoplasm scrotum
C0154012|ICD9CM|PT|222.8|Benign neoplasm of other specified sites of male genital organs
C0154012|ICD9CM|AB|222.8|Ben neo male genital NEC
C0154013|ICD9CM|HT|223|Benign neoplasm of kidney and other urinary organs
C0154014|ICD9CM|PT|223.0|Benign neoplasm of kidney, except pelvis
C0154014|ICD9CM|AB|223.0|Benign neoplasm kidney
C0154015|ICD9CM|PT|223.1|Benign neoplasm of renal pelvis
C0154015|ICD9CM|AB|223.1|Benign neo renal pelvis
C0154016|ICD9CM|PT|223.2|Benign neoplasm of ureter
C0154016|ICD9CM|AB|223.2|Benign neoplasm ureter
C0154017|ICD9CM|PT|223.3|Benign neoplasm of bladder
C0154017|ICD9CM|AB|223.3|Benign neoplasm bladder
C0154018|ICD9CM|HT|223.8|Benign neoplasm of other specified sites of urinary organs
C0154018|ICD9CM|PT|223.89|Benign neoplasm of other specified sites of urinary organs
C0154018|ICD9CM|AB|223.89|Benign neo urinary NEC
C0154019|ICD9CM|PT|223.81|Benign neoplasm of urethra
C0154019|ICD9CM|AB|223.81|Benign neoplasm urethra
C0154022|ICD9CM|PT|224.0|Benign neoplasm of eyeball, except conjunctiva, cornea, retina, and choroid
C0154022|ICD9CM|AB|224.0|Benign neoplasm eyeball
C0154023|ICD9CM|PT|224.1|Benign neoplasm of orbit
C0154023|ICD9CM|AB|224.1|Benign neoplasm orbit
C0154024|ICD9CM|PT|224.2|Benign neoplasm of lacrimal gland
C0154024|ICD9CM|AB|224.2|Ben neo lacrimal gland
C0154025|ICD9CM|PT|224.3|Benign neoplasm of conjunctiva
C0154025|ICD9CM|AB|224.3|Benign neo conjunctiva
C0154026|ICD9CM|PT|224.4|Benign neoplasm of cornea
C0154026|ICD9CM|AB|224.4|Benign neoplasm cornea
C0154027|ICD9CM|PT|224.5|Benign neoplasm of retina
C0154027|ICD9CM|AB|224.5|Benign neoplasm retina
C0154028|ICD9CM|PT|224.6|Benign neoplasm of choroid
C0154028|ICD9CM|AB|224.6|Benign neoplasm choroid
C0154029|ICD9CM|PT|224.7|Benign neoplasm of lacrimal duct
C0154029|ICD9CM|AB|224.7|Ben neo lacrimal duct
C0154030|ICD9CM|PT|224.8|Benign neoplasm of other specified parts of eye
C0154030|ICD9CM|AB|224.8|Benign neoplasm eye NEC
C0154033|ICD9CM|PT|225.2|Benign neoplasm of cerebral meninges
C0154033|ICD9CM|AB|225.2|Ben neo cerebr meninges
C0154034|ICD9CM|PT|225.3|Benign neoplasm of spinal cord
C0154034|ICD9CM|AB|225.3|Benign neo spinal cord
C0154035|ICD9CM|PT|225.4|Benign neoplasm of spinal meninges
C0154035|ICD9CM|AB|225.4|Ben neo spinal meninges
C0154036|ICD9CM|PT|225.8|Benign neoplasm of other specified sites of nervous system
C0154036|ICD9CM|AB|225.8|Benign neo nerv sys NEC
C0154038|ICD9CM|PT|226|Benign neoplasm of thyroid glands
C0154038|ICD9CM|AB|226|Benign neoplasm thyroid
C0154039|ICD9CM|HT|227|Benign neoplasm of other endocrine glands and related structures
C0154039|ICD9CM|PT|227.8|Benign neoplasm of other endocrine glands and related structures
C0154039|ICD9CM|AB|227.8|Benign neo endocrine NEC
C0154040|ICD9CM|PT|227.0|Benign neoplasm of adrenal gland
C0154040|ICD9CM|AB|227.0|Benign neoplasm adrenal
C0154041|ICD9CM|PT|227.1|Benign neoplasm of parathyroid gland
C0154041|ICD9CM|AB|227.1|Benign neo parathyroid
C0154043|ICD9CM|PT|227.4|Benign neoplasm of pineal gland
C0154043|ICD9CM|AB|227.4|Ben neopl pineal gland
C0154044|ICD9CM|PT|227.5|Benign neoplasm of carotid body
C0154044|ICD9CM|AB|227.5|Benign neo carotid body
C0154045|ICD9CM|PT|227.6|Benign neoplasm of aortic body and other paraganglia
C0154045|ICD9CM|AB|227.6|Ben neo paraganglia NEC
C0154049|ICD9CM|PT|228.01|Hemangioma of skin and subcutaneous tissue
C0154049|ICD9CM|AB|228.01|Hemangioma skin
C0154050|ICD9CM|PT|228.02|Hemangioma of intracranial structures
C0154050|ICD9CM|AB|228.02|Hemangioma intracranial
C0154051|ICD9CM|PT|228.03|Hemangioma of retina
C0154051|ICD9CM|AB|228.03|Hemangioma retina
C0154052|ICD9CM|PT|228.04|Hemangioma of intra-abdominal structures
C0154052|ICD9CM|AB|228.04|Hemangioma intra-abdom
C0154053|ICD9CM|HT|229|Benign neoplasm of other and unspecified sites
C0154054|ICD9CM|PT|229.0|Benign neoplasm of lymph nodes
C0154054|ICD9CM|AB|229.0|Benign neo lymph nodes
C0154055|ICD9CM|PT|229.8|Benign neoplasm of other specified sites
C0154055|ICD9CM|AB|229.8|Benign neoplasm NEC
C0154057|ICD9CM|HT|230|Carcinoma in situ of digestive organs
C0154058|ICD9CM|PT|230.0|Carcinoma in situ of lip, oral cavity, and pharynx
C0154058|ICD9CM|AB|230.0|Ca in situ oral cav/phar
C0154059|ICD9CM|PT|230.1|Carcinoma in situ of esophagus
C0154059|ICD9CM|AB|230.1|Ca in situ esophagus
C0154060|ICD9CM|PT|230.2|Carcinoma in situ of stomach
C0154060|ICD9CM|AB|230.2|Ca in situ stomach
C0154061|ICD9CM|PT|230.3|Carcinoma in situ of colon
C0154061|ICD9CM|AB|230.3|Ca in situ colon
C0154062|ICD9CM|PT|230.4|Carcinoma in situ of rectum
C0154062|ICD9CM|AB|230.4|Ca in situ rectum
C0154064|ICD9CM|PT|230.6|Carcinoma in situ of anus, unspecified
C0154064|ICD9CM|AB|230.6|Ca in situ anus NOS
C0154065|ICD9CM|PT|230.7|Carcinoma in situ of other and unspecified parts of intestine
C0154065|ICD9CM|AB|230.7|Ca in situ bowel NEC/NOS
C0154067|ICD9CM|PT|230.9|Carcinoma in situ of other and unspecified digestive organs
C0154067|ICD9CM|AB|230.9|Ca in situ GI NEC/NOS
C0154069|ICD9CM|PT|231.0|Carcinoma in situ of larynx
C0154069|ICD9CM|AB|231.0|Ca in situ larynx
C0154070|ICD9CM|PT|231.1|Carcinoma in situ of trachea
C0154070|ICD9CM|AB|231.1|Ca in situ trachea
C0154071|ICD9CM|PT|231.2|Carcinoma in situ of bronchus and lung
C0154071|ICD9CM|AB|231.2|Ca in situ bronchus/lung
C0154072|ICD9CM|PT|231.8|Carcinoma in situ of other specified parts of respiratory system
C0154072|ICD9CM|AB|231.8|Ca in situ resp sys NEC
C0154073|ICD9CM|HT|232|Carcinoma in situ of skin
C0154073|ICD9CM|PT|232.9|Carcinoma in situ of skin, site unspecified
C0154073|ICD9CM|AB|232.9|Ca in situ skin NOS
C0154074|ICD9CM|PT|232.0|Carcinoma in situ of skin of lip
C0154074|ICD9CM|AB|232.0|Ca in situ skin lip
C0154077|ICD9CM|PT|232.3|Carcinoma in situ of skin of other and unspecified parts of face
C0154077|ICD9CM|AB|232.3|Ca in situ skin face NEC
C0154078|ICD9CM|PT|232.4|Carcinoma in situ of scalp and skin of neck
C0154078|ICD9CM|AB|232.4|Ca in situ scalp
C0154079|ICD9CM|PT|232.5|Carcinoma in situ of skin of trunk, except scrotum
C0154079|ICD9CM|AB|232.5|Ca in situ skin trunk
C0154080|ICD9CM|PT|232.6|Carcinoma in situ of skin of upper limb, including shoulder
C0154080|ICD9CM|AB|232.6|Ca in situ skin arm
C0154081|ICD9CM|PT|232.7|Carcinoma in situ of skin of lower limb, including hip
C0154081|ICD9CM|AB|232.7|Ca in situ skin leg
C0154082|ICD9CM|PT|232.8|Carcinoma in situ of other specified sites of skin
C0154082|ICD9CM|AB|232.8|Ca in situ skin NEC
C0154083|ICD9CM|HT|233|Carcinoma in situ of breast and genitourinary system
C0154084|ICD9CM|PT|233.0|Carcinoma in situ of breast
C0154084|ICD9CM|AB|233.0|Ca in situ breast
C0154086|ICD9CM|PT|233.2|Carcinoma in situ of other and unspecified parts of uterus
C0154086|ICD9CM|AB|233.2|Ca in situ uterus NEC
C0154087|ICD9CM|HT|233.3|Carcinoma in situ of other and unspecified female genital organs
C0154088|ICD9CM|PT|233.4|Carcinoma in situ of prostate
C0154088|ICD9CM|AB|233.4|Ca in situ prostate
C0154089|ICD9CM|PT|233.5|Carcinoma in situ of penis
C0154089|ICD9CM|AB|233.5|Ca in situ penis
C0154090|ICD9CM|PT|233.6|Carcinoma in situ of other and unspecified male genital organs
C0154090|ICD9CM|AB|233.6|Ca in situ male gen NEC
C0154091|ICD9CM|PT|233.7|Carcinoma in situ of bladder
C0154091|ICD9CM|AB|233.7|Ca in situ bladder
C0154092|ICD9CM|PT|233.9|Carcinoma in situ of other and unspecified urinary organs
C0154092|ICD9CM|AB|233.9|Ca in situ urinary NEC
C0154093|ICD9CM|HT|234|Carcinoma in situ of other and unspecified sites
C0154094|ICD9CM|PT|234.0|Carcinoma in situ of eye
C0154094|ICD9CM|AB|234.0|Ca in situ eye
C0154095|ICD9CM|HT|235|Neoplasm of uncertain behavior of digestive and respiratory systems
C0154096|ICD9CM|PT|235.0|Neoplasm of uncertain behavior of major salivary glands
C0154096|ICD9CM|AB|235.0|Unc behav neo salivary
C0154097|ICD9CM|PT|235.1|Neoplasm of uncertain behavior of lip, oral cavity, and pharynx
C0154097|ICD9CM|AB|235.1|Unc behav neo oral/phar
C0154098|ICD9CM|PT|235.2|Neoplasm of uncertain behavior of stomach, intestines, and rectum
C0154098|ICD9CM|AB|235.2|Unc behav neo intestine
C0154100|ICD9CM|PT|235.4|Neoplasm of uncertain behavior of retroperitoneum and peritoneum
C0154100|ICD9CM|AB|235.4|Unc behav neo peritoneum
C0154101|ICD9CM|PT|235.5|Neoplasm of uncertain behavior of other and unspecified digestive organs
C0154101|ICD9CM|AB|235.5|Unc behav neo GI NEC
C0154103|ICD9CM|PT|235.7|Neoplasm of uncertain behavior of trachea, bronchus, and lung
C0154103|ICD9CM|AB|235.7|Unc behav neo lung
C0154104|ICD9CM|PT|235.8|Neoplasm of uncertain behavior of pleura, thymus, and mediastinum
C0154104|ICD9CM|AB|235.8|Unc behav neo pleura
C0154105|ICD9CM|PT|235.9|Neoplasm of uncertain behavior of other and unspecified respiratory organs
C0154105|ICD9CM|AB|235.9|Unc behav neo resp NEC
C0154106|ICD9CM|HT|236|Neoplasm of uncertain behavior of genitourinary organs
C0154113|ICD9CM|HT|236.9|Neoplasm of uncertain behavior of other and unspecified urinary organs
C0154115|ICD9CM|PT|236.91|Neoplasm of uncertain behavior of kidney and ureter
C0154115|ICD9CM|AB|236.91|Unc behav neo kidney
C0154116|ICD9CM|HT|237|Neoplasm of uncertain behavior of endocrine glands and nervous system
C0154117|ICD9CM|PT|237.2|Neoplasm of uncertain behavior of adrenal gland
C0154117|ICD9CM|AB|237.2|Unc behav neo adrenal
C0154118|ICD9CM|PT|237.4|Neoplasm of uncertain behavior of other and unspecified endocrine glands
C0154118|ICD9CM|AB|237.4|Uncer neo endocrine NEC
C0154119|ICD9CM|PT|237.5|Neoplasm of uncertain behavior of brain and spinal cord
C0154119|ICD9CM|AB|237.5|Unc beh neo brain/spinal
C0154120|ICD9CM|PT|237.6|Neoplasm of uncertain behavior of meninges
C0154120|ICD9CM|AB|237.6|Unc behav neo meninges
C0154123|ICD9CM|PT|237.9|Neoplasm of uncertain behavior of other and unspecified parts of nervous system
C0154123|ICD9CM|AB|237.9|Unc beh neo nerv sys NEC
C0154124|ICD9CM|HT|238|Neoplasm of uncertain behavior of other and unspecified sites and tissues
C0154125|ICD9CM|PT|238.1|Neoplasm of uncertain behavior of connective and other soft tissue
C0154125|ICD9CM|AB|238.1|Unc behav neo soft tissu
C0154127|ICD9CM|PT|238.5|Neoplasm of uncertain behavior of histiocytic and mast cells
C0154127|ICD9CM|AB|238.5|Mastocytoma NOS
C0154129|ICD9CM|HT|235-238.99|NEOPLASMS OF UNCERTAIN BEHAVIOR
C0154131|ICD9CM|PT|239.1|Neoplasm of unspecified nature of respiratory system
C0154131|ICD9CM|AB|239.1|Respiratory neoplasm NOS
C0154132|ICD9CM|PT|239.2|Neoplasm of unspecified nature of bone, soft tissue, and skin
C0154132|ICD9CM|AB|239.2|Bone/skin neoplasm NOS
C0154133|ICD9CM|PT|239.5|Neoplasm of unspecified nature of other genitourinary organs
C0154133|ICD9CM|AB|239.5|Other gu neoplasm NOS
C0154134|ICD9CM|PT|239.7|Neoplasm of unspecified nature of endocrine glands and other parts of nervous system
C0154134|ICD9CM|AB|239.7|Endocrine/nerv neo NOS
C0154135|ICD9CM|HT|239.8|Neoplasm of unspecified nature of other specified sites
C0154135|ICD9CM|PT|239.89|Neoplasms of unspecified nature, other specified sites
C0154135|ICD9CM|AB|239.89|Neoplasm other sites NOS
C0154138|ICD9CM|PT|242.00|Toxic diffuse goiter without mention of thyrotoxic crisis or storm
C0154138|ICD9CM|AB|242.00|Tox dif goiter no crisis
C0154139|ICD9CM|PT|242.01|Toxic diffuse goiter with mention of thyrotoxic crisis or storm
C0154139|ICD9CM|AB|242.01|Tox dif goiter w crisis
C0154141|ICD9CM|HT|242.1|Toxic uninodular goiter
C0154142|ICD9CM|PT|242.11|Toxic uninodular goiter with mention of thyrotoxic crisis or storm
C0154142|ICD9CM|AB|242.11|Tox uninod goit w crisis
C0154143|ICD9CM|HT|242.2|Toxic multinodular goiter
C0154144|ICD9CM|PT|242.20|Toxic multinodular goiter without mention of thyrotoxic crisis or storm
C0154144|ICD9CM|AB|242.20|Tox multnod goit no cris
C0154145|ICD9CM|PT|242.21|Toxic multinodular goiter with mention of thyrotoxic crisis or storm
C0154145|ICD9CM|AB|242.21|Tox multnod goit w cris
C0154146|ICD9CM|PT|242.30|Toxic nodular goiter, unspecified type, without mention of thyrotoxic crisis or storm
C0154146|ICD9CM|AB|242.30|Tox nod goiter no crisis
C0154147|ICD9CM|PT|242.31|Toxic nodular goiter, unspecified type, with mention of thyrotoxic crisis or storm
C0154147|ICD9CM|AB|242.31|Tox nod goiter w crisis
C0154148|ICD9CM|HT|242.4|Thyrotoxicosis from ectopic thyroid nodule
C0154151|ICD9CM|HT|242.8|Thyrotoxicosis of other specified origin
C0154152|ICD9CM|PT|242.80|Thyrotoxicosis of other specified origin without mention of thyrotoxic crisis or storm
C0154152|ICD9CM|AB|242.80|Thyrtox orig NEC no cris
C0154153|ICD9CM|PT|242.81|Thyrotoxicosis of other specified origin with mention of thyrotoxic crisis or storm
C0154153|ICD9CM|AB|242.81|Thyrotox orig NEC w cris
C0154154|ICD9CM|PT|242.90|Thyrotoxicosis without mention of goiter or other cause, and without mention of thyrotoxic crisis or storm
C0154154|ICD9CM|AB|242.90|Thyrotox NOS no crisis
C0154155|ICD9CM|PT|242.91|Thyrotoxicosis without mention of goiter or other cause, with mention of thyrotoxic crisis or storm
C0154155|ICD9CM|AB|242.91|Thyrotox NOS w crisis
C0154157|ICD9CM|PT|244.0|Postsurgical hypothyroidism
C0154157|ICD9CM|AB|244.0|Postsurgical hypothyroid
C0154158|ICD9CM|PT|244.1|Other postablative hypothyroidism
C0154158|ICD9CM|AB|244.1|Postablat hypothyr NEC
C0154159|ICD9CM|AB|244.2|Iodine hypothyroidism
C0154159|ICD9CM|PT|244.2|Iodine hypothyroidism
C0154160|ICD9CM|PT|244.3|Other iatrogenic hypothyroidism
C0154160|ICD9CM|AB|244.3|Iatrogen hypothyroid NEC
C0154161|ICD9CM|PT|244.8|Other specified acquired hypothyroidism
C0154161|ICD9CM|AB|244.8|Acquired hypothyroid NEC
C0154163|ICD9CM|AB|245.4|Iatrogenic thyroiditis
C0154163|ICD9CM|PT|245.4|Iatrogenic thyroiditis
C0154164|ICD9CM|HT|246|Other disorders of thyroid
C0154166|ICD9CM|PT|246.3|Hemorrhage and infarction of thyroid
C0154166|ICD9CM|AB|246.3|Hemorr/infarc thyroid
C0154167|ICD9CM|PT|246.8|Other specified disorders of thyroid
C0154167|ICD9CM|AB|246.8|Disorders of thyroid NEC
C0154183|ICD9CM|HT|250.8|Diabetes with other specified manifestations
C0154189|ICD9CM|HT|251|Other disorders of pancreatic internal secretion
C0154190|ICD9CM|PT|251.3|Postsurgical hypoinsulinemia
C0154190|ICD9CM|AB|251.3|Postsurg hypoinsulinemia
C0154191|ICD9CM|PT|251.4|Abnormality of secretion of glucagon
C0154191|ICD9CM|AB|251.4|Abn secretion glucagon
C0154192|ICD9CM|PT|251.8|Other specified disorders of pancreatic internal secretion
C0154192|ICD9CM|AB|251.8|Pancreatic disorder NEC
C0154195|ICD9CM|PT|252.8|Other specified disorders of parathyroid gland
C0154195|ICD9CM|AB|252.8|Parathyroid disorder NEC
C0154198|ICD9CM|PT|253.7|Iatrogenic pituitary disorders
C0154198|ICD9CM|AB|253.7|Iatrogenic pituitary dis
C0154199|ICD9CM|HT|254|Diseases of thymus gland
C0154199|ICD9CM|PT|254.9|Unspecified disease of thymus gland
C0154199|ICD9CM|AB|254.9|Disease of thymus NOS
C0154200|ICD9CM|AB|254.1|Abscess of thymus
C0154200|ICD9CM|PT|254.1|Abscess of thymus
C0154205|ICD9CM|PT|255.5|Other adrenal hypofunction
C0154205|ICD9CM|AB|255.5|Adrenal hypofunction NEC
C0154206|ICD9CM|PT|255.6|Medulloadrenal hyperfunction
C0154206|ICD9CM|AB|255.6|Medulloadrenal hyperfunc
C0154207|ICD9CM|PT|255.8|Other specified disorders of adrenal glands
C0154207|ICD9CM|AB|255.8|Adrenal disorder NEC
C0154208|ICD9CM|HT|256|Ovarian dysfunction
C0154208|ICD9CM|AB|256.9|Ovarian dysfunction NOS
C0154208|ICD9CM|PT|256.9|Unspecified ovarian dysfunction
C0154209|ICD9CM|AB|256.0|Hyperestrogenism
C0154209|ICD9CM|PT|256.0|Hyperestrogenism
C0154210|ICD9CM|PT|256.1|Other ovarian hyperfunction
C0154210|ICD9CM|AB|256.1|Ovarian hyperfunc NEC
C0154211|ICD9CM|PT|256.2|Postablative ovarian failure
C0154211|ICD9CM|AB|256.2|Postablativ ovarian fail
C0154212|ICD9CM|PT|256.8|Other ovarian dysfunction
C0154212|ICD9CM|AB|256.8|Ovarian dysfunction NEC
C0154215|ICD9CM|AB|257.0|Testicular hyperfunction
C0154215|ICD9CM|PT|257.0|Testicular hyperfunction
C0154216|ICD9CM|PT|257.1|Postablative testicular hypofunction
C0154216|ICD9CM|AB|257.1|Postablat testic hypofun
C0154218|ICD9CM|HT|258|Polyglandular dysfunction and related disorders
C0154220|ICD9CM|PT|258.1|Other combinations of endocrine dysfunction
C0154220|ICD9CM|AB|258.1|Comb endocr dysfunct NEC
C0154221|ICD9CM|PT|258.8|Other specified polyglandular dysfunction
C0154221|ICD9CM|AB|258.8|Polyglandul dysfunc NEC
C0154222|ICD9CM|PT|258.9|Polyglandular dysfunction, unspecified
C0154222|ICD9CM|AB|258.9|Polyglandul dysfunc NOS
C0154223|ICD9CM|HT|259|Other endocrine disorders
C0154227|ICD9CM|PT|263.0|Malnutrition of moderate degree
C0154227|ICD9CM|AB|263.0|Malnutrition mod degree
C0154228|ICD9CM|AB|263.1|Malnutrition mild degree
C0154228|ICD9CM|PT|263.1|Malnutrition of mild degree
C0154229|ICD9CM|PT|263.2|Arrested development following protein-calorie malnutrition
C0154229|ICD9CM|AB|263.2|Arrest devel d/t malnutr
C0154230|ICD9CM|PT|263.8|Other protein-calorie malnutrition
C0154230|ICD9CM|AB|263.8|Protein-cal malnutr NEC
C0154231|ICD9CM|PT|264.0|Vitamin A deficiency with conjunctival xerosis
C0154231|ICD9CM|AB|264.0|Vit A conjunctiv xerosis
C0154232|ICD9CM|PT|264.1|Vitamin A deficiency with conjunctival xerosis and Bitot's spot
C0154232|ICD9CM|AB|264.1|Vit A bitot's spot
C0154233|ICD9CM|PT|264.2|Vitamin A deficiency with corneal xerosis
C0154233|ICD9CM|AB|264.2|Vit A corneal xerosis
C0154234|ICD9CM|PT|264.3|Vitamin A deficiency with corneal ulceration and xerosis
C0154234|ICD9CM|AB|264.3|Vit A cornea ulcer/xeros
C0154235|ICD9CM|PT|264.4|Vitamin A deficiency with keratomalacia
C0154235|ICD9CM|AB|264.4|Vit A keratomalacia
C0154236|ICD9CM|PT|264.5|Vitamin A deficiency with night blindness
C0154236|ICD9CM|AB|264.5|Vit A night blindness
C0154237|ICD9CM|PT|264.6|Vitamin A deficiency with xerophthalmic scars of cornea
C0154237|ICD9CM|AB|264.6|Vit A def w corneal scar
C0154238|ICD9CM|PT|264.7|Other ocular manifestations of vitamin A deficiency
C0154238|ICD9CM|AB|264.7|Vit A ocular defic NEC
C0154239|ICD9CM|HT|265|Thiamine and niacin deficiency states
C0154240|ICD9CM|AB|268.1|Rickets, late effect
C0154240|ICD9CM|PT|268.1|Rickets, late effect
C0154241|ICD9CM|PT|269.8|Other nutritional deficiency
C0154241|ICD9CM|HT|269|Other nutritional deficiencies
C0154241|ICD9CM|AB|269.8|Nutrition deficiency NEC
C0154246|ICD9CM|PT|270.6|Disorders of urea cycle metabolism
C0154246|ICD9CM|AB|270.6|Dis urea cycle metabol
C0154247|ICD9CM|PT|270.7|Other disturbances of straight-chain amino-acid metabolism
C0154247|ICD9CM|AB|270.7|Straig amin-acid met NEC
C0154249|ICD9CM|HT|271|Disorders of carbohydrate transport and metabolism
C0154249|ICD9CM|PT|271.9|Unspecified disorder of carbohydrate transport and metabolism
C0154249|ICD9CM|AB|271.9|Dis carbohydr metab NOS
C0154251|ICD9CM|HT|272|Disorders of lipoid metabolism
C0154251|ICD9CM|PT|272.9|Unspecified disorder of lipoid metabolism
C0154251|ICD9CM|AB|272.9|Lipoid metabol dis NOS
C0154254|ICD9CM|PT|273.0|Polyclonal hypergammaglobulinemia
C0154254|ICD9CM|AB|273.0|Polyclon hypergammaglobu
C0154256|ICD9CM|PT|274.19|Other gouty nephropathy
C0154256|ICD9CM|AB|274.19|Gouty nephropathy NEC
C0154257|ICD9CM|HT|274.8|Gout with other specified manifestations
C0154257|ICD9CM|PT|274.89|Gout with other specified manifestations
C0154257|ICD9CM|AB|274.89|Gout w manifestation NEC
C0154258|ICD9CM|AB|274.81|Gouty tophi of ear
C0154258|ICD9CM|PT|274.81|Gouty tophi of ear
C0154259|ICD9CM|PT|274.82|Gouty tophi of other sites, except ear
C0154259|ICD9CM|AB|274.82|Gouty tophi site NEC
C0154260|ICD9CM|HT|275|Disorders of mineral metabolism
C0154260|ICD9CM|PT|275.9|Unspecified disorder of mineral metabolism
C0154260|ICD9CM|AB|275.9|Dis mineral metabol NOS
C0154261|ICD9CM|PT|275.8|Other specified disorders of mineral metabolism
C0154261|ICD9CM|AB|275.8|Dis mineral metabol NEC
C0154264|ICD9CM|PT|276.4|Mixed acid-base balance disorder
C0154264|ICD9CM|AB|276.4|Mixed acid-base bal dis
C0154270|ICD9CM|AB|278.1|Localized adiposity
C0154270|ICD9CM|PT|278.1|Localized adiposity
C0154271|ICD9CM|AB|278.3|Hypercarotinemia
C0154271|ICD9CM|PT|278.3|Hypercarotinemia
C0154275|ICD9CM|PT|279.02|Selective IgM immunodeficiency
C0154275|ICD9CM|AB|279.02|Selective IgM immunodef
C0154276|ICD9CM|PT|279.03|Other selective immunoglobulin deficiencies
C0154276|ICD9CM|AB|279.03|Selective ig defic NEC
C0154282|ICD9CM|PT|279.19|Other deficiency of cell-mediated immunity
C0154282|ICD9CM|AB|279.19|Defic cell immunity NOS
C0154286|ICD9CM|PT|280.0|Iron deficiency anemia secondary to blood loss (chronic)
C0154286|ICD9CM|AB|280.0|Chr blood loss anemia
C0154287|ICD9CM|PT|280.1|Iron deficiency anemia secondary to inadequate dietary iron intake
C0154287|ICD9CM|AB|280.1|Iron def anemia dietary
C0154288|ICD9CM|HT|281|Other deficiency anemias
C0154289|ICD9CM|PT|281.1|Other vitamin B12 deficiency anemia
C0154289|ICD9CM|AB|281.1|B12 defic anemia NEC
C0154290|ICD9CM|PT|281.4|Protein-deficiency anemia
C0154290|ICD9CM|AB|281.4|Protein defic anemia
C0154291|ICD9CM|PT|281.8|Anemia associated with other specified nutritional deficiency
C0154291|ICD9CM|AB|281.8|Nutritional anemia NEC
C0154292|ICD9CM|PT|282.3|Other hemolytic anemias due to enzyme deficiency
C0154292|ICD9CM|AB|282.3|Enzyme defic anemia NEC
C0154296|ICD9CM|PT|282.8|Other specified hereditary hemolytic anemias
C0154296|ICD9CM|AB|282.8|Hered hemolytic anem NEC
C0154298|ICD9CM|PT|285.1|Acute posthemorrhagic anemia
C0154298|ICD9CM|AB|285.1|Ac posthemorrhag anemia
C0154300|ICD9CM|HT|287|Purpura and other hemorrhagic conditions
C0154301|ICD9CM|HT|287.4|Secondary thrombocytopenia
C0154304|ICD9CM|AB|289.1|Chronic lymphadenitis
C0154304|ICD9CM|PT|289.1|Chronic lymphadenitis
C0154305|ICD9CM|HT|289.5|Other diseases of spleen
C0154305|ICD9CM|PT|289.59|Other diseases of spleen
C0154305|ICD9CM|AB|289.59|Spleen disease NEC
C0154309|ICD9CM|PT|290.11|Presenile dementia with delirium
C0154309|ICD9CM|AB|290.11|Presenile delirium
C0154310|ICD9CM|PT|290.12|Presenile dementia with delusional features
C0154310|ICD9CM|AB|290.12|Presenile delusion
C0154315|ICD9CM|PT|290.3|Senile dementia with delirium
C0154315|ICD9CM|AB|290.3|Senile delirium
C0154319|ICD9CM|PT|290.8|Other specified senile psychotic conditions
C0154319|ICD9CM|AB|290.8|Senile psychosis NEC
C0154325|ICD9CM|HT|292.8|Other specified drug-induced mental disorders
C0154325|ICD9CM|PT|292.89|Other specified drug-induced mental disorders
C0154325|ICD9CM|AB|292.89|Drug mental disorder NEC
C0154326|ICD9CM|AB|292.81|Drug-induced delirium
C0154326|ICD9CM|PT|292.81|Drug-induced delirium
C0154330|ICD9CM|PT|292.9|Unspecified drug-induced mental disorder
C0154330|ICD9CM|HT|292|Drug-induced mental disorders
C0154330|ICD9CM|AB|292.9|Drug mental disorder NOS
C0154333|ICD9CM|AB|293.1|Subacute delirium
C0154333|ICD9CM|PT|293.1|Subacute delirium
C0154334|ICD9CM|PT|293.89|Other specified transient mental disorders due to conditions classified elsewhere, other
C0154334|ICD9CM|AB|293.89|Transient mental dis NEC
C0154336|ICD9CM|HT|294|Persistent mental disorders due to conditions classified elsewhere
C0154338|ICD9CM|PT|294.8|Other persistent mental disorders due to conditions classified elsewhere
C0154338|ICD9CM|AB|294.8|Mental disor NEC oth dis
C0154339|ICD9CM|PT|295.01|Simple type schizophrenia, subchronic
C0154339|ICD9CM|AB|295.01|Simpl schizophren-subchr
C0154340|ICD9CM|PT|295.02|Simple type schizophrenia, chronic
C0154340|ICD9CM|AB|295.02|Simple schizophren-chr
C0154341|ICD9CM|PT|295.03|Simple type schizophrenia, subchronic with acute exacerbation
C0154341|ICD9CM|AB|295.03|Simp schiz-subchr/exacer
C0154342|ICD9CM|PT|295.04|Simple type schizophrenia, chronic with acute exacerbation
C0154342|ICD9CM|AB|295.04|Simpl schizo-chr/exacerb
C0154343|ICD9CM|PT|295.05|Simple type schizophrenia, in remission
C0154343|ICD9CM|AB|295.05|Simpl schizophren-remiss
C0154344|ICD9CM|AB|295.11|Hebephrenia-subchronic
C0154344|ICD9CM|PT|295.11|Disorganized type schizophrenia, subchronic
C0154345|ICD9CM|AB|295.12|Hebephrenia-chronic
C0154345|ICD9CM|PT|295.12|Disorganized type schizophrenia, chronic
C0154346|ICD9CM|PT|295.13|Disorganized type schizophrenia, subchronic with acute exacerbation
C0154346|ICD9CM|AB|295.13|Hebephren-subchr/exacerb
C0154347|ICD9CM|PT|295.14|Disorganized type schizophrenia, chronic with acute exacerbation
C0154347|ICD9CM|AB|295.14|Hebephrenia-chr/exacerb
C0154349|ICD9CM|AB|295.21|Catatonia-subchronic
C0154349|ICD9CM|PT|295.21|Catatonic type schizophrenia, subchronic
C0154350|ICD9CM|AB|295.22|Catatonia-chronic
C0154350|ICD9CM|PT|295.22|Catatonic type schizophrenia, chronic
C0154351|ICD9CM|PT|295.23|Catatonic type schizophrenia, subchronic with acute exacerbation
C0154351|ICD9CM|AB|295.23|Catatonia-subchr/exacerb
C0154352|ICD9CM|PT|295.24|Catatonic type schizophrenia, chronic with acute exacerbation
C0154352|ICD9CM|AB|295.24|Catatonia-chr/exacerb
C0154354|ICD9CM|PT|295.31|Paranoid type schizophrenia, subchronic
C0154354|ICD9CM|AB|295.31|Paranoid schizo-subchr
C0154356|ICD9CM|PT|295.33|Paranoid type schizophrenia, subchronic with acute exacerbation
C0154356|ICD9CM|AB|295.33|Paran schizo-subchr/exac
C0154357|ICD9CM|PT|295.34|Paranoid type schizophrenia, chronic with acute exacerbation
C0154357|ICD9CM|AB|295.34|Paran schizo-chr/exacerb
C0154358|ICD9CM|PT|295.35|Paranoid type schizophrenia, in remission
C0154358|ICD9CM|AB|295.35|Paranoid schizo-remiss
C0154360|ICD9CM|PT|295.41|Schizophreniform disorder, subchronic
C0154360|ICD9CM|AB|295.41|Schizophrenic dis-subchr
C0154361|ICD9CM|PT|295.42|Schizophreniform disorder, chronic
C0154361|ICD9CM|AB|295.42|Schizophren dis-chronic
C0154362|ICD9CM|AB|295.43|Schizo dis-subchr/exacer
C0154362|ICD9CM|PT|295.43|Schizophreniform disorder, subchronic with acute exacerbation
C0154363|ICD9CM|AB|295.44|Schizophr dis-chr/exacer
C0154363|ICD9CM|PT|295.44|Schizophreniform disorder, chronic with acute exacerbation
C0154364|ICD9CM|AB|295.45|Schizophrenic dis-remiss
C0154364|ICD9CM|PT|295.45|Schizophreniform disorder, in remission
C0154369|ICD9CM|PT|295.55|Latent schizophrenia, in remission
C0154369|ICD9CM|AB|295.55|Lat schizophren-remiss
C0154372|ICD9CM|PT|295.63|Schizophrenic disorders, residual type, subchronic with acute exacerbation
C0154372|ICD9CM|AB|295.63|Schizo resid subchr/exac
C0154373|ICD9CM|PT|295.64|Schizophrenic disorders, residual type, chronic with acute exacerbation
C0154373|ICD9CM|AB|295.64|Schizoph resid-chro/exac
C0154374|ICD9CM|PT|295.65|Schizophrenic disorders, residual type, in remission
C0154374|ICD9CM|AB|295.65|Schizoph dis resid-remis
C0154375|ICD9CM|PT|295.71|Schizoaffective disorder, subchronic
C0154375|ICD9CM|AB|295.71|Schizoaffectv dis-subchr
C0154376|ICD9CM|PT|295.72|Schizoaffective disorder, chronic
C0154376|ICD9CM|AB|295.72|Schizoaffective dis-chr
C0154377|ICD9CM|AB|295.73|Schizoaff dis-subch/exac
C0154377|ICD9CM|PT|295.73|Schizoaffective disorder, subchronic with acute exacerbation
C0154378|ICD9CM|AB|295.74|Schizoafftv dis-chr/exac
C0154378|ICD9CM|PT|295.74|Schizoaffective disorder, chronic with acute exacerbation
C0154380|ICD9CM|PT|295.81|Other specified types of schizophrenia, subchronic
C0154380|ICD9CM|AB|295.81|Schizophrenia NEC-subchr
C0154381|ICD9CM|PT|295.82|Other specified types of schizophrenia, chronic
C0154381|ICD9CM|AB|295.82|Schizophrenia NEC-chr
C0154382|ICD9CM|PT|295.83|Other specified types of schizophrenia, subchronic with acute exacerbation
C0154382|ICD9CM|AB|295.83|Schizo NEC-subchr/exacer
C0154383|ICD9CM|PT|295.84|Other specified types of schizophrenia, chronic with acute exacerbation
C0154383|ICD9CM|AB|295.84|Schizo NEC-chr/exacerb
C0154384|ICD9CM|PT|295.85|Other specified types of schizophrenia, in remission
C0154384|ICD9CM|AB|295.85|Schizophrenia NEC-remiss
C0154387|ICD9CM|PT|295.93|Unspecified schizophrenia, subchronic with acute exacerbation
C0154387|ICD9CM|AB|295.93|Schizo NOS-subchr/exacer
C0154388|ICD9CM|PT|295.94|Unspecified schizophrenia, chronic with acute exacerbation
C0154388|ICD9CM|AB|295.94|Schizo NOS-chr/exacerb
C0154392|ICD9CM|PT|296.03|Bipolar I disorder, single manic episode, severe, without mention of psychotic behavior
C0154392|ICD9CM|AB|296.03|Bipol I sing-sev w/o psy
C0154393|ICD9CM|PT|296.04|Bipolar I disorder, single manic episode, severe, specified as with psychotic behavior
C0154393|ICD9CM|AB|296.04|Bipo I sin man-sev w psy
C0154397|ICD9CM|PT|296.11|Manic affective disorder, recurrent episode, mild
C0154397|ICD9CM|AB|296.11|Recur manic dis-mild
C0154398|ICD9CM|PT|296.12|Manic affective disorder, recurrent episode, moderate
C0154398|ICD9CM|AB|296.12|Recur manic dis-mod
C0154399|ICD9CM|PT|296.13|Manic affective disorder, recurrent episode, severe, without mention of psychotic behavior
C0154399|ICD9CM|AB|296.13|Recur manic dis-severe
C0154400|ICD9CM|PT|296.14|Manic affective disorder, recurrent episode, severe, specified as with psychotic behavior
C0154400|ICD9CM|AB|296.14|Recur manic-sev w psycho
C0154403|ICD9CM|PT|296.21|Major depressive affective disorder, single episode, mild
C0154403|ICD9CM|AB|296.21|Depress psychosis-mild
C0154404|ICD9CM|PT|296.22|Major depressive affective disorder, single episode, moderate
C0154404|ICD9CM|AB|296.22|Depressive psychosis-mod
C0154405|ICD9CM|PT|296.23|Major depressive affective disorder, single episode, severe, without mention of psychotic behavior
C0154405|ICD9CM|AB|296.23|Depress psychosis-severe
C0154406|ICD9CM|PT|296.24|Major depressive affective disorder, single episode, severe, specified as with psychotic behavior
C0154406|ICD9CM|AB|296.24|Depr psychos-sev w psych
C0154408|ICD9CM|PT|296.26|Major depressive affective disorder, single episode, in full remission
C0154408|ICD9CM|AB|296.26|Depr psychos-full remiss
C0154409|ICD9CM|HT|296.3|Major depressive disorder, recurrent episode
C0154409|ICD9CM|PT|296.30|Major depressive affective disorder, recurrent episode, unspecified
C0154409|ICD9CM|AB|296.30|Recurr depr psychos-unsp
C0154411|ICD9CM|PT|296.32|Major depressive affective disorder, recurrent episode, moderate
C0154411|ICD9CM|AB|296.32|Recurr depr psychos-mod
C0154412|ICD9CM|PT|296.33|Major depressive affective disorder, recurrent episode, severe, without mention of psychotic behavior
C0154412|ICD9CM|AB|296.33|Recur depr psych-severe
C0154413|ICD9CM|PT|296.34|Major depressive affective disorder, recurrent episode, severe, specified as with psychotic behavior
C0154413|ICD9CM|AB|296.34|Rec depr psych-psychotic
C0154417|ICD9CM|PT|296.41|Bipolar I disorder, most recent episode (or current) manic, mild
C0154417|ICD9CM|AB|296.41|Bipol I curnt manic-mild
C0154418|ICD9CM|PT|296.42|Bipolar I disorder, most recent episode (or current) manic, moderate
C0154418|ICD9CM|AB|296.42|Bipol I currnt manic-mod
C0154419|ICD9CM|PT|296.43|Bipolar I disorder, most recent episode (or current) manic, severe, without mention of psychotic behavior
C0154419|ICD9CM|AB|296.43|Bipol I manc-sev w/o psy
C0154420|ICD9CM|PT|296.44|Bipolar I disorder, most recent episode (or current) manic, severe, specified as with psychotic behavior
C0154420|ICD9CM|AB|296.44|Bipol I manic-sev w psy
C0154421|ICD9CM|PT|296.45|Bipolar I disorder, most recent episode (or current) manic, in partial or unspecified remission
C0154421|ICD9CM|AB|296.45|Bipol I cur man part rem
C0154422|ICD9CM|PT|296.46|Bipolar I disorder, most recent episode (or current) manic, in full remission
C0154422|ICD9CM|AB|296.46|Bipol I cur man full rem
C0154424|ICD9CM|PT|296.51|Bipolar I disorder, most recent episode (or current) depressed, mild
C0154424|ICD9CM|AB|296.51|Bipol I cur depress-mild
C0154425|ICD9CM|PT|296.52|Bipolar I disorder, most recent episode (or current) depressed, moderate
C0154425|ICD9CM|AB|296.52|Bipol I cur depress-mod
C0154426|ICD9CM|PT|296.53|Bipolar I disorder, most recent episode (or current) depressed, severe, without mention of psychotic behavior
C0154426|ICD9CM|AB|296.53|Bipol I curr dep w/o psy
C0154427|ICD9CM|PT|296.54|Bipolar I disorder, most recent episode (or current) depressed, severe, specified as with psychotic behavior
C0154427|ICD9CM|AB|296.54|Bipol I currnt dep w psy
C0154428|ICD9CM|PT|296.55|Bipolar I disorder, most recent episode (or current) depressed, in partial or unspecified remission
C0154428|ICD9CM|AB|296.55|Bipol I cur dep rem NOS
C0154429|ICD9CM|PT|296.56|Bipolar I disorder, most recent episode (or current) depressed, in full remission
C0154429|ICD9CM|AB|296.56|Bipol I currnt dep remis
C0154432|ICD9CM|PT|296.63|Bipolar I disorder, most recent episode (or current) mixed, severe, without mention of psychotic behavior
C0154432|ICD9CM|AB|296.63|Bipol I cur mix w/o psy
C0154433|ICD9CM|PT|296.64|Bipolar I disorder, most recent episode (or current) mixed, severe, specified as with psychotic behavior
C0154433|ICD9CM|AB|296.64|Bipol I cur mixed w psy
C0154434|ICD9CM|PT|296.65|Bipolar I disorder, most recent episode (or current) mixed, in partial or unspecified remission
C0154434|ICD9CM|AB|296.65|Bipol I cur mix-part rem
C0154436|ICD9CM|AB|296.81|Atypical manic disorder
C0154436|ICD9CM|PT|296.81|Atypical manic disorder
C0154437|ICD9CM|PT|296.82|Atypical depressive disorder
C0154437|ICD9CM|AB|296.82|Atypical depressive dis
C0154440|ICD9CM|AB|297.0|Paranoid state, simple
C0154440|ICD9CM|PT|297.0|Paranoid state, simple
C0154441|ICD9CM|PT|297.8|Other specified paranoid states
C0154441|ICD9CM|AB|297.8|Paranoid states NEC
C0154442|ICD9CM|HT|298|Other nonorganic psychoses
C0154446|ICD9CM|PT|299.00|Autistic disorder, current or active state
C0154446|ICD9CM|AB|299.00|Autistic disord-current
C0154448|ICD9CM|PT|299.10|Childhood disintegrative disorder, current or active state
C0154448|ICD9CM|AB|299.10|Childhd disintegr-active
C0154449|ICD9CM|AB|299.11|Childhd disintegr-resid
C0154449|ICD9CM|PT|299.11|Childhood disintegrative disorder, residual state
C0154451|ICD9CM|PT|299.80|Other specified pervasive developmental disorders, current or active state
C0154451|ICD9CM|AB|299.80|Pervasv dev dis-cur NEC
C0154452|ICD9CM|PT|299.81|Other specified pervasive developmental disorders, residual state
C0154452|ICD9CM|AB|299.81|Pervasv dev dis-res NEC
C0154453|ICD9CM|PT|299.90|Unspecified pervasive developmental disorder, current or active state
C0154453|ICD9CM|AB|299.90|Pervasv dev dis-cur NOS
C0154454|ICD9CM|PT|299.91|Unspecified pervasive developmental disorder, residual state
C0154454|ICD9CM|AB|299.91|Pervasv dev dis-res NOS
C0154455|ICD9CM|PT|300.09|Other anxiety states
C0154455|ICD9CM|AB|300.09|Anxiety state NEC
C0154456|ICD9CM|PT|300.19|Other and unspecified factitious illness
C0154456|ICD9CM|AB|300.19|Factitious ill NEC/NOS
C0154459|ICD9CM|PT|301.11|Chronic hypomanic personality disorder
C0154459|ICD9CM|AB|301.11|Chronic hypomanic person
C0154462|ICD9CM|PT|302.51|Trans-sexualism with asexual history
C0154462|ICD9CM|AB|302.51|Trans-sexualism, asexual
C0154463|ICD9CM|PT|302.52|Trans-sexualism with homosexual history
C0154463|ICD9CM|AB|302.52|Trans-sexual, homosexual
C0154464|ICD9CM|PT|302.53|Trans-sexualism with heterosexual history
C0154464|ICD9CM|AB|302.53|Trans-sex, heterosexual
C0154466|ICD9CM|PT|302.76|Dyspareunia, psychogenic
C0154466|ICD9CM|AB|302.76|Dyspareunia,psychogenic
C0154467|ICD9CM|PT|302.85|Gender identity disorder in adolescents or adults
C0154467|ICD9CM|AB|302.85|Gend iden dis,adol/adult
C0154473|ICD9CM|PT|303.03|Acute alcoholic intoxication in alcoholism, in remission
C0154473|ICD9CM|AB|303.03|Ac alcohol intox-remiss
C0154474|ICD9CM|PT|303.90|Other and unspecified alcohol dependence, unspecified
C0154474|ICD9CM|HT|303.9|Other and unspecified alcohol dependence
C0154474|ICD9CM|AB|303.90|Alcoh dep NEC/NOS-unspec
C0154475|ICD9CM|PT|303.91|Other and unspecified alcohol dependence, continuous
C0154475|ICD9CM|AB|303.91|Alcoh dep NEC/NOS-contin
C0154476|ICD9CM|PT|303.92|Other and unspecified alcohol dependence, episodic
C0154476|ICD9CM|AB|303.92|Alcoh dep NEC/NOS-episod
C0154477|ICD9CM|PT|303.93|Other and unspecified alcohol dependence, in remission
C0154477|ICD9CM|AB|303.93|Alcoh dep NEC/NOS-remiss
C0154478|ICD9CM|PT|304.01|Opioid type dependence, continuous
C0154478|ICD9CM|AB|304.01|Opioid dependence-contin
C0154479|ICD9CM|PT|304.02|Opioid type dependence, episodic
C0154479|ICD9CM|AB|304.02|Opioid dependence-episod
C0154480|ICD9CM|PT|304.03|Opioid type dependence, in remission
C0154480|ICD9CM|AB|304.03|Opioid dependence-remiss
C0154482|ICD9CM|PT|304.11|Sedative, hypnotic or anxiolytic dependence, continuous
C0154482|ICD9CM|AB|304.11|Sed,hyp,anxiolyt dep-con
C0154483|ICD9CM|PT|304.12|Sedative, hypnotic or anxiolytic dependence, episodic
C0154483|ICD9CM|AB|304.12|Sed,hyp,anxiolyt dep-epi
C0154487|ICD9CM|PT|304.23|Cocaine dependence, in remission
C0154487|ICD9CM|AB|304.23|Cocaine depend-remiss
C0154490|ICD9CM|PT|304.33|Cannabis dependence, in remission
C0154490|ICD9CM|AB|304.33|Cannabis depend-remiss
C0154492|ICD9CM|PT|304.41|Amphetamine and other psychostimulant dependence, continuous
C0154492|ICD9CM|AB|304.41|Amphetamin depend-contin
C0154493|ICD9CM|PT|304.42|Amphetamine and other psychostimulant dependence, episodic
C0154493|ICD9CM|AB|304.42|Amphetamin depend-episod
C0154494|ICD9CM|PT|304.43|Amphetamine and other psychostimulant dependence, in remission
C0154494|ICD9CM|AB|304.43|Amphetamin depend-remiss
C0154497|ICD9CM|PT|304.53|Hallucinogen dependence, in remission
C0154497|ICD9CM|AB|304.53|Hallucinogen dep-remiss
C0154500|ICD9CM|PT|304.63|Other specified drug dependence, in remission
C0154500|ICD9CM|AB|304.63|Drug depend NEC-in rem
C0154501|ICD9CM|HT|304.7|Combinations of opioid type drug with any other drug dependence
C0154502|ICD9CM|PT|304.71|Combinations of opioid type drug with any other drug dependence, continuous
C0154502|ICD9CM|AB|304.71|Opioid/other dep-contin
C0154503|ICD9CM|PT|304.72|Combinations of opioid type drug with any other drug dependence, episodic
C0154503|ICD9CM|AB|304.72|Opioid/other dep-episod
C0154504|ICD9CM|PT|304.73|Combinations of opioid type drug with any other drug dependence, in remission
C0154504|ICD9CM|AB|304.73|Opioid/other dep-remiss
C0154505|ICD9CM|HT|304.8|Combinations of drug dependence excluding opioid type drug
C0154506|ICD9CM|PT|304.81|Combinations of drug dependence excluding opioid type drug, continuous
C0154506|ICD9CM|AB|304.81|Comb drug dep NEC-contin
C0154507|ICD9CM|PT|304.82|Combinations of drug dependence excluding opioid type drug, episodic
C0154507|ICD9CM|AB|304.82|Comb drug dep NEC-episod
C0154508|ICD9CM|PT|304.83|Combinations of drug dependence excluding opioid type drug, in remission
C0154508|ICD9CM|AB|304.83|Comb drug dep NEC-remiss
C0154509|ICD9CM|AB|304.91|Drug depend NOS-contin
C0154509|ICD9CM|PT|304.91|Unspecified drug dependence, continuous
C0154510|ICD9CM|AB|304.92|Drug depend NOS-episodic
C0154510|ICD9CM|PT|304.92|Unspecified drug dependence, episodic
C0154511|ICD9CM|PT|304.93|Unspecified drug dependence, in remission
C0154511|ICD9CM|AB|304.93|Drug depend NOS-remiss
C0154515|ICD9CM|AB|305.02|Alcohol abuse-episodic
C0154515|ICD9CM|PT|305.02|Alcohol abuse, episodic
C0154516|ICD9CM|PT|305.03|Alcohol abuse, in remission
C0154516|ICD9CM|AB|305.03|Alcohol abuse-in remiss
C0154520|ICD9CM|AB|305.21|Cannabis abuse-contin
C0154520|ICD9CM|PT|305.21|Cannabis abuse, continuous
C0154521|ICD9CM|AB|305.22|Cannabis abuse-episodic
C0154521|ICD9CM|PT|305.22|Cannabis abuse, episodic
C0154522|ICD9CM|PT|305.23|Cannabis abuse, in remission
C0154522|ICD9CM|AB|305.23|Cannabis abuse-in remiss
C0154523|ICD9CM|AB|305.31|Hallucinog abuse-contin
C0154523|ICD9CM|PT|305.31|Hallucinogen abuse, continuous
C0154524|ICD9CM|AB|305.32|Hallucinog abuse-episod
C0154524|ICD9CM|PT|305.32|Hallucinogen abuse, episodic
C0154525|ICD9CM|PT|305.33|Hallucinogen abuse, in remission
C0154525|ICD9CM|AB|305.33|Hallucinog abuse-remiss
C0154527|ICD9CM|PT|305.41|Sedative, hypnotic or anxiolytic abuse, continuous
C0154527|ICD9CM|AB|305.41|Sed,hyp,anxiolytc ab-con
C0154528|ICD9CM|PT|305.42|Sedative, hypnotic or anxiolytic abuse, episodic
C0154528|ICD9CM|AB|305.42|Sed,hyp,anxiolytc ab-epi
C0154529|ICD9CM|PT|305.43|Sedative, hypnotic or anxiolytic abuse, in remission
C0154529|ICD9CM|AB|305.43|Sed,hyp,anxiolytc ab-rem
C0154530|ICD9CM|AB|305.51|Opioid abuse-continuous
C0154530|ICD9CM|PT|305.51|Opioid abuse, continuous
C0154531|ICD9CM|AB|305.52|Opioid abuse-episodic
C0154531|ICD9CM|PT|305.52|Opioid abuse, episodic
C0154532|ICD9CM|PT|305.53|Opioid abuse, in remission
C0154532|ICD9CM|AB|305.53|Opioid abuse-in remiss
C0154533|ICD9CM|PT|305.61|Cocaine abuse, continuous
C0154533|ICD9CM|AB|305.61|Cocaine abuse-continuous
C0154534|ICD9CM|AB|305.62|Cocaine abuse-episodic
C0154534|ICD9CM|PT|305.62|Cocaine abuse, episodic
C0154535|ICD9CM|PT|305.63|Cocaine abuse, in remission
C0154535|ICD9CM|AB|305.63|Cocaine abuse-in remiss
C0154536|ICD9CM|HT|305.7|Amphetamine or related acting sympathomimetic abuse
C0154537|ICD9CM|PT|305.71|Amphetamine or related acting sympathomimetic abuse, continuous
C0154537|ICD9CM|AB|305.71|Amphetamine abuse-contin
C0154538|ICD9CM|PT|305.72|Amphetamine or related acting sympathomimetic abuse, episodic
C0154538|ICD9CM|AB|305.72|Amphetamine abuse-episod
C0154539|ICD9CM|PT|305.73|Amphetamine or related acting sympathomimetic abuse, in remission
C0154539|ICD9CM|AB|305.73|Amphetamine abuse-remiss
C0154540|ICD9CM|HT|305.8|Antidepressant type abuse
C0154541|ICD9CM|PT|305.81|Antidepressant type abuse, continuous
C0154541|ICD9CM|AB|305.81|Antidepress abuse-contin
C0154542|ICD9CM|PT|305.82|Antidepressant type abuse, episodic
C0154542|ICD9CM|AB|305.82|Antidepress abuse-episod
C0154543|ICD9CM|PT|305.83|Antidepressant type abuse, in remission
C0154543|ICD9CM|AB|305.83|Antidepress abuse-remiss
C0154544|ICD9CM|PT|305.90|Other, mixed, or unspecified drug abuse, unspecified
C0154544|ICD9CM|HT|305.9|Other, mixed, or unspecified drug abuse
C0154544|ICD9CM|AB|305.90|Drug abuse NEC-unspec
C0154545|ICD9CM|PT|305.91|Other, mixed, or unspecified drug abuse, continuous
C0154545|ICD9CM|AB|305.91|Drug abuse NEC-contin
C0154546|ICD9CM|PT|305.92|Other, mixed, or unspecified drug abuse, episodic
C0154546|ICD9CM|AB|305.92|Drug abuse NEC-episodic
C0154547|ICD9CM|PT|305.93|Other, mixed, or unspecified drug abuse, in remission
C0154547|ICD9CM|AB|305.93|Drug abuse NEC-in remiss
C0154548|ICD9CM|HT|306|Physiological malfunction arising from mental factors
C0154549|ICD9CM|PT|306.0|Musculoskeletal malfunction arising from mental factors
C0154549|ICD9CM|AB|306.0|Psychogen musculskel dis
C0154551|ICD9CM|PT|306.3|Skin disorder arising from mental factors
C0154551|ICD9CM|AB|306.3|Psychogenic skin disease
C0154552|ICD9CM|HT|306.5|Genitourinary malfunction arising from mental factors
C0154555|ICD9CM|AB|306.52|Psychogenic dysmenorrhea
C0154555|ICD9CM|PT|306.52|Psychogenic dysmenorrhea
C0154557|ICD9CM|PT|306.59|Other genitourinary malfunction arising from mental factors
C0154557|ICD9CM|AB|306.59|Psychogenic gu dis NEC
C0154558|ICD9CM|PT|306.6|Endocrine disorder arising from mental factors
C0154558|ICD9CM|AB|306.6|Psychogen endocrine dis
C0154559|ICD9CM|PT|306.7|Disorder of organs of special sense arising from mental factors
C0154559|ICD9CM|AB|306.7|Psychogenic sensory dis
C0154564|ICD9CM|HT|307.4|Specific disorders of sleep of nonorganic origin
C0154565|ICD9CM|PT|307.40|Nonorganic sleep disorder, unspecified
C0154565|ICD9CM|AB|307.40|Nonorganic sleep dis NOS
C0154566|ICD9CM|PT|307.41|Transient disorder of initiating or maintaining sleep
C0154566|ICD9CM|AB|307.41|Transient insomnia
C0154568|ICD9CM|PT|307.43|Transient disorder of initiating or maintaining wakefulness
C0154568|ICD9CM|AB|307.43|Transient hypersomnia
C0154569|ICD9CM|PT|307.44|Persistent disorder of initiating or maintaining wakefulness
C0154569|ICD9CM|AB|307.44|Persistent hypersomnia
C0154571|ICD9CM|PT|307.47|Other dysfunctions of sleep stages or arousal from sleep
C0154571|ICD9CM|AB|307.47|Sleep stage dysfunc NEC
C0154572|ICD9CM|PT|307.48|Repetitive intrusions of sleep
C0154572|ICD9CM|AB|307.48|Repetit sleep intrusion
C0154573|ICD9CM|PT|307.49|Other specific disorders of sleep of nonorganic origin
C0154573|ICD9CM|AB|307.49|Nonorganic sleep dis NEC
C0154575|ICD9CM|AB|307.53|Rumination disorder
C0154575|ICD9CM|PT|307.53|Rumination disorder
C0154578|ICD9CM|PT|308.0|Predominant disturbance of emotions
C0154578|ICD9CM|AB|308.0|Stress react, emotional
C0154579|ICD9CM|PT|308.1|Predominant disturbance of consciousness
C0154579|ICD9CM|AB|308.1|Stress reaction, fugue
C0154580|ICD9CM|PT|308.2|Predominant psychomotor disturbance
C0154580|ICD9CM|AB|308.2|Stress react, psychomot
C0154581|ICD9CM|PT|308.4|Mixed disorders as reaction to stress
C0154581|ICD9CM|AB|308.4|Stress react, mixed dis
C0154583|ICD9CM|PT|309.1|Prolonged depressive reaction
C0154583|ICD9CM|AB|309.1|Prolong depressive react
C0154584|ICD9CM|HT|309.2|Adjustment reaction with predominant disturbance of other emotions
C0154585|ICD9CM|PT|309.22|Emancipation disorder of adolescence and early adult life
C0154585|ICD9CM|AB|309.22|Emancipation disorder
C0154586|ICD9CM|PT|309.23|Specific academic or work inhibition
C0154586|ICD9CM|AB|309.23|Academic/work inhibition
C0154587|ICD9CM|PT|309.24|Adjustment disorder with anxiety
C0154587|ICD9CM|AB|309.24|Adjustment dis w anxiety
C0154588|ICD9CM|PT|309.28|Adjustment disorder with mixed anxiety and depressed mood
C0154588|ICD9CM|AB|309.28|Adjust dis w anxiety/dep
C0154589|ICD9CM|PT|309.29|Other adjustment reactions with predominant disturbance of other emotions
C0154589|ICD9CM|AB|309.29|Adj react-emotion NEC
C0154592|ICD9CM|HT|309.8|Other specified adjustment reactions
C0154592|ICD9CM|PT|309.89|Other specified adjustment reactions
C0154592|ICD9CM|AB|309.89|Adjustment reaction NEC
C0154594|ICD9CM|PT|309.82|Adjustment reaction with physical symptoms
C0154594|ICD9CM|AB|309.82|Adjust react-phys sympt
C0154595|ICD9CM|PT|309.83|Adjustment reaction with withdrawal
C0154595|ICD9CM|AB|309.83|Adjust react-withdrawal
C0154598|ICD9CM|HT|310.8|Other specified nonpsychotic mental disorders following organic brain damage
C0154598|ICD9CM|PT|310.89|Other specified nonpsychotic mental disorders following organic brain damage
C0154598|ICD9CM|AB|310.89|Nonpsych mntl disord NEC
C0154600|ICD9CM|PT|312.01|Undersocialized conduct disorder, aggressive type, mild
C0154600|ICD9CM|AB|312.01|Unsocial aggression-mild
C0154601|ICD9CM|PT|312.02|Undersocialized conduct disorder, aggressive type, moderate
C0154601|ICD9CM|AB|312.02|Unsocial aggression-mod
C0154602|ICD9CM|PT|312.03|Undersocialized conduct disorder, aggressive type, severe
C0154602|ICD9CM|AB|312.03|Unsocial aggress-severe
C0154603|ICD9CM|HT|312.1|Undersocialized conduct disorder, unaggressive type
C0154604|ICD9CM|PT|312.11|Undersocialized conduct disorder, unaggressive type, mild
C0154604|ICD9CM|AB|312.11|Unsocial unaggress-mild
C0154605|ICD9CM|PT|312.12|Undersocialized conduct disorder, unaggressive type, moderate
C0154605|ICD9CM|AB|312.12|Unsocial unaggress-mod
C0154606|ICD9CM|PT|312.13|Undersocialized conduct disorder, unaggressive type, severe
C0154606|ICD9CM|AB|312.13|Unsocial unaggr-severe
C0154610|ICD9CM|PT|312.35|Isolated explosive disorder
C0154610|ICD9CM|AB|312.35|Isolated explosive dis
C0154613|ICD9CM|HT|313|Disturbance of emotions specific to childhood and adolescence
C0154614|ICD9CM|PT|313.1|Misery and unhappiness disorder specific to childhood and adolescence
C0154614|ICD9CM|AB|313.1|Misery & unhappiness dis
C0154615|ICD9CM|HT|313.2|Sensitivity, shyness, and social withdrawal disorder specific to childhood and adolescence
C0154616|ICD9CM|PT|313.21|Shyness disorder of childhood
C0154616|ICD9CM|AB|313.21|Shyness disorder-child
C0154618|ICD9CM|PT|313.3|Relationship problems specific to childhood and adolescence
C0154618|ICD9CM|AB|313.3|Relationship problems
C0154619|ICD9CM|HT|313.8|Other or mixed emotional disturbances of childhood or adolescence
C0154621|ICD9CM|PT|313.83|Academic underachievement disorder of childhood or adolescence
C0154621|ICD9CM|AB|313.83|Academic underachievment
C0154622|ICD9CM|PT|313.89|Other emotional disturbances of childhood or adolescence
C0154622|ICD9CM|AB|313.89|Emotional dis child NEC
C0154623|ICD9CM|PT|313.9|Unspecified emotional disturbance of childhood or adolescence
C0154623|ICD9CM|AB|313.9|Emotional dis child NOS
C0154627|ICD9CM|PT|314.1|Hyperkinesis with developmental delay
C0154627|ICD9CM|AB|314.1|Hyperkinet w devel delay
C0154628|ICD9CM|PT|314.2|Hyperkinetic conduct disorder
C0154628|ICD9CM|AB|314.2|Hyperkinetic conduct dis
C0154629|ICD9CM|PT|314.8|Other specified manifestations of hyperkinetic syndrome
C0154629|ICD9CM|AB|314.8|Other hyperkinetic synd
C0154631|ICD9CM|PT|315.09|Other specific developmental reading disorder
C0154631|ICD9CM|AB|315.09|Reading disorder NEC
C0154632|ICD9CM|HT|315.3|Developmental speech or language disorder
C0154633|ICD9CM|PT|315.39|Other developmental speech or language disorder
C0154633|ICD9CM|AB|315.39|Speech/language dis NEC
C0154634|ICD9CM|PT|315.5|Mixed development disorder
C0154634|ICD9CM|AB|315.5|Mixed development dis
C0154635|ICD9CM|PT|315.8|Other specified delays in development
C0154635|ICD9CM|AB|315.8|Development delays NEC
C0154637|ICD9CM|PT|316|Psychic factors associated with diseases classified elsewhere
C0154637|ICD9CM|AB|316|Psychic factor w oth dis
C0154639|ICD9CM|AB|320.2|Streptococcal meningitis
C0154639|ICD9CM|PT|320.2|Streptococcal meningitis
C0154640|ICD9CM|PT|320.3|Staphylococcal meningitis
C0154640|ICD9CM|AB|320.3|Staphylococc meningitis
C0154641|ICD9CM|PT|320.7|Meningitis in other bacterial diseases classified elsewhere
C0154641|ICD9CM|AB|320.7|Mening in oth bact dis
C0154642|ICD9CM|HT|320.8|Meningitis due to other specified bacteria
C0154642|ICD9CM|PT|320.89|Meningitis due to other specified bacteria
C0154642|ICD9CM|AB|320.89|Meningitis oth spcf bact
C0154644|ICD9CM|HT|321|Meningitis due to other organisms
C0154645|ICD9CM|PT|321.1|Meningitis in other fungal diseases
C0154645|ICD9CM|AB|321.1|Mening in oth fungal dis
C0154648|ICD9CM|PT|321.4|Meningitis in sarcoidosis
C0154648|ICD9CM|AB|321.4|Meningit d/t sarcoidosis
C0154649|ICD9CM|PT|321.8|Meningitis due to other nonbacterial organisms classified elsewhere
C0154649|ICD9CM|AB|321.8|Mening in oth nonbac dis
C0154651|ICD9CM|AB|322.0|Nonpyogenic meningitis
C0154651|ICD9CM|PT|322.0|Nonpyogenic meningitis
C0154652|ICD9CM|AB|322.1|Eosinophilic meningitis
C0154652|ICD9CM|PT|322.1|Eosinophilic meningitis
C0154653|ICD9CM|AB|322.2|Chronic meningitis
C0154653|ICD9CM|PT|322.2|Chronic meningitis
C0154660|ICD9CM|HT|324|Intracranial and intraspinal abscess
C0154660|ICD9CM|PT|324.9|Intracranial and intraspinal abscess of unspecified site
C0154660|ICD9CM|AB|324.9|Cns abscess NOS
C0154661|ICD9CM|AB|324.1|Intraspinal abscess
C0154661|ICD9CM|PT|324.1|Intraspinal abscess
C0154662|ICD9CM|PT|325|Phlebitis and thrombophlebitis of intracranial venous sinuses
C0154662|ICD9CM|AB|325|Phlebitis intrcran sinus
C0154663|ICD9CM|PT|326|Late effects of intracranial abscess or pyogenic infection
C0154663|ICD9CM|AB|326|Late eff cns abscess
C0154664|ICD9CM|HT|330|Cerebral degenerations usually manifest in childhood
C0154666|ICD9CM|PT|330.3|Cerebral degeneration of childhood in other diseases classified elsewhere
C0154666|ICD9CM|AB|330.3|Cerb deg chld in oth dis
C0154667|ICD9CM|PT|330.9|Unspecified cerebral degeneration in childhood
C0154667|ICD9CM|AB|330.9|Cereb degen in child NOS
C0154668|ICD9CM|HT|331.8|Other cerebral degeneration
C0154668|ICD9CM|PT|331.89|Other cerebral degeneration
C0154668|ICD9CM|HT|331|Other cerebral degenerations
C0154668|ICD9CM|AB|331.89|Cereb degeneration NEC
C0154669|ICD9CM|PT|331.2|Senile degeneration of brain
C0154669|ICD9CM|AB|331.2|Senile degenerat brain
C0154671|ICD9CM|PT|331.9|Cerebral degeneration, unspecified
C0154671|ICD9CM|AB|331.9|Cereb degeneration NOS
C0154675|ICD9CM|HT|333.8|Fragments of torsion dystonia
C0154676|ICD9CM|AB|333.84|Organic writers' cramp
C0154676|ICD9CM|PT|333.84|Organic writers' cramp
C0154677|ICD9CM|PT|333.89|Other fragments of torsion dystonia
C0154677|ICD9CM|AB|333.89|Fragm torsion dyston NEC
C0154678|ICD9CM|PT|333.99|Other extrapyramidal diseases and abnormal movement disorders
C0154678|ICD9CM|HT|333|Other extrapyramidal disease and abnormal movement disorders
C0154678|ICD9CM|HT|333.9|Other and unspecified extrapyramidal diseases and abnormal movement disorders
C0154678|ICD9CM|AB|333.99|Extrapyramidal dis NEC
C0154681|ICD9CM|HT|335|Anterior horn cell disease
C0154681|ICD9CM|PT|335.9|Anterior horn cell disease, unspecified
C0154681|ICD9CM|AB|335.9|Ant horn cell dis NOS
C0154682|ICD9CM|PT|335.24|Primary lateral sclerosis
C0154682|ICD9CM|AB|335.24|Prim lateral sclerosis
C0154683|ICD9CM|PT|335.29|Other motor neuron disease
C0154683|ICD9CM|AB|335.29|Motor neuron disease NEC
C0154684|ICD9CM|PT|335.8|Other anterior horn cell diseases
C0154684|ICD9CM|AB|335.8|Ant horn cell dis NEC
C0154685|ICD9CM|AB|336.1|Vascular myelopathies
C0154685|ICD9CM|PT|336.1|Vascular myelopathies
C0154686|ICD9CM|PT|336.2|Subacute combined degeneration of spinal cord in diseases classified elsewhere
C0154686|ICD9CM|AB|336.2|Comb deg cord in oth dis
C0154687|ICD9CM|PT|336.3|Myelopathy in other diseases classified elsewhere
C0154687|ICD9CM|AB|336.3|Myelopathy in oth dis
C0154688|ICD9CM|HT|336|Other diseases of spinal cord
C0154690|ICD9CM|HT|337.0|Idiopathic peripheral autonomic neuropathy
C0154691|ICD9CM|PT|337.1|Peripheral autonomic neuropathy in disorders classified elsewhere
C0154691|ICD9CM|AB|337.1|Aut neuropthy in oth dis
C0154692|ICD9CM|HT|341|Other demyelinating diseases of central nervous system
C0154692|ICD9CM|PT|341.8|Other demyelinating diseases of central nervous system
C0154692|ICD9CM|AB|341.8|Cns demyelination NEC
C0154693|ICD9CM|HT|342.0|Flaccid hemiplegia
C0154693|ICD9CM|PT|342.00|Flaccid hemiplegia and hemiparesis affecting unspecified side
C0154693|ICD9CM|AB|342.00|Flccd hmiplga unspf side
C0154694|ICD9CM|HT|342.1|Spastic hemiplegia
C0154694|ICD9CM|PT|342.10|Spastic hemiplegia and hemiparesis affecting unspecified side
C0154694|ICD9CM|AB|342.10|Spstc hmiplga unspf side
C0154695|ICD9CM|AB|343.0|Congenital diplegia
C0154695|ICD9CM|PT|343.0|Congenital diplegia
C0154697|ICD9CM|AB|343.2|Congenital quadriplegia
C0154697|ICD9CM|PT|343.2|Congenital quadriplegia
C0154698|ICD9CM|AB|343.3|Congenital monoplegia
C0154698|ICD9CM|PT|343.3|Congenital monoplegia
C0154700|ICD9CM|HT|344|Other paralytic syndromes
C0154701|ICD9CM|AB|344.2|Diplegia of upper limbs
C0154701|ICD9CM|PT|344.2|Diplegia of upper limbs
C0154702|ICD9CM|HT|344.3|Monoplegia of lower limb
C0154703|ICD9CM|HT|344.4|Monoplegia of upper limb
C0154703|ICD9CM|PT|344.40|Monoplegia of upper limb affecting unspecified side
C0154703|ICD9CM|AB|344.40|Monplga upr lmb unsp sde
C0154706|ICD9CM|HT|344.8|Other specified paralytic syndromes
C0154706|ICD9CM|PT|344.89|Other specified paralytic syndrome
C0154706|ICD9CM|AB|344.89|Oth spcf paralytic synd
C0154707|ICD9CM|PT|345.00|Generalized nonconvulsive epilepsy, without mention of intractable epilepsy
C0154707|ICD9CM|AB|345.00|Gen noncv ep w/o intr ep
C0154709|ICD9CM|PT|345.10|Generalized convulsive epilepsy, without mention of intractable epilepsy
C0154709|ICD9CM|AB|345.10|Gen cnv epil w/o intr ep
C0154710|ICD9CM|PT|345.11|Generalized convulsive epilepsy, with intractable epilepsy
C0154710|ICD9CM|AB|345.11|Gen cnv epil w intr epil
C0154712|ICD9CM|PT|345.51|Localization-related (focal) (partial) epilepsy and epileptic syndromes with simple partial seizures, with intractable epilepsy
C0154712|ICD9CM|AB|345.51|Part epil w intr epil
C0154713|ICD9CM|PT|345.41|Localization-related (focal) (partial) epilepsy and epileptic syndromes with complex partial seizures, with intractable epilepsy
C0154713|ICD9CM|AB|345.41|Psymotr epil w intr epil
C0154714|ICD9CM|PT|345.50|Localization-related (focal) (partial) epilepsy and epileptic syndromes with simple partial seizures, without mention of intractable epilepsy
C0154714|ICD9CM|AB|345.50|Part epil w/o intr epil
C0154715|ICD9CM|PT|345.60|Infantile spasms, without mention of intractable epilepsy
C0154715|ICD9CM|AB|345.60|Inf spasm w/o intr epil
C0154716|ICD9CM|PT|345.61|Infantile spasms, with intractable epilepsy
C0154716|ICD9CM|AB|345.61|Inf spasm w intract epil
C0154717|ICD9CM|PT|345.70|Epilepsia partialis continua, without mention of intractable epilepsy
C0154717|ICD9CM|AB|345.70|Epil par cont w/o int ep
C0154718|ICD9CM|PT|345.71|Epilepsia partialis continua, with intractable epilepsy
C0154718|ICD9CM|AB|345.71|Epil par cont w intr epi
C0154719|ICD9CM|PT|345.80|Other forms of epilepsy and recurrent seizures, without mention of intractable epilepsy
C0154719|ICD9CM|AB|345.80|Epilep NEC w/o intr epil
C0154720|ICD9CM|PT|345.81|Other forms of epilepsy and recurrent seizures, with intractable epilepsy
C0154720|ICD9CM|AB|345.81|Epilepsy NEC w intr epil
C0154721|ICD9CM|PT|345.90|Epilepsy, unspecified, without mention of intractable epilepsy
C0154721|ICD9CM|AB|345.90|Epilep NOS w/o intr epil
C0154722|ICD9CM|PT|345.91|Epilepsy, unspecified, with intractable epilepsy
C0154722|ICD9CM|AB|345.91|Epilepsy NOS w intr epil
C0154723|ICD9CM|HT|346.0|Migraine with aura
C0154724|ICD9CM|AB|348.0|Cerebral cysts
C0154724|ICD9CM|PT|348.0|Cerebral cysts
C0154725|ICD9CM|HT|349|Other and unspecified disorders of the nervous system
C0154727|ICD9CM|PT|349.1|Nervous system complications from surgically implanted device
C0154727|ICD9CM|AB|349.1|Complication cns device
C0154729|ICD9CM|AB|350.2|Atypical face pain
C0154729|ICD9CM|PT|350.2|Atypical face pain
C0154730|ICD9CM|HT|352|Disorders of other cranial nerves
C0154731|ICD9CM|PT|352.1|Glossopharyngeal neuralgia
C0154731|ICD9CM|AB|352.1|Glossopharyng neuralgia
C0154733|ICD9CM|PT|352.6|Multiple cranial nerve palsies
C0154733|ICD9CM|AB|352.6|Mult cranial nerve palsy
C0154735|ICD9CM|PT|353.1|Lumbosacral plexus lesions
C0154735|ICD9CM|AB|353.1|Lumbosacral plex lesion
C0154739|ICD9CM|PT|353.8|Other nerve root and plexus disorders
C0154739|ICD9CM|AB|353.8|Nerv root/plexus dis NEC
C0154741|ICD9CM|HT|354|Mononeuritis of upper limb and mononeuritis multiplex
C0154742|ICD9CM|PT|354.1|Other lesion of median nerve
C0154742|ICD9CM|AB|354.1|Median nerve lesion NEC
C0154744|ICD9CM|PT|354.3|Lesion of radial nerve
C0154744|ICD9CM|AB|354.3|Radial nerve lesion
C0154745|ICD9CM|PT|354.8|Other mononeuritis of upper limb
C0154745|ICD9CM|AB|354.8|Mononeuritis arm NEC
C0154746|ICD9CM|PT|354.9|Mononeuritis of upper limb, unspecified
C0154746|ICD9CM|AB|354.9|Mononeuritis arm NOS
C0154747|ICD9CM|HT|355|Mononeuritis of lower limb
C0154747|ICD9CM|PT|355.8|Mononeuritis of lower limb, unspecified
C0154747|ICD9CM|AB|355.8|Mononeuritis leg NOS
C0154748|ICD9CM|PT|355.0|Lesion of sciatic nerve
C0154748|ICD9CM|AB|355.0|Sciatic nerve lesion
C0154749|ICD9CM|PT|355.2|Other lesion of femoral nerve
C0154749|ICD9CM|AB|355.2|Femoral nerve lesion NEC
C0154752|ICD9CM|AB|355.6|Plantar nerve lesion
C0154752|ICD9CM|PT|355.6|Lesion of plantar nerve
C0154753|ICD9CM|HT|355.7|Other mononeuritis of lower limb
C0154753|ICD9CM|PT|355.79|Other mononeuritis of lower limb
C0154753|ICD9CM|AB|355.79|Oth mononeur lower limb
C0154754|ICD9CM|HT|356|Hereditary and idiopathic peripheral neuropathy
C0154756|ICD9CM|PT|356.4|Idiopathic progressive polyneuropathy
C0154756|ICD9CM|AB|356.4|Idio prog polyneuropathy
C0154757|ICD9CM|PT|356.8|Other specified idiopathic peripheral neuropathy
C0154757|ICD9CM|AB|356.8|Idio periph neurpthy NEC
C0154758|ICD9CM|HT|357|Inflammatory and toxic neuropathy
C0154758|ICD9CM|PT|357.9|Unspecified inflammatory and toxic neuropathy
C0154758|ICD9CM|AB|357.9|Inflam/tox neuropthy NOS
C0154759|ICD9CM|PT|357.1|Polyneuropathy in collagen vascular disease
C0154759|ICD9CM|AB|357.1|Neurpthy in col vasc dis
C0154761|ICD9CM|PT|357.4|Polyneuropathy in other diseases classified elsewhere
C0154761|ICD9CM|AB|357.4|Neuropathy in other dis
C0154762|ICD9CM|PT|357.6|Polyneuropathy due to drugs
C0154762|ICD9CM|AB|357.6|Neuropathy due to drugs
C0154763|ICD9CM|PT|357.7|Polyneuropathy due to other toxic agents
C0154763|ICD9CM|AB|357.7|Neurpthy toxic agent NEC
C0154764|ICD9CM|PT|357.89|Other inflammatory and toxic neuropathy
C0154764|ICD9CM|HT|357.8|Other inflammatory and toxic neuropathies
C0154764|ICD9CM|AB|357.89|Inflam/tox neuropthy NEC
C0154769|ICD9CM|AB|359.4|Toxic myopathy
C0154769|ICD9CM|PT|359.4|Toxic myopathy
C0154770|ICD9CM|PT|359.5|Myopathy in endocrine diseases classified elsewhere
C0154770|ICD9CM|AB|359.5|Myopathy in endocrin dis
C0154771|ICD9CM|PT|359.6|Symptomatic inflammatory myopathy in diseases classified elsewhere
C0154771|ICD9CM|AB|359.6|Infl myopathy in oth dis
C0154773|ICD9CM|AB|360.01|Acute endophthalmitis
C0154773|ICD9CM|PT|360.01|Acute endophthalmitis
C0154774|ICD9CM|AB|360.03|Chronic endophthalmitis
C0154774|ICD9CM|PT|360.03|Chronic endophthalmitis
C0154775|ICD9CM|AB|360.14|Ophthalmia nodosa
C0154775|ICD9CM|PT|360.14|Ophthalmia nodosa
C0154777|ICD9CM|HT|360.4|Degenerated conditions of globe
C0154777|ICD9CM|PT|360.40|Degenerated globe or eye, unspecified
C0154777|ICD9CM|PT|360.20|Degenerative disorder of globe, unspecified
C0154777|ICD9CM|HT|360.2|Degenerative disorders of globe
C0154777|ICD9CM|AB|360.40|Degeneration of eye NOS
C0154777|ICD9CM|AB|360.20|Degenerat globe dis NOS
C0154778|ICD9CM|PT|360.21|Progressive high (degenerative) myopia
C0154778|ICD9CM|AB|360.21|Progressive high myopia
C0154780|ICD9CM|PT|360.29|Other degenerative disorders of globe
C0154780|ICD9CM|AB|360.29|Degenerative globe NEC
C0154782|ICD9CM|PT|360.31|Primary hypotony of eye
C0154782|ICD9CM|AB|360.31|Primary hypotony
C0154783|ICD9CM|PT|360.32|Ocular fistula causing hypotony
C0154783|ICD9CM|AB|360.32|Hypotony due to fistula
C0154784|ICD9CM|PT|360.33|Hypotony associated with other ocular disorders
C0154784|ICD9CM|AB|360.33|Hypotony w eye dis NEC
C0154788|ICD9CM|AB|360.41|Blind hypotensive eye
C0154788|ICD9CM|PT|360.41|Blind hypotensive eye
C0154789|ICD9CM|AB|360.42|Blind hypertensive eye
C0154789|ICD9CM|PT|360.42|Blind hypertensive eye
C0154792|ICD9CM|PT|360.51|Foreign body, magnetic, in anterior chamber of eye
C0154792|ICD9CM|AB|360.51|Old magnet fb, ant chamb
C0154793|ICD9CM|PT|360.52|Foreign body, magnetic, in iris or ciliary body
C0154793|ICD9CM|AB|360.52|Old magnet fb, iris
C0154794|ICD9CM|PT|360.53|Foreign body, magnetic, in lens
C0154794|ICD9CM|AB|360.53|Old magnet fb, lens
C0154795|ICD9CM|PT|360.54|Foreign body, magnetic, in vitreous
C0154795|ICD9CM|AB|360.54|Old magnet fb, vitreous
C0154796|ICD9CM|PT|360.55|Foreign body, magnetic, in posterior wall
C0154796|ICD9CM|AB|360.55|Old magnet fb, post wall
C0154797|ICD9CM|PT|360.59|Intraocular foreign body, magnetic, in other or multiple sites
C0154797|ICD9CM|AB|360.59|Old magnet fb, eye NEC
C0154799|ICD9CM|PT|360.61|Foreign body in anterior chamber
C0154799|ICD9CM|AB|360.61|FB in anterior chamber
C0154800|ICD9CM|PT|360.62|Foreign body in iris or ciliary body
C0154800|ICD9CM|AB|360.62|FB in iris or ciliary
C0154801|ICD9CM|AB|360.63|Foreign body in lens
C0154801|ICD9CM|PT|360.63|Foreign body in lens
C0154802|ICD9CM|AB|360.64|Foreign body in vitreous
C0154802|ICD9CM|PT|360.64|Foreign body in vitreous
C0154803|ICD9CM|PT|360.65|Foreign body in posterior wall of eye
C0154803|ICD9CM|AB|360.65|FB in posterior wall
C0154804|ICD9CM|PT|360.69|Intraocular foreign body in other or multiple sites
C0154804|ICD9CM|AB|360.69|Intraocular FB NEC
C0154805|ICD9CM|HT|360.8|Other disorders of globe
C0154805|ICD9CM|PT|360.89|Other disorders of globe
C0154805|ICD9CM|AB|360.89|Disorder of globe NEC
C0154806|ICD9CM|AB|360.81|Luxation of globe
C0154806|ICD9CM|PT|360.81|Luxation of globe
C0154808|ICD9CM|HT|361.0|Retinal detachment with retinal defect
C0154808|ICD9CM|PT|361.00|Retinal detachment with retinal defect, unspecified
C0154808|ICD9CM|AB|361.00|Detachmnt w defect NOS
C0154809|ICD9CM|PT|361.01|Recent retinal detachment, partial, with single defect
C0154809|ICD9CM|AB|361.01|Part detach-singl defec
C0154810|ICD9CM|PT|361.02|Recent retinal detachment, partial, with multiple defects
C0154810|ICD9CM|AB|361.02|Part detach-mult defect
C0154811|ICD9CM|PT|361.03|Recent retinal detachment, partial, with giant tear
C0154811|ICD9CM|AB|361.03|Part detach-giant tear
C0154812|ICD9CM|PT|361.04|Recent retinal detachment, partial, with retinal dialysis
C0154812|ICD9CM|AB|361.04|Part detach-dialysis
C0154813|ICD9CM|PT|361.05|Recent retinal detachment, total or subtotal
C0154813|ICD9CM|AB|361.05|Recent detachment, total
C0154814|ICD9CM|PT|361.06|Old retinal detachment, partial
C0154814|ICD9CM|AB|361.06|Old detachment, partial
C0154815|ICD9CM|PT|361.07|Old retinal detachment, total or subtotal
C0154815|ICD9CM|AB|361.07|Old detachment, total
C0154816|ICD9CM|HT|361.1|Retinoschisis and retinal cysts
C0154817|ICD9CM|AB|361.11|Flat retinoschisis
C0154817|ICD9CM|PT|361.11|Flat retinoschisis
C0154819|ICD9CM|AB|361.13|Primary retinal cysts
C0154819|ICD9CM|PT|361.13|Primary retinal cysts
C0154820|ICD9CM|AB|361.14|Secondary retinal cysts
C0154820|ICD9CM|PT|361.14|Secondary retinal cysts
C0154821|ICD9CM|PT|361.19|Other retinoschisis and retinal cysts
C0154821|ICD9CM|AB|361.19|Retinoshisis or cyst NEC
C0154822|ICD9CM|PT|361.2|Serous retinal detachment
C0154822|ICD9CM|AB|361.2|Serous retina detachment
C0154823|ICD9CM|AB|361.30|Retinal defect NOS
C0154823|ICD9CM|PT|361.30|Retinal defect, unspecified
C0154825|ICD9CM|PT|361.31|Round hole of retina without detachment
C0154825|ICD9CM|AB|361.31|Round hole of retina
C0154826|ICD9CM|PT|361.32|Horseshoe tear of retina without detachment
C0154826|ICD9CM|AB|361.32|Horseshoe tear of retina
C0154827|ICD9CM|PT|361.33|Multiple defects of retina without detachment
C0154827|ICD9CM|AB|361.33|Mult defects of retina
C0154828|ICD9CM|PT|361.81|Traction detachment of retina
C0154828|ICD9CM|AB|361.81|Retinal traction detach
C0154830|ICD9CM|PT|362.02|Proliferative diabetic retinopathy
C0154830|ICD9CM|AB|362.02|Prolif diab retinopathy
C0154831|ICD9CM|HT|362.1|Other background retinopathy and retinal vascular changes
C0154832|ICD9CM|AB|362.12|Exudative retinopathy
C0154832|ICD9CM|PT|362.12|Exudative retinopathy
C0154834|ICD9CM|PT|362.14|Retinal microaneurysms NOS
C0154834|ICD9CM|AB|362.14|Retina microaneurysm NOS
C0154835|ICD9CM|AB|362.15|Retinal telangiectasia
C0154835|ICD9CM|PT|362.15|Retinal telangiectasia
C0154836|ICD9CM|PT|362.17|Other intraretinal microvascular abnormalities
C0154836|ICD9CM|AB|362.17|Retinal varices
C0154837|ICD9CM|HT|362.2|Other proliferative retinopathy
C0154838|ICD9CM|PT|362.29|Other nondiabetic proliferative retinopathy
C0154838|ICD9CM|AB|362.29|Prolif retinopathy NEC
C0154839|ICD9CM|PT|362.33|Partial retinal arterial occlusion
C0154839|ICD9CM|AB|362.33|Part arterial occlusion
C0154840|ICD9CM|PT|362.34|Transient retinal arterial occlusion
C0154840|ICD9CM|AB|362.34|Transient arterial occlu
C0154841|ICD9CM|PT|362.35|Central retinal vein occlusion
C0154841|ICD9CM|AB|362.35|Cent retinal vein occlus
C0154842|ICD9CM|PT|362.36|Venous tributary (branch) occlusion
C0154842|ICD9CM|AB|362.36|Venous tributary occlus
C0154843|ICD9CM|PT|362.37|Venous engorgement
C0154843|ICD9CM|AB|362.37|Retina venous engorgemnt
C0154844|ICD9CM|HT|362.4|Separation of retinal layers
C0154844|ICD9CM|PT|362.40|Retinal layer separation, unspecified
C0154844|ICD9CM|AB|362.40|Retina layer separat NOS
C0154845|ICD9CM|PT|362.42|Serous detachment of retinal pigment epithelium
C0154845|ICD9CM|AB|362.42|Serous detach pigm epith
C0154846|ICD9CM|PT|362.43|Hemorrhagic detachment of retinal pigment epithelium
C0154846|ICD9CM|AB|362.43|Hem detach pigmnt epith
C0154850|ICD9CM|PT|362.53|Cystoid macular degeneration
C0154850|ICD9CM|AB|362.53|Cystoid macular degen
C0154854|ICD9CM|PT|362.61|Paving stone degeneration
C0154854|ICD9CM|AB|362.61|Paving stone degenerat
C0154855|ICD9CM|PT|362.62|Microcystoid degeneration
C0154855|ICD9CM|AB|362.62|Microcystoid degenerat
C0154856|ICD9CM|AB|362.63|Lattice degeneration
C0154856|ICD9CM|PT|362.63|Lattice degeneration
C0154857|ICD9CM|PT|362.64|Senile reticular degeneration
C0154857|ICD9CM|AB|362.64|Senile reticular degen
C0154858|ICD9CM|AB|362.65|Secondry pigment degen
C0154858|ICD9CM|PT|362.65|Secondary pigmentary degeneration
C0154859|ICD9CM|PT|362.66|Secondary vitreoretinal degenerations
C0154859|ICD9CM|AB|362.66|Sec vitreoretina degen
C0154860|ICD9CM|HT|362.7|Hereditary retinal dystrophies
C0154860|ICD9CM|PT|362.70|Hereditary retinal dystrophy, unspecified
C0154860|ICD9CM|AB|362.70|Hered retin dystrphy NOS
C0154861|ICD9CM|PT|362.71|Retinal dystrophy in systemic or cerebroretinal lipidoses
C0154861|ICD9CM|AB|362.71|Ret dystrph in lipidoses
C0154862|ICD9CM|PT|362.72|Retinal dystrophy in other systemic disorders and syndromes
C0154862|ICD9CM|AB|362.72|Ret dystrph in syst dis
C0154863|ICD9CM|AB|362.73|Vitreoretinal dystrophy
C0154863|ICD9CM|PT|362.73|Vitreoretinal dystrophies
C0154864|ICD9CM|PT|362.75|Other dystrophies primarily involving the sensory retina
C0154864|ICD9CM|AB|362.75|Sensory retina dystrophy
C0154865|ICD9CM|PT|362.76|Dystrophies primarily involving the retinal pigment epithelium
C0154865|ICD9CM|AB|362.76|Vitelliform dystrophy
C0154866|ICD9CM|PT|362.77|Dystrophies primarily involving Bruch's membrane
C0154866|ICD9CM|AB|362.77|Bruch membrane dystrophy
C0154867|ICD9CM|PT|362.82|Retinal exudates and deposits
C0154867|ICD9CM|AB|362.82|Retina exudates/deposits
C0154870|ICD9CM|HT|363.0|Focal chorioretinitis and focal retinochoroiditis
C0154870|ICD9CM|PT|363.00|Focal chorioretinitis, unspecified
C0154870|ICD9CM|AB|363.00|Focal chorioretinit NOS
C0154871|ICD9CM|PT|363.01|Focal choroiditis and chorioretinitis, juxtapapillary
C0154871|ICD9CM|AB|363.01|Juxtapap foc choroiditis
C0154872|ICD9CM|PT|363.03|Focal choroiditis and chorioretinitis of other posterior pole
C0154872|ICD9CM|AB|363.03|Foc choroiditis post NEC
C0154875|ICD9CM|PT|363.06|Focal retinitis and retinochoroiditis, macular or paramacular
C0154875|ICD9CM|AB|363.06|Macular focal retinitis
C0154876|ICD9CM|PT|363.07|Focal retinitis and retinochoroiditis of other posterior pole
C0154876|ICD9CM|AB|363.07|Foc retinitis post NEC
C0154877|ICD9CM|PT|363.08|Focal retinitis and retinochoroiditis, peripheral
C0154877|ICD9CM|AB|363.08|Periph focal retinitis
C0154879|ICD9CM|HT|363.1|Disseminated chorioretinitis and disseminated retinochoroiditis
C0154879|ICD9CM|PT|363.10|Disseminated chorioretinitis, unspecified
C0154879|ICD9CM|AB|363.10|Dissem chorioretinit NOS
C0154880|ICD9CM|PT|363.11|Disseminated choroiditis and chorioretinitis, posterior pole
C0154880|ICD9CM|AB|363.11|Dissem choroiditis, post
C0154881|ICD9CM|PT|363.12|Disseminated choroiditis and chorioretinitis, peripheral
C0154881|ICD9CM|AB|363.12|Periph disem choroiditis
C0154882|ICD9CM|PT|363.13|Disseminated choroiditis and chorioretinitis, generalized
C0154882|ICD9CM|AB|363.13|Gen dissem choroiditis
C0154883|ICD9CM|PT|363.14|Disseminated retinitis and retinochoroiditis, metastatic
C0154883|ICD9CM|AB|363.14|Metastat dissem retinit
C0154884|ICD9CM|PT|363.15|Disseminated retinitis and retinochoroiditis, pigment epitheliopathy
C0154884|ICD9CM|AB|363.15|Pigment epitheliopathy
C0154888|ICD9CM|PT|363.34|Peripheral scars
C0154888|ICD9CM|AB|363.34|Peripheral retinal scars
C0154889|ICD9CM|PT|363.35|Disseminated scars
C0154889|ICD9CM|AB|363.35|Disseminated retina scar
C0154891|ICD9CM|PT|363.41|Senile atrophy of choroid
C0154891|ICD9CM|AB|363.41|Senile atrophy, choroid
C0154892|ICD9CM|PT|363.42|Diffuse secondary atrophy of choroid
C0154892|ICD9CM|AB|363.42|Difus sec atroph choroid
C0154893|ICD9CM|HT|363.5|Hereditary choroidal dystrophies
C0154893|ICD9CM|PT|363.50|Hereditary choroidal dystrophy or atrophy, unspecified
C0154893|ICD9CM|AB|363.50|Hered choroid atroph NOS
C0154895|ICD9CM|PT|363.51|Circumpapillary dystrophy of choroid, partial
C0154895|ICD9CM|AB|363.51|Prt circmpap choroid dys
C0154896|ICD9CM|PT|363.52|Circumpapillary dystrophy of choroid, total
C0154896|ICD9CM|AB|363.52|Tot circmpap choroid dys
C0154898|ICD9CM|PT|363.54|Central choroidal atrophy, total
C0154898|ICD9CM|AB|363.54|Tot cent choroid atrophy
C0154899|ICD9CM|PT|363.56|Other diffuse or generalized dystrophy of choroid, partial
C0154899|ICD9CM|AB|363.56|Prt gen choroid dyst NEC
C0154900|ICD9CM|PT|363.57|Other diffuse or generalized dystrophy of choroid, total
C0154900|ICD9CM|AB|363.57|Tot gen choroid dyst NEC
C0154901|ICD9CM|HT|363.6|Choroidal hemorrhage and rupture
C0154902|ICD9CM|PT|363.62|Expulsive choroidal hemorrhage
C0154902|ICD9CM|AB|363.62|Expulsive choroid hemorr
C0154903|ICD9CM|AB|363.63|Choroidal rupture
C0154903|ICD9CM|PT|363.63|Choroidal rupture
C0154904|ICD9CM|PT|363.71|Serous choroidal detachment
C0154904|ICD9CM|AB|363.71|Serous choroid detachmnt
C0154905|ICD9CM|PT|363.72|Hemorrhagic choroidal detachment
C0154905|ICD9CM|AB|363.72|Hemorr choroid detachmnt
C0154906|ICD9CM|PT|363.8|Other disorders of choroid
C0154906|ICD9CM|AB|363.8|Disorders of choroid NEC
C0154907|ICD9CM|HT|364|Disorders of iris and ciliary body
C0154907|ICD9CM|PT|364.9|Unspecified disorder of iris and ciliary body
C0154907|ICD9CM|AB|364.9|Iris/ciliary dis NOS
C0154908|ICD9CM|HT|364.0|Acute and subacute iridocyclitis
C0154908|ICD9CM|AB|364.00|Acute iridocyclitis NOS
C0154908|ICD9CM|PT|364.00|Acute and subacute iridocyclitis, unspecified
C0154909|ICD9CM|AB|364.01|Primary iridocyclitis
C0154909|ICD9CM|PT|364.01|Primary iridocyclitis
C0154910|ICD9CM|AB|364.02|Recurrent iridocyclitis
C0154910|ICD9CM|PT|364.02|Recurrent iridocyclitis
C0154911|ICD9CM|PT|364.03|Secondary iridocyclitis, infectious
C0154911|ICD9CM|AB|364.03|Secondry iritis, infect
C0154915|ICD9CM|HT|364.4|Vascular disorders of iris and ciliary body
C0154916|ICD9CM|AB|364.42|Rubeosis iridis
C0154916|ICD9CM|PT|364.42|Rubeosis iridis
C0154917|ICD9CM|HT|364.5|Degenerations of iris and ciliary body
C0154919|ICD9CM|AB|364.52|Iridoschisis
C0154919|ICD9CM|PT|364.52|Iridoschisis
C0154921|ICD9CM|PT|364.54|Degeneration of pupillary margin
C0154921|ICD9CM|AB|364.54|Pupillary margin degen
C0154922|ICD9CM|PT|364.55|Miotic cysts of pupillary margin
C0154922|ICD9CM|AB|364.55|Miotic cyst pupil margin
C0154923|ICD9CM|PT|364.56|Degenerative changes of chamber angle
C0154923|ICD9CM|AB|364.56|Degen chamber angle
C0154924|ICD9CM|PT|364.57|Degenerative changes of ciliary body
C0154924|ICD9CM|AB|364.57|Degen ciliary body
C0154925|ICD9CM|PT|364.59|Other iris atrophy
C0154925|ICD9CM|AB|364.59|Iris atrophy NEC
C0154926|ICD9CM|HT|364.6|Cysts of iris, ciliary body, and anterior chamber
C0154927|ICD9CM|PT|364.60|Idiopathic cysts of iris, ciliary body, and anterior chamber
C0154927|ICD9CM|AB|364.60|Idiopathic cysts
C0154929|ICD9CM|PT|364.62|Exudative cysts of iris or anterior chamber
C0154929|ICD9CM|AB|364.62|Exud cyst iris/ant chamb
C0154930|ICD9CM|PT|364.63|Primary cyst of pars plana
C0154930|ICD9CM|AB|364.63|Primary cyst pars plana
C0154931|ICD9CM|PT|364.64|Exudative cyst of pars plana
C0154931|ICD9CM|AB|364.64|Exudat cyst pars plana
C0154932|ICD9CM|HT|364.7|Adhesions and disruptions of iris and ciliary body
C0154933|ICD9CM|AB|364.70|Adhesions of iris NOS
C0154933|ICD9CM|PT|364.70|Adhesions of iris, unspecified
C0154934|ICD9CM|AB|364.73|Goniosynechiae
C0154934|ICD9CM|PT|364.73|Goniosynechiae
C0154935|ICD9CM|PT|364.74|Adhesions and disruptions of pupillary membranes
C0154935|ICD9CM|AB|364.74|Pupillary membranes
C0154936|ICD9CM|AB|364.75|Pupillary abnormalities
C0154936|ICD9CM|PT|364.75|Pupillary abnormalities
C0154937|ICD9CM|PT|364.77|Recession of chamber angle of eye
C0154937|ICD9CM|AB|364.77|Recession, chamber angle
C0154941|ICD9CM|PT|365.02|Anatomical narrow angle borderline glaucoma
C0154941|ICD9CM|AB|365.02|Anatomical narrow angle
C0154944|ICD9CM|PT|365.15|Residual stage of open angle glaucoma
C0154944|ICD9CM|AB|365.15|Residual opn ang glaucma
C0154945|ICD9CM|PT|365.21|Intermittent angle-closure glaucoma
C0154945|ICD9CM|AB|365.21|Intermit angl-clos glauc
C0154946|ICD9CM|PT|365.22|Acute angle-closure glaucoma
C0154946|ICD9CM|AB|365.22|Acute angl-clos glaucoma
C0154947|ICD9CM|PT|365.23|Chronic angle-closure glaucoma
C0154947|ICD9CM|AB|365.23|Chr angle-clos glaucoma
C0154948|ICD9CM|PT|365.24|Residual stage of angle-closure glaucoma
C0154948|ICD9CM|AB|365.24|Residual angl-clos glauc
C0154952|ICD9CM|HT|365.4|Glaucoma associated with congenital anomalies, dystrophies, and systemic syndromes
C0154953|ICD9CM|PT|365.41|Glaucoma associated with chamber angle anomalies
C0154953|ICD9CM|AB|365.41|Glauc w chamb angle anom
C0154954|ICD9CM|PT|365.42|Glaucoma associated with anomalies of iris
C0154954|ICD9CM|AB|365.42|Glaucoma w iris anomaly
C0154955|ICD9CM|PT|365.43|Glaucoma associated with other anterior segment anomalies
C0154955|ICD9CM|AB|365.43|Glauc w ant seg anom NEC
C0154956|ICD9CM|PT|365.44|Glaucoma associated with systemic syndromes
C0154956|ICD9CM|AB|365.44|Glaucoma w systemic synd
C0154959|ICD9CM|PT|365.59|Glaucoma associated with other lens disorders
C0154959|ICD9CM|AB|365.59|Glaucoma w lens dis NEC
C0154960|ICD9CM|HT|365.6|Glaucoma associated with other ocular disorders
C0154961|ICD9CM|PT|365.60|Glaucoma associated with unspecified ocular disorder
C0154961|ICD9CM|AB|365.60|Glauc w ocular dis NOS
C0154964|ICD9CM|PT|365.63|Glaucoma associated with vascular disorders
C0154964|ICD9CM|AB|365.63|Glaucoma w vascular dis
C0154965|ICD9CM|PT|365.64|Glaucoma associated with tumors or cysts
C0154965|ICD9CM|AB|365.64|Glaucoma w tumor or cyst
C0154968|ICD9CM|AB|365.81|Hypersecretion glaucoma
C0154968|ICD9CM|PT|365.81|Hypersecretion glaucoma
C0154970|ICD9CM|HT|366.0|Infantile, juvenile, and presenile cataract
C0154974|ICD9CM|AB|366.03|Cortical cataract
C0154974|ICD9CM|PT|366.03|Cortical, lamellar, or zonular cataract
C0154976|ICD9CM|PT|366.09|Other and combined forms of nonsenile cataract
C0154976|ICD9CM|AB|366.09|Nonsenile cataract NEC
C0154978|ICD9CM|PT|366.13|Anterior subcapsular polar senile cataract
C0154978|ICD9CM|AB|366.13|Ant subcaps senile catar
C0154979|ICD9CM|PT|366.14|Posterior subcapsular polar senile cataract
C0154979|ICD9CM|AB|366.14|Post subcap senile catar
C0154980|ICD9CM|AB|366.15|Cortical senile cataract
C0154980|ICD9CM|PT|366.15|Cortical senile cataract
C0154982|ICD9CM|PT|366.19|Other and combined forms of senile cataract
C0154982|ICD9CM|AB|366.19|Senile cataract NEC
C0154983|ICD9CM|HT|366.2|Traumatic cataract
C0154983|ICD9CM|AB|366.20|Traumatic cataract NOS
C0154983|ICD9CM|PT|366.20|Traumatic cataract, unspecified
C0154984|ICD9CM|PT|366.21|Localized traumatic opacities
C0154984|ICD9CM|AB|366.21|Local traumatic opacity
C0154985|ICD9CM|AB|366.22|Total traumatic cataract
C0154985|ICD9CM|PT|366.22|Total traumatic cataract
C0154986|ICD9CM|PT|366.23|Partially resolved traumatic cataract
C0154986|ICD9CM|AB|366.23|Part resolv traum catar
C0154989|ICD9CM|PT|366.31|Glaucomatous flecks (subcapsular)
C0154989|ICD9CM|AB|366.31|Glaucomatous flecks
C0154990|ICD9CM|PT|366.32|Cataract in inflammatory ocular disorders
C0154990|ICD9CM|AB|366.32|Cataract in inflam dis
C0154992|ICD9CM|PT|366.34|Cataract in degenerative ocular disorders
C0154992|ICD9CM|AB|366.34|Cataract in degen dis
C0154994|ICD9CM|PT|366.44|Cataract associated with other syndromes
C0154994|ICD9CM|HT|366.4|Cataract associated with other disorders
C0154994|ICD9CM|AB|366.44|Cataract w syndrome NEC
C0154995|ICD9CM|AB|366.45|Toxic cataract
C0154995|ICD9CM|PT|366.45|Toxic cataract
C0154996|ICD9CM|PT|366.46|Cataract associated with radiation and other physical influences
C0154996|ICD9CM|AB|366.46|Cataract w radiation
C0154997|ICD9CM|PT|366.52|Other after-cataract, not obscuring vision
C0154997|ICD9CM|AB|366.52|After-cataract NEC
C0154998|ICD9CM|PT|366.53|After-cataract, obscuring vision
C0154998|ICD9CM|AB|366.53|Aftr-catar obscur vision
C0154999|ICD9CM|HT|367.3|Anisometropia and aniseikonia
C0155000|ICD9CM|PT|367.81|Transient refractive change
C0155000|ICD9CM|AB|367.81|Transient refract change
C0155001|ICD9CM|HT|368.1|Subjective visual disturbances
C0155001|ICD9CM|PT|368.10|Subjective visual disturbance, unspecified
C0155001|ICD9CM|AB|368.10|Subj visual disturb NOS
C0155002|ICD9CM|AB|368.11|Sudden visual loss
C0155002|ICD9CM|PT|368.11|Sudden visual loss
C0155003|ICD9CM|AB|368.12|Transient visual loss
C0155003|ICD9CM|PT|368.12|Transient visual loss
C0155004|ICD9CM|PT|368.14|Visual distortions of shape and size
C0155004|ICD9CM|AB|368.14|Distortion of shape/size
C0155005|ICD9CM|PT|368.15|Other visual distortions and entoptic phenomena
C0155005|ICD9CM|AB|368.15|Visual distortions NEC
C0155006|ICD9CM|PT|368.16|Psychophysical visual disturbances
C0155006|ICD9CM|AB|368.16|Psychophysic visual dist
C0155007|ICD9CM|HT|368.3|Other disorders of binocular vision
C0155008|ICD9CM|PT|368.32|Simultaneous visual perception without fusion
C0155008|ICD9CM|AB|368.32|Visual percept w/o fusn
C0155009|ICD9CM|PT|368.33|Fusion with defective stereopsis
C0155009|ICD9CM|AB|368.33|Fusion w def stereopsis
C0155010|ICD9CM|PT|368.34|Abnormal retinal correspondence
C0155010|ICD9CM|AB|368.34|Abn retina correspond
C0155012|ICD9CM|PT|368.45|Generalized visual field contraction or constriction
C0155012|ICD9CM|AB|368.45|Gen visual contraction
C0155015|ICD9CM|AB|368.51|Protan defect
C0155015|ICD9CM|PT|368.51|Protan defect
C0155016|ICD9CM|AB|368.52|Deutan defect
C0155016|ICD9CM|PT|368.52|Deutan defect
C0155017|ICD9CM|AB|368.53|Tritan defect
C0155017|ICD9CM|PT|368.53|Tritan defect
C0155018|ICD9CM|PT|368.55|Acquired color vision deficiencies
C0155018|ICD9CM|AB|368.55|Acq color deficiency
C0155019|ICD9CM|PT|368.63|Abnormal dark adaptation curve
C0155019|ICD9CM|AB|368.63|Abn dark adaptat curve
C0155020|ICD9CM|HT|369|Blindness and low vision
C0155021|ICD9CM|HT|369.0|Profound vision impairment, both eyes
C0155022|ICD9CM|PT|369.01|Better eye: total vision impairment; lesser eye: total vision impairment
C0155022|ICD9CM|AB|369.01|Tot impairment-both eyes
C0155040|ICD9CM|HT|369.2|Moderate or severe vision impairment, both eyes
C0155047|ICD9CM|PT|369.3|Unqualified visual loss, both eyes
C0155047|ICD9CM|AB|369.3|Blindness NOS, both eyes
C0155049|ICD9CM|HT|369.6|Profound vision impairment, one eye
C0155058|ICD9CM|HT|369.7|Moderate or severe vision impairment, one eye
C0155066|ICD9CM|PT|369.8|Unqualified visual loss, one eye
C0155066|ICD9CM|AB|369.8|Visual loss, one eye NOS
C0155067|ICD9CM|AB|370.01|Marginal corneal ulcer
C0155067|ICD9CM|PT|370.01|Marginal corneal ulcer
C0155068|ICD9CM|AB|370.02|Ring corneal ulcer
C0155068|ICD9CM|PT|370.02|Ring corneal ulcer
C0155069|ICD9CM|AB|370.03|Central corneal ulcer
C0155069|ICD9CM|PT|370.03|Central corneal ulcer
C0155070|ICD9CM|AB|370.04|Hypopyon ulcer
C0155070|ICD9CM|PT|370.04|Hypopyon ulcer
C0155071|ICD9CM|AB|370.05|Mycotic corneal ulcer
C0155071|ICD9CM|PT|370.05|Mycotic corneal ulcer
C0155072|ICD9CM|AB|370.07|Mooren's ulcer
C0155072|ICD9CM|PT|370.07|Mooren's ulcer
C0155073|ICD9CM|HT|370.2|Superficial keratitis without conjunctivitis
C0155074|ICD9CM|PT|370.20|Superficial keratitis, unspecified
C0155074|ICD9CM|AB|370.20|Superfic keratitis NOS
C0155076|ICD9CM|AB|370.22|Macular keratitis
C0155076|ICD9CM|PT|370.22|Macular keratitis
C0155077|ICD9CM|AB|370.23|Filamentary keratitis
C0155077|ICD9CM|PT|370.23|Filamentary keratitis
C0155078|ICD9CM|AB|370.24|Photokeratitis
C0155078|ICD9CM|PT|370.24|Photokeratitis
C0155079|ICD9CM|HT|370.3|Certain types of keratoconjunctivitis
C0155080|ICD9CM|PT|370.31|Phlyctenular keratoconjunctivitis
C0155080|ICD9CM|AB|370.31|Phlycten keratoconjunct
C0155081|ICD9CM|PT|370.32|Limbar and corneal involvement in vernal conjunctivitis
C0155081|ICD9CM|AB|370.32|Limbar keratoconjunctiv
C0155082|ICD9CM|PT|370.33|Keratoconjunctivitis sicca, not specified as Sjogren's
C0155082|ICD9CM|AB|370.33|Keratoconjunctivit sicca
C0155084|ICD9CM|PT|370.35|Neurotrophic keratoconjunctivitis
C0155084|ICD9CM|AB|370.35|Neurotroph keratoconjunc
C0155085|ICD9CM|HT|370.4|Other and unspecified keratoconjunctivitis
C0155086|ICD9CM|PT|370.44|Keratitis or keratoconjunctivitis in exanthema
C0155086|ICD9CM|AB|370.44|Keratitis in exanthema
C0155087|ICD9CM|HT|370.5|Interstitial and deep keratitis
C0155088|ICD9CM|PT|370.50|Interstitial keratitis, unspecified
C0155088|ICD9CM|AB|370.50|Interstit keratitis NOS
C0155089|ICD9CM|PT|370.52|Diffuse interstitial keratitis
C0155089|ICD9CM|AB|370.52|Diffus interstit keratit
C0155090|ICD9CM|AB|370.54|Sclerosing keratitis
C0155090|ICD9CM|PT|370.54|Sclerosing keratitis
C0155091|ICD9CM|AB|370.55|Corneal abscess
C0155091|ICD9CM|PT|370.55|Corneal abscess
C0155092|ICD9CM|PT|370.59|Other interstitial and deep keratitis
C0155092|ICD9CM|AB|370.59|Interstit keratitis NEC
C0155093|ICD9CM|PT|370.61|Localized vascularization of cornea
C0155093|ICD9CM|AB|370.61|Local vasculariza cornea
C0155094|ICD9CM|AB|370.62|Corneal pannus
C0155094|ICD9CM|PT|370.62|Pannus (corneal)
C0155095|ICD9CM|PT|370.63|Deep vascularization of cornea
C0155095|ICD9CM|AB|370.63|Deep vasculariza cornea
C0155096|ICD9CM|AB|370.64|Corneal ghost vessels
C0155096|ICD9CM|PT|370.64|Ghost vessels (corneal)
C0155097|ICD9CM|HT|371|Corneal opacity and other disorders of cornea
C0155098|ICD9CM|HT|371.0|Corneal scars and opacities
C0155099|ICD9CM|AB|371.01|Minor opacity of cornea
C0155099|ICD9CM|PT|371.01|Minor opacity of cornea
C0155100|ICD9CM|PT|371.02|Peripheral opacity of cornea
C0155100|ICD9CM|AB|371.02|Periph opacity of cornea
C0155102|ICD9CM|AB|371.05|Phthisical cornea
C0155102|ICD9CM|PT|371.05|Phthisical cornea
C0155104|ICD9CM|PT|371.11|Anterior corneal pigmentations
C0155104|ICD9CM|AB|371.11|Ant cornea pigmentation
C0155105|ICD9CM|PT|371.12|Stromal corneal pigmentations
C0155105|ICD9CM|AB|371.12|Stromal cornea pigment
C0155106|ICD9CM|PT|371.13|Posterior corneal pigmentations
C0155106|ICD9CM|AB|371.13|Post cornea pigmentation
C0155107|ICD9CM|PT|371.15|Other corneal deposits associated with metabolic disorders
C0155107|ICD9CM|AB|371.15|Oth deposit w metab dis
C0155108|ICD9CM|PT|371.16|Argentous corneal deposits
C0155108|ICD9CM|AB|371.16|Argentous cornea deposit
C0155109|ICD9CM|AB|371.21|Idiopathic corneal edema
C0155109|ICD9CM|PT|371.21|Idiopathic corneal edema
C0155110|ICD9CM|AB|371.22|Secondary corneal edema
C0155110|ICD9CM|PT|371.22|Secondary corneal edema
C0155111|ICD9CM|AB|371.23|Bullous keratopathy
C0155111|ICD9CM|PT|371.23|Bullous keratopathy
C0155114|ICD9CM|HT|371.3|Changes of corneal membranes
C0155114|ICD9CM|PT|371.30|Corneal membrane change, unspecified
C0155114|ICD9CM|AB|371.30|Cornea memb change NOS
C0155115|ICD9CM|PT|371.31|Folds and rupture of bowman's membrane
C0155115|ICD9CM|AB|371.31|Fold of bowman membrane
C0155116|ICD9CM|PT|371.32|Folds in descemet's membrane
C0155116|ICD9CM|AB|371.32|Fold in descemet membran
C0155117|ICD9CM|PT|371.33|Rupture in descemet's membrane
C0155117|ICD9CM|AB|371.33|Rupture descemet membran
C0155118|ICD9CM|HT|371.4|Corneal degenerations
C0155118|ICD9CM|AB|371.40|Corneal degeneration NOS
C0155118|ICD9CM|PT|371.40|Corneal degeneration, unspecified
C0155119|ICD9CM|PT|371.42|Recurrent erosion of cornea
C0155119|ICD9CM|AB|371.42|Recurrent cornea erosion
C0155120|ICD9CM|AB|371.43|Band-shaped keratopathy
C0155120|ICD9CM|PT|371.43|Band-shaped keratopathy
C0155121|ICD9CM|PT|371.44|Other calcerous degenerations of cornea
C0155121|ICD9CM|AB|371.44|Calcer cornea degen NEC
C0155122|ICD9CM|PT|371.46|Nodular degeneration of cornea
C0155122|ICD9CM|AB|371.46|Nodular cornea degen
C0155123|ICD9CM|PT|371.48|Peripheral degenerations of cornea
C0155123|ICD9CM|AB|371.48|Peripheral cornea degen
C0155124|ICD9CM|PT|371.49|Other corneal degenerations
C0155124|ICD9CM|AB|371.49|Cornea degeneration NEC
C0155126|ICD9CM|PT|371.52|Other anterior corneal dystrophies
C0155126|ICD9CM|AB|371.52|Ant cornea dystrophy NEC
C0155127|ICD9CM|PT|371.54|Lattice corneal dystrophy
C0155127|ICD9CM|AB|371.54|Lattice cornea dystrophy
C0155128|ICD9CM|PT|371.56|Other stromal corneal dystrophies
C0155128|ICD9CM|AB|371.56|Strom cornea dystrph NEC
C0155130|ICD9CM|PT|371.58|Other posterior corneal dystrophies
C0155130|ICD9CM|AB|371.58|Post cornea dystrphy NEC
C0155131|ICD9CM|PT|371.61|Keratoconus, stable condition
C0155131|ICD9CM|AB|371.61|Keratoconus, stable
C0155133|ICD9CM|HT|371.7|Other corneal deformities
C0155135|ICD9CM|AB|371.71|Corneal ectasia
C0155135|ICD9CM|PT|371.71|Corneal ectasia
C0155136|ICD9CM|AB|371.72|Descemetocele
C0155136|ICD9CM|PT|371.72|Descemetocele
C0155137|ICD9CM|HT|371.8|Other corneal disorders
C0155137|ICD9CM|PT|371.89|Other corneal disorders
C0155137|ICD9CM|AB|371.89|Corneal disorder NEC
C0155138|ICD9CM|PT|371.81|Corneal anesthesia and hypoesthesia
C0155138|ICD9CM|AB|371.81|Corneal anesthesia
C0155141|ICD9CM|HT|372.0|Acute conjunctivitis
C0155141|ICD9CM|AB|372.00|Acute conjunctivitis NOS
C0155141|ICD9CM|PT|372.00|Acute conjunctivitis, unspecified
C0155142|ICD9CM|PT|372.01|Serous conjunctivitis, except viral
C0155142|ICD9CM|AB|372.01|Serous conjunctivitis
C0155143|ICD9CM|PT|372.02|Acute follicular conjunctivitis
C0155143|ICD9CM|AB|372.02|Ac follic conjunctivitis
C0155144|ICD9CM|PT|372.04|Pseudomembranous conjunctivitis
C0155144|ICD9CM|AB|372.04|Pseudomemb conjunctivit
C0155145|ICD9CM|HT|372.1|Chronic conjunctivitis
C0155145|ICD9CM|PT|372.10|Chronic conjunctivitis, unspecified
C0155145|ICD9CM|AB|372.10|Chr conjunctivitis NOS
C0155146|ICD9CM|PT|372.11|Simple chronic conjunctivitis
C0155146|ICD9CM|AB|372.11|Simpl chr conjunctivitis
C0155147|ICD9CM|PT|372.12|Chronic follicular conjunctivitis
C0155147|ICD9CM|AB|372.12|Chr follic conjunctivit
C0155148|ICD9CM|AB|372.15|Parasitic conjunctivitis
C0155148|ICD9CM|PT|372.15|Parasitic conjunctivitis
C0155149|ICD9CM|PT|372.21|Angular blepharoconjunctivitis
C0155149|ICD9CM|AB|372.21|Angular blepharoconjunct
C0155150|ICD9CM|PT|372.22|Contact blepharoconjunctivitis
C0155150|ICD9CM|AB|372.22|Contact blepharoconjunct
C0155152|ICD9CM|AB|372.31|Rosacea conjunctivitis
C0155152|ICD9CM|PT|372.31|Rosacea conjunctivitis
C0155153|ICD9CM|PT|372.33|Conjunctivitis in mucocutaneous disease
C0155153|ICD9CM|AB|372.33|Mucocutan dis conjunctiv
C0155154|ICD9CM|PT|372.41|Peripheral pterygium, stationary
C0155154|ICD9CM|AB|372.41|Periph station pterygium
C0155155|ICD9CM|PT|372.42|Peripheral pterygium, progressive
C0155155|ICD9CM|AB|372.42|Periph progess pterygium
C0155156|ICD9CM|AB|372.43|Central pterygium
C0155156|ICD9CM|PT|372.43|Central pterygium
C0155157|ICD9CM|AB|372.44|Double pterygium
C0155157|ICD9CM|PT|372.44|Double pterygium
C0155158|ICD9CM|AB|372.45|Recurrent pterygium
C0155158|ICD9CM|PT|372.45|Recurrent pterygium
C0155159|ICD9CM|HT|372.5|Conjunctival degenerations and deposits
C0155160|ICD9CM|PT|372.50|Conjunctival degeneration, unspecified
C0155160|ICD9CM|AB|372.50|Conjunctival degen NOS
C0155161|ICD9CM|AB|372.52|Pseudopterygium
C0155161|ICD9CM|PT|372.52|Pseudopterygium
C0155162|ICD9CM|AB|372.54|Conjunctival concretions
C0155162|ICD9CM|PT|372.54|Conjunctival concretions
C0155163|ICD9CM|PT|372.55|Conjunctival pigmentations
C0155163|ICD9CM|AB|372.55|Conjunctiva pigmentation
C0155164|ICD9CM|HT|372.6|Conjunctival scars
C0155164|ICD9CM|AB|372.64|Scarring of conjunctiva
C0155164|ICD9CM|PT|372.64|Scarring of conjunctiva
C0155165|ICD9CM|AB|372.61|Granuloma of conjunctiva
C0155165|ICD9CM|PT|372.61|Granuloma of conjunctiva
C0155166|ICD9CM|PT|372.62|Localized adhesions and strands of conjunctiva
C0155166|ICD9CM|AB|372.62|Local conjunctiva adhes
C0155168|ICD9CM|HT|372.7|Conjunctival vascular disorders and cysts
C0155170|ICD9CM|AB|372.75|Conjunctival cysts
C0155170|ICD9CM|PT|372.75|Conjunctival cysts
C0155171|ICD9CM|HT|372.8|Other disorders of conjunctiva
C0155171|ICD9CM|PT|372.89|Other disorders of conjunctiva
C0155171|ICD9CM|AB|372.89|Conjunctiva disorder NEC
C0155173|ICD9CM|AB|373.01|Ulcerative blepharitis
C0155173|ICD9CM|PT|373.01|Ulcerative blepharitis
C0155174|ICD9CM|AB|373.02|Squamous blepharitis
C0155174|ICD9CM|PT|373.02|Squamous blepharitis
C0155175|ICD9CM|AB|373.13|Abscess of eyelid
C0155175|ICD9CM|PT|373.13|Abscess of eyelid
C0155176|ICD9CM|HT|373.3|Noninfectious dermatoses of eyelid
C0155177|ICD9CM|PT|373.31|Eczematous dermatitis of eyelid
C0155177|ICD9CM|AB|373.31|Eczem dermatitis eyelid
C0155178|ICD9CM|PT|373.32|Contact and allergic dermatitis of eyelid
C0155178|ICD9CM|AB|373.32|Contact dermatit eyelid
C0155179|ICD9CM|AB|373.33|Xeroderma of eyelid
C0155179|ICD9CM|PT|373.33|Xeroderma of eyelid
C0155180|ICD9CM|PT|373.34|Discoid lupus erythematosus of eyelid
C0155180|ICD9CM|AB|373.34|Disc lup erythematos lid
C0155181|ICD9CM|PT|373.4|Infective dermatitis of eyelid of types resulting in deformity
C0155181|ICD9CM|AB|373.4|Infect derm lid w deform
C0155182|ICD9CM|PT|373.5|Other infective dermatitis of eyelid
C0155182|ICD9CM|AB|373.5|Infec dermatitis lid NEC
C0155183|ICD9CM|PT|373.6|Parasitic infestation of eyelid
C0155183|ICD9CM|AB|373.6|Parasitic infest eyelid
C0155184|ICD9CM|PT|373.8|Other inflammations of eyelids
C0155184|ICD9CM|AB|373.8|Inflammation eyelid NEC
C0155186|ICD9CM|HT|374.8|Other disorders of eyelid
C0155186|ICD9CM|PT|374.89|Other disorders of eyelid
C0155186|ICD9CM|HT|374|Other disorders of eyelids
C0155186|ICD9CM|AB|374.89|Disorders of eyelid NEC
C0155188|ICD9CM|AB|374.01|Senile entropion
C0155188|ICD9CM|PT|374.01|Senile entropion
C0155189|ICD9CM|AB|374.02|Mechanical entropion
C0155189|ICD9CM|PT|374.02|Mechanical entropion
C0155190|ICD9CM|AB|374.03|Spastic entropion
C0155190|ICD9CM|PT|374.03|Spastic entropion
C0155191|ICD9CM|AB|374.04|Cicatricial entropion
C0155191|ICD9CM|PT|374.04|Cicatricial entropion
C0155193|ICD9CM|AB|374.11|Senile ectropion
C0155193|ICD9CM|PT|374.11|Senile ectropion
C0155194|ICD9CM|AB|374.12|Mechanical ectropion
C0155194|ICD9CM|PT|374.12|Mechanical ectropion
C0155195|ICD9CM|AB|374.13|Spastic ectropion
C0155195|ICD9CM|PT|374.13|Spastic ectropion
C0155196|ICD9CM|AB|374.14|Cicatricial ectropion
C0155196|ICD9CM|PT|374.14|Cicatricial ectropion
C0155197|ICD9CM|AB|374.21|Paralytic lagophthalmos
C0155197|ICD9CM|PT|374.21|Paralytic lagophthalmos
C0155198|ICD9CM|AB|374.22|Mechanical lagophthalmos
C0155198|ICD9CM|PT|374.22|Mechanical lagophthalmos
C0155199|ICD9CM|PT|374.23|Cicatricial lagophthalmos
C0155199|ICD9CM|AB|374.23|Cicatricial lagophthalm
C0155201|ICD9CM|AB|374.32|Myogenic ptosis
C0155201|ICD9CM|PT|374.32|Myogenic ptosis
C0155202|ICD9CM|AB|374.33|Mechanical ptosis
C0155202|ICD9CM|PT|374.33|Mechanical ptosis
C0155203|ICD9CM|HT|374.4|Other disorders affecting eyelid function
C0155204|ICD9CM|AB|374.41|Lid retraction or lag
C0155204|ICD9CM|PT|374.41|Lid retraction or lag
C0155206|ICD9CM|PT|374.44|Sensory disorders of eyelid
C0155206|ICD9CM|AB|374.44|Sensory disorders, lid
C0155207|ICD9CM|PT|374.45|Other sensorimotor disorders of eyelid
C0155207|ICD9CM|AB|374.45|Sensormotr disor lid NEC
C0155208|ICD9CM|HT|374.5|Degenerative disorders of eyelid and periocular area
C0155209|ICD9CM|PT|374.50|Degenerative disorder of eyelid, unspecified
C0155209|ICD9CM|AB|374.50|Degen disorder NOS, lid
C0155210|ICD9CM|PT|374.51|Xanthelasma of eyelid
C0155210|ICD9CM|AB|374.51|Xanthelasma
C0155211|ICD9CM|PT|374.52|Hyperpigmentation of eyelid
C0155211|ICD9CM|AB|374.52|Hyperpigmentation lid
C0155212|ICD9CM|PT|374.53|Hypopigmentation of eyelid
C0155212|ICD9CM|AB|374.53|Hypopigmentation lid
C0155213|ICD9CM|AB|374.54|Hypertrichosis of eyelid
C0155213|ICD9CM|PT|374.54|Hypertrichosis of eyelid
C0155214|ICD9CM|AB|374.55|Hypotrichosis of eyelid
C0155214|ICD9CM|PT|374.55|Hypotrichosis of eyelid
C0155215|ICD9CM|PT|374.56|Other degenerative disorders of skin affecting eyelid
C0155215|ICD9CM|AB|374.56|Degen dis eyelid NEC
C0155216|ICD9CM|AB|374.81|Hemorrhage of eyelid
C0155216|ICD9CM|PT|374.81|Hemorrhage of eyelid
C0155217|ICD9CM|AB|374.83|Elephantiasis of eyelid
C0155217|ICD9CM|PT|374.83|Elephantiasis of eyelid
C0155218|ICD9CM|AB|374.84|Cysts of eyelids
C0155218|ICD9CM|PT|374.84|Cysts of eyelids
C0155219|ICD9CM|PT|374.85|Vascular anomalies of eyelid
C0155219|ICD9CM|AB|374.85|Vascular anomaly, eyelid
C0155223|ICD9CM|HT|375.0|Dacryoadenitis
C0155223|ICD9CM|AB|375.00|Dacryoadenitis NOS
C0155223|ICD9CM|PT|375.00|Dacryoadenitis, unspecified
C0155224|ICD9CM|AB|375.02|Chronic dacryoadenitis
C0155224|ICD9CM|PT|375.02|Chronic dacryoadenitis
C0155226|ICD9CM|HT|375.1|Other disorders of lacrimal gland
C0155227|ICD9CM|AB|375.11|Dacryops
C0155227|ICD9CM|PT|375.11|Dacryops
C0155228|ICD9CM|PT|375.12|Other lacrimal cysts and cystic degeneration
C0155228|ICD9CM|AB|375.12|Lacrimal gland cyst NEC
C0155229|ICD9CM|AB|375.13|Primary lacrimal atrophy
C0155229|ICD9CM|PT|375.13|Primary lacrimal atrophy
C0155231|ICD9CM|PT|375.16|Dislocation of lacrimal gland
C0155231|ICD9CM|AB|375.16|Lacrimal gland dislocat
C0155233|ICD9CM|PT|375.21|Epiphora due to excess lacrimation
C0155233|ICD9CM|AB|375.21|Epiphora d/t excess tear
C0155234|ICD9CM|PT|375.22|Epiphora due to insufficient drainage
C0155234|ICD9CM|AB|375.22|Epiphora d/t insuf drain
C0155237|ICD9CM|AB|375.32|Acute dacryocystitis
C0155237|ICD9CM|PT|375.32|Acute dacryocystitis
C0155238|ICD9CM|PT|375.33|Phlegmonous dacryocystitis
C0155238|ICD9CM|AB|375.33|Phlegmon dacryocystitis
C0155239|ICD9CM|HT|375.4|Chronic inflammation of lacrimal passages
C0155240|ICD9CM|AB|375.41|Chronic canaliculitis
C0155240|ICD9CM|PT|375.41|Chronic canaliculitis
C0155241|ICD9CM|AB|375.43|Lacrimal mucocele
C0155241|ICD9CM|PT|375.43|Lacrimal mucocele
C0155242|ICD9CM|HT|375.5|Stenosis and insufficiency of lacrimal passages
C0155243|ICD9CM|PT|375.51|Eversion of lacrimal punctum
C0155243|ICD9CM|AB|375.51|Lacriml punctum eversion
C0155244|ICD9CM|PT|375.52|Stenosis of lacrimal punctum
C0155244|ICD9CM|AB|375.52|Lacriml punctum stenosis
C0155245|ICD9CM|PT|375.53|Stenosis of lacrimal canaliculi
C0155245|ICD9CM|AB|375.53|Lacrim canalic stenosis
C0155246|ICD9CM|PT|375.54|Stenosis of lacrimal sac
C0155246|ICD9CM|AB|375.54|Lacrimal sac stenosis
C0155248|ICD9CM|PT|375.56|Stenosis of nasolacrimal duct, acquired
C0155248|ICD9CM|AB|375.56|Acq nasolacrml stenosis
C0155249|ICD9CM|AB|375.57|Dacryolith
C0155249|ICD9CM|PT|375.57|Dacryolith
C0155250|ICD9CM|HT|375.6|Other changes of lacrimal passages
C0155250|ICD9CM|PT|375.69|Other changes of lacrimal passages
C0155250|ICD9CM|AB|375.69|Lacrim passge change NEC
C0155251|ICD9CM|AB|375.61|Lacrimal fistula
C0155251|ICD9CM|PT|375.61|Lacrimal fistula
C0155252|ICD9CM|HT|375.8|Other disorders of lacrimal system
C0155252|ICD9CM|PT|375.89|Other disorders of lacrimal system
C0155252|ICD9CM|AB|375.89|Lacrimal syst dis NEC
C0155253|ICD9CM|PT|375.81|Granuloma of lacrimal passages
C0155253|ICD9CM|AB|375.81|Lacrim passage granuloma
C0155256|ICD9CM|HT|376.0|Acute inflammation of orbit
C0155256|ICD9CM|PT|376.00|Acute inflammation of orbit, unspecified
C0155256|ICD9CM|AB|376.00|Acute inflam NOS, orbit
C0155257|ICD9CM|AB|376.02|Orbital periostitis
C0155257|ICD9CM|PT|376.02|Orbital periostitis
C0155258|ICD9CM|AB|376.03|Orbital osteomyelitis
C0155258|ICD9CM|PT|376.03|Orbital osteomyelitis
C0155259|ICD9CM|AB|376.04|Orbital tenonitis
C0155259|ICD9CM|PT|376.04|Orbital tenonitis
C0155261|ICD9CM|HT|376.1|Chronic inflammatory disorders of orbit
C0155261|ICD9CM|PT|376.10|Chronic inflammation of orbit, unspecified
C0155261|ICD9CM|AB|376.10|Chr inflam NOS, orbit
C0155262|ICD9CM|AB|376.11|Orbital granuloma
C0155262|ICD9CM|PT|376.11|Orbital granuloma
C0155263|ICD9CM|PT|376.13|Parasitic infestation of orbit
C0155263|ICD9CM|AB|376.13|Parasite infest, orbit
C0155264|ICD9CM|HT|376.2|Endocrine exophthalmos
C0155265|ICD9CM|AB|376.21|Thyrotoxic exophthalmos
C0155265|ICD9CM|PT|376.21|Thyrotoxic exophthalmos
C0155266|ICD9CM|HT|376.3|Other exophthalmic conditions
C0155267|ICD9CM|AB|376.31|Constant exophthalmos
C0155267|ICD9CM|PT|376.31|Constant exophthalmos
C0155268|ICD9CM|AB|376.32|Orbital hemorrhage
C0155268|ICD9CM|PT|376.32|Orbital hemorrhage
C0155270|ICD9CM|PT|376.34|Intermittent exophthalmos
C0155270|ICD9CM|AB|376.34|Intermittnt exophthalmos
C0155271|ICD9CM|AB|376.35|Pulsating exophthalmos
C0155271|ICD9CM|PT|376.35|Pulsating exophthalmos
C0155272|ICD9CM|PT|376.36|Lateral displacement of globe
C0155272|ICD9CM|AB|376.36|Lateral globe displacmnt
C0155275|ICD9CM|AB|376.42|Exostosis of orbit
C0155275|ICD9CM|PT|376.42|Exostosis of orbit
C0155276|ICD9CM|PT|376.43|Local deformities of orbit due to bone disease
C0155276|ICD9CM|AB|376.43|Orbt deform d/t bone dis
C0155277|ICD9CM|PT|376.44|Orbital deformities associated with craniofacial deformities
C0155277|ICD9CM|AB|376.44|Craniofacial-orbit defor
C0155278|ICD9CM|AB|376.45|Atrophy of orbit
C0155278|ICD9CM|PT|376.45|Atrophy of orbit
C0155279|ICD9CM|AB|376.46|Enlargement of orbit
C0155279|ICD9CM|PT|376.46|Enlargement of orbit
C0155280|ICD9CM|PT|376.47|Deformity of orbit due to trauma or surgery
C0155280|ICD9CM|AB|376.47|Orbit deform d/t trauma
C0155281|ICD9CM|PT|376.51|Enophthalmos due to atrophy of orbital tissue
C0155281|ICD9CM|AB|376.51|Enophth d/t orbit atrphy
C0155282|ICD9CM|PT|376.52|Enophthalmos due to trauma or surgery
C0155282|ICD9CM|AB|376.52|Enophthalmos d/t trauma
C0155283|ICD9CM|PT|376.6|Retained (old) foreign body following penetrating wound of orbit
C0155283|ICD9CM|AB|376.6|Old foreign body, orbit
C0155284|ICD9CM|HT|376.8|Other orbital disorders
C0155285|ICD9CM|AB|376.81|Orbital cysts
C0155285|ICD9CM|PT|376.81|Orbital cysts
C0155286|ICD9CM|PT|376.82|Myopathy of extraocular muscles
C0155286|ICD9CM|AB|376.82|Extraocul muscl myopathy
C0155288|ICD9CM|PT|377.01|Papilledema associated with increased intracranial pressure
C0155288|ICD9CM|AB|377.01|Papilledema w incr press
C0155290|ICD9CM|PT|377.03|Papilledema associated with retinal disorder
C0155290|ICD9CM|AB|377.03|Papilledema w retina dis
C0155291|ICD9CM|AB|377.11|Primary optic atrophy
C0155291|ICD9CM|PT|377.11|Primary optic atrophy
C0155292|ICD9CM|PT|377.12|Postinflammatory optic atrophy
C0155292|ICD9CM|AB|377.12|Postinflam optic atrophy
C0155293|ICD9CM|PT|377.13|Optic atrophy associated with retinal dystrophies
C0155293|ICD9CM|AB|377.13|Optic atrph w retin dyst
C0155295|ICD9CM|AB|377.15|Partial optic atrophy
C0155295|ICD9CM|PT|377.15|Partial optic atrophy
C0155296|ICD9CM|HT|377.2|Other disorders of optic disc
C0155298|ICD9CM|PT|377.22|Crater-like holes of optic disc
C0155298|ICD9CM|AB|377.22|Crater-like hole op disc
C0155299|ICD9CM|AB|377.23|Coloboma of optic disc
C0155299|ICD9CM|PT|377.23|Coloboma of optic disc
C0155300|ICD9CM|AB|377.24|Pseudopapilledema
C0155300|ICD9CM|PT|377.24|Pseudopapilledema
C0155301|ICD9CM|PT|377.32|Retrobulbar neuritis (acute)
C0155301|ICD9CM|AB|377.32|Retrobulbar neuritis
C0155302|ICD9CM|PT|377.33|Nutritional optic neuropathy
C0155302|ICD9CM|AB|377.33|Nutrition optc neuropthy
C0155303|ICD9CM|AB|377.34|Toxic optic neuropathy
C0155303|ICD9CM|PT|377.34|Toxic optic neuropathy
C0155304|ICD9CM|HT|377.4|Other disorders of optic nerve
C0155304|ICD9CM|PT|377.49|Other disorders of optic nerve
C0155304|ICD9CM|AB|377.49|Optic nerve disorder NEC
C0155305|ICD9CM|PT|377.41|Ischemic optic neuropathy
C0155305|ICD9CM|AB|377.41|Ischemic optic neuropthy
C0155306|ICD9CM|PT|377.42|Hemorrhage in optic nerve sheaths
C0155306|ICD9CM|AB|377.42|Optic nerve sheath hemor
C0155307|ICD9CM|HT|377.5|Disorders of optic chiasm
C0155308|ICD9CM|PT|377.51|Disorders of optic chiasm associated with pituitary neoplasms and disorders
C0155308|ICD9CM|AB|377.51|Opt chiasm w pituit dis
C0155311|ICD9CM|PT|377.54|Disorders of optic chiasm associated with inflammatory disorders
C0155311|ICD9CM|AB|377.54|Op chiasm dis w infl dis
C0155312|ICD9CM|HT|377.6|Disorders of other visual pathways
C0155313|ICD9CM|PT|377.61|Disorders of other visual pathways associated with neoplasms
C0155313|ICD9CM|AB|377.61|Vis path dis w neoplasms
C0155314|ICD9CM|PT|377.62|Disorders of other visual pathways associated with vascular disorders
C0155314|ICD9CM|AB|377.62|Vis path dis w vasc dis
C0155315|ICD9CM|PT|377.63|Disorders of other visual pathways associated with inflammatory disorders
C0155315|ICD9CM|AB|377.63|Vis path dis w infl dis
C0155320|ICD9CM|AB|377.75|Cortical blindness
C0155320|ICD9CM|PT|377.75|Cortical blindness
C0155322|ICD9CM|PT|378.02|Monocular esotropia with A pattern
C0155322|ICD9CM|AB|378.02|Monoc esotrop w a pattrn
C0155323|ICD9CM|PT|378.03|Monocular esotropia with V pattern
C0155323|ICD9CM|AB|378.03|Monoc esotrop w v pattrn
C0155324|ICD9CM|PT|378.04|Monocular esotropia with other noncomitancies
C0155324|ICD9CM|AB|378.04|Monoc esotrop w x/y pat
C0155325|ICD9CM|PT|378.06|Alternating esotropia with A pattern
C0155325|ICD9CM|AB|378.06|Alt esotropia w a pattrn
C0155326|ICD9CM|PT|378.07|Alternating esotropia with V pattern
C0155326|ICD9CM|AB|378.07|Alt esotropia w v pattrn
C0155327|ICD9CM|PT|378.08|Alternating esotropia with other noncomitancies
C0155327|ICD9CM|AB|378.08|Alt esotrop w x/y pattrn
C0155328|ICD9CM|PT|378.12|Monocular exotropia with A pattern
C0155328|ICD9CM|AB|378.12|Monoc exotrop w a pattrn
C0155329|ICD9CM|PT|378.13|Monocular exotropia with V pattern
C0155329|ICD9CM|AB|378.13|Monoc exotrop w v pattrn
C0155330|ICD9CM|PT|378.14|Monocular exotropia with other noncomitancies
C0155330|ICD9CM|AB|378.14|Monoc exotrop w x/y pat
C0155331|ICD9CM|PT|378.16|Alternating exotropia with A pattern
C0155331|ICD9CM|AB|378.16|Alt exotropia w a pattrn
C0155332|ICD9CM|PT|378.17|Alternating exotropia with V pattern
C0155332|ICD9CM|AB|378.17|Alt exotropia w v pattrn
C0155333|ICD9CM|PT|378.18|Alternating exotropia with other noncomitancies
C0155333|ICD9CM|AB|378.18|Alt exotrop w x/y pattrn
C0155334|ICD9CM|HT|378.3|Other and unspecified heterotropia
C0155336|ICD9CM|PT|378.35|Accommodative component in esotropia
C0155336|ICD9CM|AB|378.35|Accommodative esotropia
C0155338|ICD9CM|AB|378.56|Total ophthalmoplegia
C0155338|ICD9CM|PT|378.56|Total ophthalmoplegia
C0155339|ICD9CM|PT|378.61|Brown's (tendon) sheath syndrome
C0155339|ICD9CM|AB|378.61|Brown's sheath syndrome
C0155340|ICD9CM|PT|378.62|Mechanical strabismus from other musculofascial disorders
C0155340|ICD9CM|AB|378.62|Mech strab d/t muscl dis
C0155341|ICD9CM|PT|378.63|Limited duction associated with other conditions
C0155341|ICD9CM|AB|378.63|Mech strab w oth conditn
C0155342|ICD9CM|PT|378.73|Strabismus in other neuromuscular disorders
C0155342|ICD9CM|AB|378.73|Neuromuscle dis strabism
C0155343|ICD9CM|HT|378.8|Other disorders of binocular eye movements
C0155344|ICD9CM|AB|378.82|Spasm of conjugate gaze
C0155344|ICD9CM|PT|378.82|Spasm of conjugate gaze
C0155345|ICD9CM|PT|378.83|Convergence insufficiency or palsy
C0155345|ICD9CM|AB|378.83|Convergenc insufficiency
C0155346|ICD9CM|PT|378.84|Convergence excess or spasm
C0155346|ICD9CM|AB|378.84|Convergence excess
C0155347|ICD9CM|AB|378.85|Anomalies of divergence
C0155347|ICD9CM|PT|378.85|Anomalies of divergence
C0155351|ICD9CM|PT|379.01|Episcleritis periodica fugax
C0155351|ICD9CM|AB|379.01|Episclerit periodic fugx
C0155352|ICD9CM|AB|379.02|Nodular episcleritis
C0155352|ICD9CM|PT|379.02|Nodular episcleritis
C0155353|ICD9CM|AB|379.03|Anterior scleritis
C0155353|ICD9CM|PT|379.03|Anterior scleritis
C0155354|ICD9CM|AB|379.04|Scleromalacia perforans
C0155354|ICD9CM|PT|379.04|Scleromalacia perforans
C0155355|ICD9CM|PT|379.05|Scleritis with corneal involvement
C0155355|ICD9CM|AB|379.05|Scleritis w cornea invol
C0155356|ICD9CM|AB|379.06|Brawny scleritis
C0155356|ICD9CM|PT|379.06|Brawny scleritis
C0155357|ICD9CM|AB|379.07|Posterior scleritis
C0155357|ICD9CM|PT|379.07|Posterior scleritis
C0155358|ICD9CM|PT|379.19|Other disorders of sclera
C0155358|ICD9CM|HT|379.1|Other disorders of sclera
C0155358|ICD9CM|AB|379.19|Disorder of sclera NEC
C0155360|ICD9CM|AB|379.12|Staphyloma posticum
C0155360|ICD9CM|PT|379.12|Staphyloma posticum
C0155361|ICD9CM|AB|379.13|Equatorial staphyloma
C0155361|ICD9CM|PT|379.13|Equatorial staphyloma
C0155362|ICD9CM|PT|379.14|Anterior staphyloma, localized
C0155362|ICD9CM|AB|379.14|Local anterior staphylma
C0155363|ICD9CM|AB|379.15|Ring staphyloma
C0155363|ICD9CM|PT|379.15|Ring staphyloma
C0155364|ICD9CM|PT|379.16|Other degenerative disorders of sclera
C0155364|ICD9CM|AB|379.16|Scleral degen dis NEC
C0155365|ICD9CM|HT|379.2|Disorders of vitreous body
C0155366|ICD9CM|AB|379.21|Vitreous degeneration
C0155366|ICD9CM|PT|379.21|Vitreous degeneration
C0155367|ICD9CM|PT|379.22|Crystalline deposits in vitreous
C0155367|ICD9CM|AB|379.22|Crystal deposit vitreous
C0155368|ICD9CM|PT|379.25|Vitreous membranes and strands
C0155368|ICD9CM|AB|379.25|Vitreous membranes
C0155369|ICD9CM|AB|379.26|Vitreous prolapse
C0155369|ICD9CM|PT|379.26|Vitreous prolapse
C0155370|ICD9CM|PT|379.29|Other disorders of vitreous
C0155370|ICD9CM|AB|379.29|Vitreous disorders NEC
C0155371|ICD9CM|HT|379.3|Aphakia and other disorders of lens
C0155372|ICD9CM|PT|379.33|Anterior dislocation of lens
C0155372|ICD9CM|AB|379.33|Ant dislocation of lens
C0155373|ICD9CM|PT|379.34|Posterior dislocation of lens
C0155373|ICD9CM|AB|379.34|Post dislocation of lens
C0155375|ICD9CM|PT|379.45|Argyll Robertson pupil, atypical
C0155375|ICD9CM|AB|379.45|Argyll robertson pupil
C0155376|ICD9CM|PT|379.49|Other anomalies of pupillary function
C0155376|ICD9CM|AB|379.49|Pupil funct anomaly NEC
C0155379|ICD9CM|PT|379.54|Nystagmus associated with disorders of the vestibular system
C0155379|ICD9CM|AB|379.54|Nystagms w vestibulr dis
C0155380|ICD9CM|AB|379.55|Dissociated nystagmus
C0155380|ICD9CM|PT|379.55|Dissociated nystagmus
C0155382|ICD9CM|PT|379.58|Deficiencies of smooth pursuit movements
C0155382|ICD9CM|AB|379.58|Smooth pursuit mvmnt def
C0155383|ICD9CM|PT|379.59|Other irregularities of eye movements
C0155383|ICD9CM|AB|379.59|Irregular eye mvmnts NEC
C0155384|ICD9CM|PT|379.8|Other specified disorders of eye and adnexa
C0155384|ICD9CM|AB|379.8|Eye disorders NEC
C0155386|ICD9CM|AB|379.92|Swelling or mass of eye
C0155386|ICD9CM|PT|379.92|Swelling or mass of eye
C0155387|ICD9CM|PT|379.99|Other ill-defined disorders of eye
C0155387|ICD9CM|AB|379.99|Ill-defined eye dis NEC
C0155388|ICD9CM|HT|380|Disorders of external ear
C0155388|ICD9CM|PT|380.9|Unspecified disorder of external ear
C0155388|ICD9CM|AB|380.9|Dis external ear NOS
C0155389|ICD9CM|AB|380.00|Perichondritis pinna NOS
C0155389|ICD9CM|PT|380.00|Perichondritis of pinna, unspecified
C0155389|ICD9CM|HT|380.0|Perichondritis and chondritis of pinna
C0155390|ICD9CM|PT|380.01|Acute perichondritis of pinna
C0155390|ICD9CM|AB|380.01|Ac perichondritis pinna
C0155391|ICD9CM|PT|380.02|Chronic perichondritis of pinna
C0155391|ICD9CM|AB|380.02|Chr perichondritis pinna
C0155392|ICD9CM|AB|380.11|Acute infection of pinna
C0155392|ICD9CM|PT|380.11|Acute infection of pinna
C0155394|ICD9CM|PT|380.13|Other acute infections of external ear
C0155394|ICD9CM|AB|380.13|Ac infect extern ear NEC
C0155395|ICD9CM|AB|380.14|Malignant otitis externa
C0155395|ICD9CM|PT|380.14|Malignant otitis externa
C0155396|ICD9CM|PT|380.15|Chronic mycotic otitis externa
C0155396|ICD9CM|AB|380.15|Chr mycot otitis externa
C0155397|ICD9CM|PT|380.16|Other chronic infective otitis externa
C0155397|ICD9CM|AB|380.16|Chr inf otit externa NEC
C0155398|ICD9CM|PT|380.21|Cholesteatoma of external ear
C0155398|ICD9CM|AB|380.21|Cholesteatoma extern ear
C0155399|ICD9CM|PT|380.22|Other acute otitis externa
C0155399|ICD9CM|AB|380.22|Acute otitis externa NEC
C0155400|ICD9CM|PT|380.23|Other chronic otitis externa
C0155400|ICD9CM|AB|380.23|Chr otitis externa NEC
C0155402|ICD9CM|AB|380.30|Disorder of pinna NOS
C0155402|ICD9CM|PT|380.30|Disorder of pinna, unspecified
C0155404|ICD9CM|PT|380.39|Other noninfectious disorders of pinna
C0155404|ICD9CM|AB|380.39|Noninfect dis pinna NEC
C0155405|ICD9CM|HT|380.5|Acquired stenosis of external ear canal
C0155405|ICD9CM|PT|380.50|Acquired stenosis of external ear canal, unspecified as to cause
C0155405|ICD9CM|AB|380.50|Acq stenos ear canal NOS
C0155410|ICD9CM|HT|380.8|Other disorders of external ear
C0155410|ICD9CM|PT|380.89|Other disorders of external ear
C0155410|ICD9CM|AB|380.89|Dis external ear NEC
C0155411|ICD9CM|PT|380.81|Exostosis of external ear canal
C0155411|ICD9CM|AB|380.81|Exostosis ext ear canal
C0155413|ICD9CM|HT|381|Nonsuppurative otitis media and Eustachian tube disorders
C0155415|ICD9CM|PT|381.01|Acute serous otitis media
C0155415|ICD9CM|AB|381.01|Ac serous otitis media
C0155418|ICD9CM|PT|381.04|Acute allergic serous otitis media
C0155418|ICD9CM|AB|381.04|Ac allergic serous OM
C0155419|ICD9CM|PT|381.05|Acute allergic mucoid otitis media
C0155419|ICD9CM|AB|381.05|Ac allergic mucoid OM
C0155420|ICD9CM|PT|381.06|Acute allergic sanguinous otitis media
C0155420|ICD9CM|AB|381.06|Ac allerg sanguinous OM
C0155421|ICD9CM|HT|381.1|Chronic serous otitis media
C0155422|ICD9CM|PT|381.10|Chronic serous otitis media, simple or unspecified
C0155422|ICD9CM|AB|381.10|Chr serous OM simp/NOS
C0155423|ICD9CM|PT|381.19|Other chronic serous otitis media
C0155423|ICD9CM|AB|381.19|Chr serous OM NEC
C0155426|ICD9CM|PT|381.29|Other chronic mucoid otitis media
C0155426|ICD9CM|AB|381.29|Chr mucoid OM NEC
C0155427|ICD9CM|PT|381.3|Other and unspecified chronic nonsuppurative otitis media
C0155427|ICD9CM|AB|381.3|Chr nonsup OM NOS/NEC
C0155428|ICD9CM|HT|381.5|Eustachian salpingitis
C0155428|ICD9CM|PT|381.50|Eustachian salpingitis, unspecified
C0155428|ICD9CM|AB|381.50|Eustachian salping NOS
C0155429|ICD9CM|PT|381.51|Acute Eustachian salpingitis
C0155429|ICD9CM|AB|381.51|Ac eustachian salping
C0155430|ICD9CM|PT|381.52|Chronic Eustachian salpingitis
C0155430|ICD9CM|AB|381.52|Chr eustachian salping
C0155431|ICD9CM|PT|381.61|Osseous obstruction of Eustachian tube
C0155431|ICD9CM|AB|381.61|Osseous eustachian obstr
C0155433|ICD9CM|PT|381.63|Extrinsic cartilagenous obstruction of Eustachian tube
C0155433|ICD9CM|AB|381.63|Extrinsic eustach obstr
C0155434|ICD9CM|AB|381.7|Patulous eustachian tube
C0155434|ICD9CM|PT|381.7|Patulous Eustachian tube
C0155435|ICD9CM|HT|381.8|Other disorders of Eustachian tube
C0155435|ICD9CM|PT|381.89|Other disorders of Eustachian tube
C0155435|ICD9CM|AB|381.89|Eustachian tube dis NEC
C0155439|ICD9CM|PT|382.02|Acute suppurative otitis media in diseases classified elsewhere
C0155439|ICD9CM|AB|382.02|Ac supp OM in oth dis
C0155440|ICD9CM|PT|382.1|Chronic tubotympanic suppurative otitis media
C0155440|ICD9CM|AB|382.1|Chr tubotympan suppur OM
C0155441|ICD9CM|PT|382.2|Chronic atticoantral suppurative otitis media
C0155441|ICD9CM|AB|382.2|Chr atticoantral sup OM
C0155442|ICD9CM|HT|383|Mastoiditis and related conditions
C0155445|ICD9CM|PT|383.01|Subperiosteal abscess of mastoid
C0155445|ICD9CM|AB|383.01|Subperi mastoid abscess
C0155446|ICD9CM|PT|383.02|Acute mastoiditis with other complications
C0155446|ICD9CM|AB|383.02|Ac mastoiditis-compl NEC
C0155447|ICD9CM|AB|383.1|Chronic mastoiditis
C0155447|ICD9CM|PT|383.1|Chronic mastoiditis
C0155448|ICD9CM|HT|383.2|Petrositis
C0155448|ICD9CM|AB|383.20|Petrositis NOS
C0155448|ICD9CM|PT|383.20|Petrositis, unspecified
C0155449|ICD9CM|AB|383.21|Acute petrositis
C0155449|ICD9CM|PT|383.21|Acute petrositis
C0155450|ICD9CM|AB|383.22|Chronic petrositis
C0155450|ICD9CM|PT|383.22|Chronic petrositis
C0155452|ICD9CM|HT|383.3|Complications following mastoidectomy
C0155452|ICD9CM|PT|383.30|Postmastoidectomy complication, unspecified
C0155452|ICD9CM|AB|383.30|Postmastoid compl NOS
C0155453|ICD9CM|PT|383.31|Mucosal cyst of postmastoidectomy cavity
C0155453|ICD9CM|AB|383.31|Postmastoid mucosal cyst
C0155454|ICD9CM|PT|383.32|Recurrent cholesteatoma of postmastoidectomy cavity
C0155454|ICD9CM|AB|383.32|Postmastoid cholesteatma
C0155455|ICD9CM|PT|383.33|Granulations of postmastoidectomy cavity
C0155455|ICD9CM|AB|383.33|Postmastoid granulations
C0155456|ICD9CM|HT|383.8|Other disorders of mastoid
C0155456|ICD9CM|PT|383.89|Other disorders of mastoid
C0155456|ICD9CM|AB|383.89|Disorders of mastoid NEC
C0155458|ICD9CM|HT|384|Other disorders of tympanic membrane
C0155459|ICD9CM|HT|384.0|Acute myringitis without mention of otitis media
C0155460|ICD9CM|AB|384.00|Acute myringitis NOS
C0155460|ICD9CM|PT|384.00|Acute myringitis, unspecified
C0155461|ICD9CM|AB|384.01|Bullous myringitis
C0155461|ICD9CM|PT|384.01|Bullous myringitis
C0155462|ICD9CM|PT|384.09|Other acute myringitis without mention of otitis media
C0155462|ICD9CM|AB|384.09|Acute myringitis NEC
C0155464|ICD9CM|PT|384.21|Central perforation of tympanic membrane
C0155464|ICD9CM|AB|384.21|Cent perf tympanic memb
C0155465|ICD9CM|PT|384.22|Attic perforation of tympanic membrane
C0155465|ICD9CM|AB|384.22|Attic perf tympanic memb
C0155466|ICD9CM|PT|384.23|Other marginal perforation of tympanic membrane
C0155466|ICD9CM|AB|384.23|Marginal perf tymp NEC
C0155467|ICD9CM|PT|384.24|Multiple perforations of tympanic membrane
C0155467|ICD9CM|AB|384.24|Mult perf tympanic memb
C0155468|ICD9CM|PT|384.25|Total perforation of tympanic membrane
C0155468|ICD9CM|AB|384.25|Total perf tympanic memb
C0155469|ICD9CM|HT|384.8|Other specified disorders of tympanic membrane
C0155470|ICD9CM|PT|384.81|Atrophic flaccid tympanic membrane
C0155470|ICD9CM|AB|384.81|Atrophic flaccid tympan
C0155471|ICD9CM|PT|384.82|Atrophic nonflaccid tympanic membrane
C0155471|ICD9CM|AB|384.82|Atrophic nonflaccid tymp
C0155472|ICD9CM|HT|385|Other disorders of middle ear and mastoid
C0155472|ICD9CM|HT|385.8|Other disorders of middle ear and mastoid
C0155472|ICD9CM|PT|385.89|Other disorders of middle ear and mastoid
C0155472|ICD9CM|AB|385.89|Dis mid ear/mastoid NEC
C0155477|ICD9CM|PT|385.09|Tympanosclerosis involving other combination of structures
C0155477|ICD9CM|AB|385.09|Tympnsclr-oth site comb
C0155478|ICD9CM|HT|385.1|Adhesive middle ear disease
C0155478|ICD9CM|PT|385.10|Adhesive middle ear disease, unspecified as to involvement
C0155478|ICD9CM|AB|385.10|Adhesive mid ear dis NOS
C0155480|ICD9CM|PT|385.11|Adhesions of drum head to incus
C0155480|ICD9CM|AB|385.11|Adhesion tympanum-incus
C0155481|ICD9CM|PT|385.12|Adhesions of drum head to stapes
C0155481|ICD9CM|AB|385.12|Adhesion tympanum-stapes
C0155482|ICD9CM|PT|385.13|Adhesions of drum head to promontorium
C0155482|ICD9CM|AB|385.13|Adhesion tymp-promontor
C0155483|ICD9CM|PT|385.19|Other middle ear adhesions and combinations
C0155483|ICD9CM|AB|385.19|Adhesive mid ear dis NEC
C0155484|ICD9CM|HT|385.2|Other acquired abnormality of ear ossicles
C0155486|ICD9CM|PT|385.22|Impaired mobility of other ear ossicles
C0155486|ICD9CM|AB|385.22|Ankylosis ear ossicl NEC
C0155487|ICD9CM|PT|385.23|Discontinuity or dislocation of ear ossicles
C0155487|ICD9CM|AB|385.23|Dislocation ear ossicle
C0155488|ICD9CM|PT|385.24|Partial loss or necrosis of ear ossicles
C0155488|ICD9CM|AB|385.24|Partial loss ear ossicle
C0155489|ICD9CM|AB|385.31|Cholesteatoma of attic
C0155489|ICD9CM|PT|385.31|Cholesteatoma of attic
C0155490|ICD9CM|AB|385.32|Cholesteatoma middle ear
C0155490|ICD9CM|PT|385.32|Cholesteatoma of middle ear
C0155491|ICD9CM|PT|385.35|Diffuse cholesteatosis of middle ear and mastoid
C0155491|ICD9CM|AB|385.35|Diffuse cholesteatosis
C0155493|ICD9CM|PT|385.83|Retained foreign body of middle ear
C0155493|ICD9CM|AB|385.83|Foreign body middle ear
C0155494|ICD9CM|PT|385.9|Unspecified disorder of middle ear and mastoid
C0155494|ICD9CM|AB|385.9|Dis mid ear/mastoid NOS
C0155496|ICD9CM|PT|386.01|Active Ménière's disease, cochleovestibular
C0155496|ICD9CM|AB|386.01|Actv Meniere,cochlvestib
C0155497|ICD9CM|PT|386.02|Active Ménière's disease, cochlear
C0155497|ICD9CM|AB|386.02|Active Meniere, cochlear
C0155498|ICD9CM|PT|386.03|Active Ménière's disease, vestibular
C0155498|ICD9CM|AB|386.03|Actv Meniere, vestibular
C0155499|ICD9CM|PT|386.04|Inactive Ménière's disease
C0155499|ICD9CM|AB|386.04|Inactive Meniere's dis
C0155501|ICD9CM|AB|386.10|Peripheral vertigo NOS
C0155501|ICD9CM|PT|386.10|Peripheral vertigo, unspecified
C0155502|ICD9CM|PT|386.11|Benign paroxysmal positional vertigo
C0155502|ICD9CM|AB|386.11|Benign parxysmal vertigo
C0155503|ICD9CM|AB|386.2|Central origin vertigo
C0155503|ICD9CM|PT|386.2|Vertigo of central origin
C0155504|ICD9CM|AB|386.31|Serous labyrinthitis
C0155504|ICD9CM|PT|386.31|Serous labyrinthitis
C0155505|ICD9CM|PT|386.32|Circumscribed labyrinthitis
C0155505|ICD9CM|AB|386.32|Circumscri labyrinthitis
C0155506|ICD9CM|PT|386.33|Suppurative labyrinthitis
C0155506|ICD9CM|AB|386.33|Suppurativ labyrinthitis
C0155507|ICD9CM|AB|386.34|Toxic labyrinthitis
C0155507|ICD9CM|PT|386.34|Toxic labyrinthitis
C0155508|ICD9CM|AB|386.35|Viral labyrinthitis
C0155508|ICD9CM|PT|386.35|Viral labyrinthitis
C0155509|ICD9CM|HT|386.4|Labyrinthine fistula
C0155509|ICD9CM|AB|386.40|Labyrinthine fistula NOS
C0155509|ICD9CM|PT|386.40|Labyrinthine fistula, unspecified
C0155512|ICD9CM|PT|386.43|Semicircular canal fistula
C0155512|ICD9CM|AB|386.43|Semicircul canal fistula
C0155513|ICD9CM|PT|386.48|Labyrinthine fistula of combined sites
C0155513|ICD9CM|AB|386.48|Labyrinth fistula comb
C0155514|ICD9CM|HT|386.5|Labyrinthine dysfunction
C0155514|ICD9CM|PT|386.50|Labyrinthine dysfunction, unspecified
C0155514|ICD9CM|AB|386.50|Labyrinthine dysfunc NOS
C0155515|ICD9CM|PT|386.51|Hyperactive labyrinth, unilateral
C0155515|ICD9CM|AB|386.51|Hypract labyrinth unilat
C0155516|ICD9CM|PT|386.52|Hyperactive labyrinth, bilateral
C0155516|ICD9CM|AB|386.52|Hyperact labyrinth bilat
C0155517|ICD9CM|PT|386.53|Hypoactive labyrinth, unilateral
C0155517|ICD9CM|AB|386.53|Hypoact labyrinth unilat
C0155518|ICD9CM|PT|386.54|Hypoactive labyrinth, bilateral
C0155518|ICD9CM|AB|386.54|Hypoact labyrinth bilat
C0155519|ICD9CM|PT|386.55|Loss of labyrinthine reactivity, unilateral
C0155519|ICD9CM|AB|386.55|Loss labyrn react unilat
C0155520|ICD9CM|PT|386.56|Loss of labyrinthine reactivity, bilateral
C0155520|ICD9CM|AB|386.56|Loss labyrin react bilat
C0155521|ICD9CM|PT|386.58|Other forms and combinations of labyrinthine dysfunction
C0155521|ICD9CM|AB|386.58|Labyrinthine dysfunc NEC
C0155522|ICD9CM|PT|386.8|Other disorders of labyrinth
C0155522|ICD9CM|AB|386.8|Disorders labyrinth NEC
C0155523|ICD9CM|PT|386.9|Unspecified vertiginous syndromes and labyrinthine disorders
C0155523|ICD9CM|HT|386|Vertiginous syndromes and other disorders of vestibular system
C0155523|ICD9CM|AB|386.9|Vertiginous synd NOS
C0155524|ICD9CM|PT|387.0|Otosclerosis involving oval window, nonobliterative
C0155524|ICD9CM|AB|387.0|Otoscler-oval wnd nonobl
C0155525|ICD9CM|PT|387.1|Otosclerosis involving oval window, obliterative
C0155525|ICD9CM|AB|387.1|Otoscler-oval wndw oblit
C0155526|ICD9CM|AB|387.2|Cochlear otosclerosis
C0155526|ICD9CM|PT|387.2|Cochlear otosclerosis
C0155527|ICD9CM|HT|388|Other disorders of ear
C0155527|ICD9CM|PT|388.8|Other disorders of ear
C0155527|ICD9CM|AB|388.8|Disorders of ear NEC
C0155528|ICD9CM|HT|388.0|Degenerative and vascular disorders of ear
C0155528|ICD9CM|PT|388.00|Degenerative and vascular disorders, unspecified
C0155528|ICD9CM|AB|388.00|Degen/vascul dis ear NOS
C0155530|ICD9CM|PT|388.02|Transient ischemic deafness
C0155530|ICD9CM|AB|388.02|Trans ischemic deafness
C0155531|ICD9CM|HT|388.1|Noise effects on inner ear
C0155531|ICD9CM|PT|388.10|Noise effects on inner ear, unspecified
C0155531|ICD9CM|AB|388.10|Noise effect-ear/NOS
C0155532|ICD9CM|PT|388.11|Acoustic trauma (explosive) to ear
C0155532|ICD9CM|AB|388.11|Acoustic trauma
C0155533|ICD9CM|AB|388.31|Subjective tinnitus
C0155533|ICD9CM|PT|388.31|Subjective tinnitus
C0155534|ICD9CM|AB|388.32|Objective tinnitus
C0155534|ICD9CM|PT|388.32|Objective tinnitus
C0155535|ICD9CM|HT|388.4|Other abnormal auditory perception
C0155537|ICD9CM|PT|388.43|Impairment of auditory discrimination
C0155537|ICD9CM|AB|388.43|Impairm auditory discrim
C0155540|ICD9CM|HT|388.6|Otorrhea
C0155540|ICD9CM|AB|388.60|Otorrhea NOS
C0155540|ICD9CM|PT|388.60|Otorrhea, unspecified
C0155541|ICD9CM|PT|388.69|Other otorrhea
C0155541|ICD9CM|AB|388.69|Otorrhea NEC
C0155542|ICD9CM|AB|388.71|Otogenic pain
C0155542|ICD9CM|PT|388.71|Otogenic pain
C0155544|ICD9CM|PT|389.01|Conductive hearing loss, external ear
C0155544|ICD9CM|AB|389.01|Conduc hear loss ext ear
C0155545|ICD9CM|PT|389.02|Conductive hearing loss, tympanic membrane
C0155545|ICD9CM|AB|389.02|Conduct hear loss tympan
C0155546|ICD9CM|PT|389.03|Conductive hearing loss, middle ear
C0155546|ICD9CM|AB|389.03|Conduc hear loss mid ear
C0155547|ICD9CM|PT|389.04|Conductive hearing loss, inner ear
C0155547|ICD9CM|AB|389.04|Cond hear loss inner ear
C0155548|ICD9CM|PT|389.08|Conductive hearing loss of combined types
C0155548|ICD9CM|AB|389.08|Cond hear loss comb type
C0155552|ICD9CM|HT|389.2|Mixed conductive and sensorineural hearing loss
C0155552|ICD9CM|AB|389.20|Mixed hearing loss NOS
C0155552|ICD9CM|PT|389.20|Mixed hearing loss, unspecified
C0155555|ICD9CM|PT|391.0|Acute rheumatic pericarditis
C0155555|ICD9CM|AB|391.0|Acute rheumatic pericard
C0155556|ICD9CM|PT|391.1|Acute rheumatic endocarditis
C0155556|ICD9CM|AB|391.1|Acute rheumatic endocard
C0155557|ICD9CM|PT|391.2|Acute rheumatic myocarditis
C0155557|ICD9CM|AB|391.2|Ac rheumatic myocarditis
C0155558|ICD9CM|PT|391.8|Other acute rheumatic heart disease
C0155558|ICD9CM|AB|391.8|Ac rheumat hrt dis NEC
C0155559|ICD9CM|PT|392.0|Rheumatic chorea with heart involvement
C0155559|ICD9CM|AB|392.0|Rheum chorea w hrt invol
C0155561|ICD9CM|PT|393|Chronic rheumatic pericarditis
C0155561|ICD9CM|AB|393|Chr rheumatic pericard
C0155563|ICD9CM|PT|394.1|Rheumatic mitral insufficiency
C0155563|ICD9CM|AB|394.1|Rheumatic mitral insuff
C0155567|ICD9CM|PT|395.0|Rheumatic aortic stenosis
C0155567|ICD9CM|AB|395.0|Rheumat aortic stenosis
C0155568|ICD9CM|PT|395.1|Rheumatic aortic insufficiency
C0155568|ICD9CM|AB|395.1|Rheumatic aortic insuff
C0155569|ICD9CM|PT|395.2|Rheumatic aortic stenosis with insufficiency
C0155569|ICD9CM|AB|395.2|Rheum aortic sten/insuff
C0155570|ICD9CM|PT|395.9|Other and unspecified rheumatic aortic diseases
C0155570|ICD9CM|AB|395.9|Rheum aortic dis NEC/NOS
C0155572|ICD9CM|PT|396.0|Mitral valve stenosis and aortic valve stenosis
C0155572|ICD9CM|AB|396.0|Mitral/aortic stenosis
C0155576|ICD9CM|PT|396.8|Multiple involvement of mitral and aortic valves
C0155576|ICD9CM|AB|396.8|Mitr/aortic mult involv
C0155578|ICD9CM|HT|397|Diseases of other endocardial structures
C0155579|ICD9CM|PT|397.1|Rheumatic diseases of pulmonary valve
C0155579|ICD9CM|AB|397.1|Rheum pulmon valve dis
C0155582|ICD9CM|PT|398.91|Rheumatic heart failure (congestive)
C0155582|ICD9CM|AB|398.91|Rheumatic heart failure
C0155583|ICD9CM|PT|401.1|Benign essential hypertension
C0155583|ICD9CM|AB|401.1|Benign hypertension
C0155584|ICD9CM|HT|402.0|Malignant hypertensive heart disease
C0155587|ICD9CM|HT|402.1|Benign hypertensive heart disease
C0155596|ICD9CM|HT|403.1|Hypertensive renal disease, benign
C0155596|ICD9CM|PT|403.10|Hypertensive chronic kidney disease, benign, with chronic kidney disease stage I through stage IV, or unspecified
C0155596|ICD9CM|AB|403.10|Ben hy kid w cr kid I-IV
C0155598|ICD9CM|PT|403.11|Hypertensive chronic kidney disease, benign, with chronic kidney disease stage V or end stage renal disease
C0155598|ICD9CM|AB|403.11|Ben hyp kid w cr kid V
C0155601|ICD9CM|HT|404.9|Hypertensive heart and renal disease, unspecified
C0155607|ICD9CM|HT|404.1|Hypertensive heart and renal disease, benign
C0155608|ICD9CM|PT|404.10|Hypertensive heart and chronic kidney disease, benign, without heart failure and with chronic kidney disease stage I through stage IV, or unspecified
C0155608|ICD9CM|AB|404.10|Ben hy ht/kd I-IV w/o hf
C0155609|ICD9CM|PT|404.11|Hypertensive heart and chronic kidney disease, benign, with heart failure and with chronic kidney disease stage I through stage IV, or unspecified
C0155609|ICD9CM|AB|404.11|Ben hyp ht/kd I-IV w hf
C0155610|ICD9CM|PT|404.12|Hypertensive heart and chronic kidney disease, benign, without heart failure and with chronic kidney disease stage V or end stage renal disease
C0155610|ICD9CM|AB|404.12|Ben hy ht/kd st V w/o hf
C0155611|ICD9CM|PT|404.13|Hypertensive heart and chronic kidney disease, benign, with heart failure and chronic kidney disease stage V or end stage renal disease
C0155611|ICD9CM|AB|404.13|Ben hyp ht/kd stg V w hf
C0155612|ICD9CM|PT|404.90|Hypertensive heart and chronic kidney disease, unspecified, without heart failure and with chronic kidney disease stage I through stage IV, or unspecified
C0155612|ICD9CM|AB|404.90|Hy ht/kd NOS I-IV w/o hf
C0155616|ICD9CM|HT|405|Secondary hypertension
C0155616|ICD9CM|HT|405.9|Unspecified secondary hypertension
C0155617|ICD9CM|HT|405.0|Malignant secondary hypertension
C0155619|ICD9CM|PT|405.09|Other malignant secondary hypertension
C0155619|ICD9CM|AB|405.09|Mal second hyperten NEC
C0155620|ICD9CM|HT|405.1|Benign secondary hypertension
C0155621|ICD9CM|PT|405.11|Benign renovascular hypertension
C0155621|ICD9CM|AB|405.11|Benign renovasc hyperten
C0155622|ICD9CM|PT|405.19|Other benign secondary hypertension
C0155622|ICD9CM|AB|405.19|Benign second hypert NEC
C0155624|ICD9CM|PT|405.91|Unspecified renovascular hypertension
C0155624|ICD9CM|AB|405.91|Renovasc hypertension
C0155626|ICD9CM|HT|410|Acute myocardial infarction
C0155626|ICD9CM|PT|410.90|Acute myocardial infarction of unspecified site, episode of care unspecified
C0155626|ICD9CM|HT|410.9|Acute myocardial infarction, unspecified site
C0155626|ICD9CM|AB|410.90|AMI NOS, unspecified
C0155627|ICD9CM|HT|410.0|Acute myocardial infarction, of anterolateral wall
C0155628|ICD9CM|PT|410.00|Acute myocardial infarction of anterolateral wall, episode of care unspecified
C0155628|ICD9CM|AB|410.00|AMI anterolateral,unspec
C0155629|ICD9CM|PT|410.01|Acute myocardial infarction of anterolateral wall, initial episode of care
C0155629|ICD9CM|AB|410.01|AMI anterolateral, init
C0155630|ICD9CM|PT|410.02|Acute myocardial infarction of anterolateral wall, subsequent episode of care
C0155630|ICD9CM|AB|410.02|AMI anterolateral,subseq
C0155631|ICD9CM|HT|410.1|Acute myocardial infarction, of other anterior wall
C0155632|ICD9CM|PT|410.10|Acute myocardial infarction of other anterior wall, episode of care unspecified
C0155632|ICD9CM|AB|410.10|AMI anterior wall,unspec
C0155633|ICD9CM|PT|410.11|Acute myocardial infarction of other anterior wall, initial episode of care
C0155633|ICD9CM|AB|410.11|AMI anterior wall, init
C0155634|ICD9CM|PT|410.12|Acute myocardial infarction of other anterior wall, subsequent episode of care
C0155634|ICD9CM|AB|410.12|AMI anterior wall,subseq
C0155636|ICD9CM|PT|410.20|Acute myocardial infarction of inferolateral wall, episode of care unspecified
C0155636|ICD9CM|AB|410.20|AMI inferolateral,unspec
C0155637|ICD9CM|PT|410.21|Acute myocardial infarction of inferolateral wall, initial episode of care
C0155637|ICD9CM|AB|410.21|AMI inferolateral, init
C0155638|ICD9CM|PT|410.22|Acute myocardial infarction of inferolateral wall, subsequent episode of care
C0155638|ICD9CM|AB|410.22|AMI inferolateral,subseq
C0155640|ICD9CM|PT|410.30|Acute myocardial infarction of inferoposterior wall, episode of care unspecified
C0155640|ICD9CM|AB|410.30|AMI inferopost, unspec
C0155641|ICD9CM|PT|410.31|Acute myocardial infarction of inferoposterior wall, initial episode of care
C0155641|ICD9CM|AB|410.31|AMI inferopost, initial
C0155642|ICD9CM|PT|410.32|Acute myocardial infarction of inferoposterior wall, subsequent episode of care
C0155642|ICD9CM|AB|410.32|AMI inferopost, subseq
C0155643|ICD9CM|HT|410.4|Acute myocardial infarction, of other inferior wall
C0155644|ICD9CM|PT|410.40|Acute myocardial infarction of other inferior wall, episode of care unspecified
C0155644|ICD9CM|AB|410.40|AMI inferior wall,unspec
C0155645|ICD9CM|PT|410.41|Acute myocardial infarction of other inferior wall, initial episode of care
C0155645|ICD9CM|AB|410.41|AMI inferior wall, init
C0155646|ICD9CM|PT|410.42|Acute myocardial infarction of other inferior wall, subsequent episode of care
C0155646|ICD9CM|AB|410.42|AMI inferior wall,subseq
C0155647|ICD9CM|HT|410.5|Acute myocardial infarction, of other lateral wall
C0155648|ICD9CM|PT|410.50|Acute myocardial infarction of other lateral wall, episode of care unspecified
C0155648|ICD9CM|AB|410.50|AMI lateral NEC, unspec
C0155649|ICD9CM|PT|410.51|Acute myocardial infarction of other lateral wall, initial episode of care
C0155649|ICD9CM|AB|410.51|AMI lateral NEC, initial
C0155650|ICD9CM|PT|410.52|Acute myocardial infarction of other lateral wall, subsequent episode of care
C0155650|ICD9CM|AB|410.52|AMI lateral NEC, subseq
C0155652|ICD9CM|PT|410.60|True posterior wall infarction, episode of care unspecified
C0155652|ICD9CM|AB|410.60|True post infarct,unspec
C0155653|ICD9CM|PT|410.61|True posterior wall infarction, initial episode of care
C0155653|ICD9CM|AB|410.61|True post infarct, init
C0155654|ICD9CM|PT|410.62|True posterior wall infarction, subsequent episode of care
C0155654|ICD9CM|AB|410.62|True post infarct,subseq
C0155655|ICD9CM|HT|410.7|Acute myocardial infarction, subendocardial infarction
C0155657|ICD9CM|PT|410.71|Subendocardial infarction, initial episode of care
C0155657|ICD9CM|AB|410.71|Subendo infarct, initial
C0155658|ICD9CM|PT|410.72|Subendocardial infarction, subsequent episode of care
C0155658|ICD9CM|AB|410.72|Subendo infarct, subseq
C0155659|ICD9CM|HT|410.8|Acute myocardial infarction, of other specified sites
C0155660|ICD9CM|PT|410.80|Acute myocardial infarction of other specified sites, episode of care unspecified
C0155660|ICD9CM|AB|410.80|AMI NEC, unspecified
C0155661|ICD9CM|PT|410.81|Acute myocardial infarction of other specified sites, initial episode of care
C0155661|ICD9CM|AB|410.81|AMI NEC, initial
C0155662|ICD9CM|PT|410.82|Acute myocardial infarction of other specified sites, subsequent episode of care
C0155662|ICD9CM|AB|410.82|AMI NEC, subsequent
C0155664|ICD9CM|PT|410.91|Acute myocardial infarction of unspecified site, initial episode of care
C0155664|ICD9CM|AB|410.91|AMI NOS, initial
C0155665|ICD9CM|PT|410.92|Acute myocardial infarction of unspecified site, subsequent episode of care
C0155665|ICD9CM|AB|410.92|AMI NOS, subsequent
C0155668|ICD9CM|PT|412|Old myocardial infarction
C0155668|ICD9CM|AB|412|Old myocardial infarct
C0155669|ICD9CM|HT|414|Other forms of chronic ischemic heart disease
C0155670|ICD9CM|PT|414.8|Other specified forms of chronic ischemic heart disease
C0155670|ICD9CM|AB|414.8|Chr ischemic hrt dis NEC
C0155671|ICD9CM|HT|415|Acute pulmonary heart disease
C0155672|ICD9CM|AB|415.0|Acute cor pulmonale
C0155672|ICD9CM|PT|415.0|Acute cor pulmonale
C0155673|ICD9CM|PT|416.8|Other chronic pulmonary heart diseases
C0155673|ICD9CM|AB|416.8|Chr pulmon heart dis NEC
C0155674|ICD9CM|HT|417|Other diseases of pulmonary circulation
C0155675|ICD9CM|PT|417.0|Arteriovenous fistula of pulmonary vessels
C0155675|ICD9CM|AB|417.0|Arterioven fistu pul ves
C0155676|ICD9CM|PT|417.1|Aneurysm of pulmonary artery
C0155676|ICD9CM|AB|417.1|Pulmon artery aneurysm
C0155677|ICD9CM|PT|417.8|Other specified diseases of pulmonary circulation
C0155677|ICD9CM|AB|417.8|Pulmon circulat dis NEC
C0155679|ICD9CM|HT|420|Acute pericarditis
C0155679|ICD9CM|AB|420.90|Acute pericarditis NOS
C0155679|ICD9CM|PT|420.90|Acute pericarditis, unspecified
C0155680|ICD9CM|HT|420.9|Other and unspecified acute pericarditis
C0155681|ICD9CM|PT|420.91|Acute idiopathic pericarditis
C0155681|ICD9CM|AB|420.91|Ac idiopath pericarditis
C0155683|ICD9CM|HT|421|Acute and subacute endocarditis
C0155686|ICD9CM|HT|422|Acute myocarditis
C0155686|ICD9CM|AB|422.90|Acute myocarditis NOS
C0155686|ICD9CM|PT|422.90|Acute myocarditis, unspecified
C0155687|ICD9CM|PT|422.0|Acute myocarditis in diseases classified elsewhere
C0155687|ICD9CM|AB|422.0|Ac myocardit in oth dis
C0155689|ICD9CM|AB|422.91|Idiopathic myocarditis
C0155689|ICD9CM|PT|422.91|Idiopathic myocarditis
C0155690|ICD9CM|AB|422.92|Septic myocarditis
C0155690|ICD9CM|PT|422.92|Septic myocarditis
C0155691|ICD9CM|AB|422.93|Toxic myocarditis
C0155691|ICD9CM|PT|422.93|Toxic myocarditis
C0155692|ICD9CM|PT|422.99|Other acute myocarditis
C0155692|ICD9CM|HT|422.9|Other and unspecified acute myocarditis
C0155692|ICD9CM|AB|422.99|Acute myocarditis NEC
C0155694|ICD9CM|PT|423.8|Other specified diseases of pericardium
C0155694|ICD9CM|AB|423.8|Pericardial disease NEC
C0155695|ICD9CM|HT|424|Other diseases of endocardium
C0155699|ICD9CM|PT|425.8|Cardiomyopathy in other diseases classified elsewhere
C0155699|ICD9CM|AB|425.8|Cardiomyopath in oth dis
C0155700|ICD9CM|PT|426.12|Mobitz (type) II atrioventricular block
C0155700|ICD9CM|AB|426.12|Atrioven block-mobitz ii
C0155702|ICD9CM|PT|426.2|Left bundle branch hemiblock
C0155702|ICD9CM|AB|426.2|Left bb hemiblock
C0155703|ICD9CM|PT|426.3|Other left bundle branch block
C0155703|ICD9CM|AB|426.3|Left bb block NEC
C0155704|ICD9CM|PT|426.51|Right bundle branch block and left posterior fascicular block
C0155704|ICD9CM|AB|426.51|Rt bbb/lft post fasc blk
C0155705|ICD9CM|PT|426.52|Right bundle branch block and left anterior fascicular block
C0155705|ICD9CM|AB|426.52|Rt bbb/lft ant fasc blk
C0155706|ICD9CM|PT|426.53|Other bilateral bundle branch block
C0155706|ICD9CM|AB|426.53|Bilat bb block NEC
C0155707|ICD9CM|AB|426.54|Trifascicular block
C0155707|ICD9CM|PT|426.54|Trifascicular block
C0155708|ICD9CM|HT|426.8|Other specified conduction disorders
C0155708|ICD9CM|PT|426.89|Other specified conduction disorders
C0155708|ICD9CM|AB|426.89|Conduction disorder NEC
C0155709|ICD9CM|HT|427.3|Atrial fibrillation and flutter
C0155710|ICD9CM|HT|427.4|Ventricular fibrillation and flutter
C0155711|ICD9CM|HT|429|Ill-defined descriptions and complications of heart disease
C0155712|ICD9CM|PT|429.5|Rupture of chordae tendineae
C0155712|ICD9CM|AB|429.5|Chordae tendinae rupture
C0155713|ICD9CM|PT|429.6|Rupture of papillary muscle
C0155713|ICD9CM|AB|429.6|Papillary muscle rupture
C0155717|ICD9CM|HT|429.8|Other ill-defined heart diseases
C0155717|ICD9CM|PT|429.89|Other ill-defined heart diseases
C0155717|ICD9CM|AB|429.89|Ill-defined hrt dis NEC
C0155718|ICD9CM|PT|429.81|Other disorders of papillary muscle
C0155718|ICD9CM|AB|429.81|Papillary muscle dis NEC
C0155719|ICD9CM|HT|432|Other and unspecified intracranial hemorrhage
C0155724|ICD9CM|HT|433.2|Occlusion and stenosis of vertebral artery
C0155725|ICD9CM|HT|433.3|Occlusion and stenosis of multiple and bilateral precerebral arteries
C0155726|ICD9CM|HT|433.8|Occlusion and stenosis of other specified precerebral artery
C0155727|ICD9CM|HT|433.9|Occlusion and stenosis of unspecified precerebral artery
C0155727|ICD9CM|HT|433|Occlusion and stenosis of precerebral arteries
C0155728|ICD9CM|PT|435.8|Other specified transient cerebral ischemias
C0155728|ICD9CM|AB|435.8|Trans cereb ischemia NEC
C0155729|ICD9CM|PT|437.8|Other ill-defined cerebrovascular disease
C0155729|ICD9CM|HT|437|Other and ill-defined cerebrovascular disease
C0155729|ICD9CM|AB|437.8|Cerebrovasc disease NEC
C0155730|ICD9CM|PT|437.3|Cerebral aneurysm, nonruptured
C0155730|ICD9CM|AB|437.3|Nonrupt cerebral aneurym
C0155731|ICD9CM|PT|437.6|Nonpyogenic thrombosis of intracranial venous sinus
C0155731|ICD9CM|AB|437.6|Nonpyogen thrombos sinus
C0155732|ICD9CM|HT|438|Late effects of cerebrovascular disease
C0155732|ICD9CM|PT|438.9|Unspecified late effects of cerebrovascular disease
C0155732|ICD9CM|AB|438.9|Late effect CV dis NOS
C0155733|ICD9CM|PT|440.0|Atherosclerosis of aorta
C0155733|ICD9CM|AB|440.0|Aortic atherosclerosis
C0155734|ICD9CM|PT|440.1|Atherosclerosis of renal artery
C0155734|ICD9CM|AB|440.1|Renal artery atheroscler
C0155740|ICD9CM|HT|442|Other aneurysm
C0155741|ICD9CM|PT|442.0|Aneurysm of artery of upper extremity
C0155741|ICD9CM|AB|442.0|Upper extremity aneurysm
C0155742|ICD9CM|PT|442.1|Aneurysm of renal artery
C0155742|ICD9CM|AB|442.1|Renal artery aneurysm
C0155744|ICD9CM|PT|442.3|Aneurysm of artery of lower extremity
C0155744|ICD9CM|AB|442.3|Lower extremity aneurysm
C0155745|ICD9CM|PT|442.81|Aneurysm of artery of neck
C0155745|ICD9CM|AB|442.81|Aneurysm of neck
C0155746|ICD9CM|PT|442.82|Aneurysm of subclavian artery
C0155746|ICD9CM|AB|442.82|Subclavian aneurysm
C0155747|ICD9CM|PT|442.83|Aneurysm of splenic artery
C0155747|ICD9CM|AB|442.83|Splenic artery aneurysm
C0155748|ICD9CM|PT|442.84|Aneurysm of other visceral artery
C0155748|ICD9CM|AB|442.84|Visceral aneurysm NEC
C0155749|ICD9CM|HT|444|Arterial embolism and thrombosis
C0155750|ICD9CM|PT|444.1|Embolism and thrombosis of thoracic aorta
C0155750|ICD9CM|AB|444.1|Thoracic aortic embolism
C0155754|ICD9CM|HT|444.8|Embolism and thrombosis of other specified artery
C0155755|ICD9CM|PT|444.81|Embolism and thrombosis of iliac artery
C0155755|ICD9CM|AB|444.81|Iliac artery embolism
C0155757|ICD9CM|HT|446|Polyarteritis nodosa and allied conditions
C0155758|ICD9CM|PT|446.29|Other specified hypersensitivity angiitis
C0155758|ICD9CM|AB|446.29|Hypersensit angiitis NEC
C0155759|ICD9CM|HT|447|Other disorders of arteries and arterioles
C0155760|ICD9CM|AB|447.2|Rupture of artery
C0155760|ICD9CM|PT|447.2|Rupture of artery
C0155761|ICD9CM|AB|447.3|Renal artery hyperplasia
C0155761|ICD9CM|PT|447.3|Hyperplasia of renal artery
C0155762|ICD9CM|AB|447.5|Necrosis of artery
C0155762|ICD9CM|PT|447.5|Necrosis of artery
C0155763|ICD9CM|PT|447.8|Other specified disorders of arteries and arterioles
C0155763|ICD9CM|AB|447.8|Arterial disease NEC
C0155764|ICD9CM|PT|447.9|Unspecified disorders of arteries and arterioles
C0155764|ICD9CM|AB|447.9|Arterial disease NOS
C0155765|ICD9CM|HT|448|Disease of capillaries
C0155770|ICD9CM|PT|451.19|Phlebitis and thrombophlebitis of deep veins of lower extremities, other
C0155770|ICD9CM|AB|451.19|Deep phlebitis-leg NEC
C0155772|ICD9CM|PT|451.81|Phlebitis and thrombophlebitis of iliac vein
C0155772|ICD9CM|AB|451.81|Iliac thrombophlebitis
C0155773|ICD9CM|AB|452|Portal vein thrombosis
C0155773|ICD9CM|PT|452|Portal vein thrombosis
C0155774|ICD9CM|HT|453|Other venous embolism and thrombosis
C0155776|ICD9CM|AB|453.3|Renal vein thrombosis
C0155776|ICD9CM|PT|453.3|Other venous embolism and thrombosis of renal vein
C0155778|ICD9CM|HT|454|Varicose veins of lower extremities
C0155779|ICD9CM|PT|454.2|Varicose veins of lower extremities with ulcer and inflammation
C0155779|ICD9CM|AB|454.2|Varicos leg ulcer/inflam
C0155781|ICD9CM|PT|455.1|Internal thrombosed hemorrhoids
C0155781|ICD9CM|AB|455.1|Int thrombos hemorrhoid
C0155782|ICD9CM|PT|455.2|Internal hemorrhoids with other complication
C0155782|ICD9CM|AB|455.2|Int hemrrhoid w comp NEC
C0155784|ICD9CM|PT|455.4|External thrombosed hemorrhoids
C0155784|ICD9CM|AB|455.4|Ext thrombos hemorrhoid
C0155785|ICD9CM|PT|455.5|External hemorrhoids with other complication
C0155785|ICD9CM|AB|455.5|Ext hemrrhoid w comp NEC
C0155787|ICD9CM|PT|455.8|Unspecified hemorrhoids with other complication
C0155787|ICD9CM|AB|455.8|Hemrrhoid NOS w comp NEC
C0155788|ICD9CM|PT|455.9|Residual hemorrhoidal skin tags
C0155788|ICD9CM|AB|455.9|Residual hemorrhoid tags
C0155789|ICD9CM|PT|456.0|Esophageal varices with bleeding
C0155789|ICD9CM|AB|456.0|Esophag varices w bleed
C0155791|ICD9CM|HT|456.2|Esophageal varices in diseases classified elsewhere
C0155792|ICD9CM|PT|456.20|Esophageal varices in diseases classified elsewhere, with bleeding
C0155792|ICD9CM|AB|456.20|Bleed esoph var oth dis
C0155793|ICD9CM|PT|456.21|Esophageal varices in diseases classified elsewhere, without mention of bleeding
C0155793|ICD9CM|AB|456.21|Esoph varice oth dis NOS
C0155794|ICD9CM|AB|456.3|Sublingual varices
C0155794|ICD9CM|PT|456.3|Sublingual varices
C0155795|ICD9CM|AB|456.5|Pelvic varices
C0155795|ICD9CM|PT|456.5|Pelvic varices
C0155796|ICD9CM|AB|456.6|Vulval varices
C0155796|ICD9CM|PT|456.6|Vulval varices
C0155797|ICD9CM|AB|456.8|Varices of other sites
C0155797|ICD9CM|PT|456.8|Varices of other sites
C0155797|ICD9CM|HT|456|Varicose veins of other sites
C0155799|ICD9CM|HT|457|Noninfectious disorders of lymphatic channels
C0155799|ICD9CM|PT|457.9|Unspecified noninfectious disorder of lymphatic channels
C0155799|ICD9CM|AB|457.9|Noninfect lymph dis NOS
C0155800|ICD9CM|AB|458.1|Chronic hypotension
C0155800|ICD9CM|PT|458.1|Chronic hypotension
C0155802|ICD9CM|AB|459.2|Compression of vein
C0155802|ICD9CM|PT|459.2|Compression of vein
C0155803|ICD9CM|HT|459.8|Other specified disorders of circulatory system
C0155803|ICD9CM|PT|459.89|Other specified disorders of circulatory system
C0155803|ICD9CM|AB|459.89|Circulatory disease NEC
C0155804|ICD9CM|PT|461.0|Acute maxillary sinusitis
C0155804|ICD9CM|AB|461.0|Ac maxillary sinusitis
C0155805|ICD9CM|PT|461.1|Acute frontal sinusitis
C0155805|ICD9CM|AB|461.1|Ac frontal sinusitis
C0155806|ICD9CM|PT|461.2|Acute ethmoidal sinusitis
C0155806|ICD9CM|AB|461.2|Ac ethmoidal sinusitis
C0155807|ICD9CM|PT|461.3|Acute sphenoidal sinusitis
C0155807|ICD9CM|AB|461.3|Ac sphenoidal sinusitis
C0155808|ICD9CM|AB|461.8|Other acute sinusitis
C0155808|ICD9CM|PT|461.8|Other acute sinusitis
C0155810|ICD9CM|PT|464.11|Acute tracheitis with obstruction
C0155810|ICD9CM|AB|464.11|Ac tracheitis w obstruct
C0155811|ICD9CM|HT|464|Acute laryngitis and tracheitis
C0155811|ICD9CM|HT|464.2|Acute laryngotracheitis
C0155813|ICD9CM|PT|464.21|Acute laryngotracheitis with obstruction
C0155813|ICD9CM|AB|464.21|Ac laryngotrach w obstr
C0155814|ICD9CM|HT|464.3|Acute epiglottitis
C0155815|ICD9CM|PT|464.31|Acute epiglottitis with obstruction
C0155815|ICD9CM|AB|464.31|Ac epiglottitis w obstr
C0155816|ICD9CM|HT|465|Acute upper respiratory infections of multiple or unspecified sites
C0155817|ICD9CM|AB|465.0|Acute laryngopharyngitis
C0155817|ICD9CM|PT|465.0|Acute laryngopharyngitis
C0155818|ICD9CM|PT|465.8|Acute upper respiratory infections of other multiple sites
C0155818|ICD9CM|AB|465.8|Acute uri mult sites NEC
C0155820|ICD9CM|HT|466|Acute bronchitis and bronchiolitis
C0155822|ICD9CM|PT|471.1|Polypoid sinus degeneration
C0155822|ICD9CM|AB|471.1|Polypoid sinus degen
C0155823|ICD9CM|PT|471.8|Other polyp of sinus
C0155823|ICD9CM|AB|471.8|Nasal sinus polyp NEC
C0155824|ICD9CM|HT|472|Chronic pharyngitis and nasopharyngitis
C0155825|ICD9CM|AB|472.1|Chronic pharyngitis
C0155825|ICD9CM|PT|472.1|Chronic pharyngitis
C0155826|ICD9CM|AB|472.2|Chronic nasopharyngitis
C0155826|ICD9CM|PT|472.2|Chronic nasopharyngitis
C0155828|ICD9CM|PT|474.9|Unspecified chronic disease of tonsils and adenoids
C0155828|ICD9CM|HT|474|Chronic disease of tonsils and adenoids
C0155828|ICD9CM|AB|474.9|Chr T & A dis NOS
C0155829|ICD9CM|HT|474.1|Hypertrophy of tonsils and adenoids
C0155829|ICD9CM|PT|474.10|Hypertrophy of tonsil with adenoids
C0155829|ICD9CM|AB|474.10|Hypertrophy T and A
C0155831|ICD9CM|PT|474.11|Hypertrophy of tonsils alone
C0155831|ICD9CM|AB|474.11|Hypertrophy tonsils
C0155833|ICD9CM|AB|474.2|Adenoid vegetations
C0155833|ICD9CM|PT|474.2|Adenoid vegetations
C0155834|ICD9CM|PT|474.8|Other chronic disease of tonsils and adenoids
C0155834|ICD9CM|AB|474.8|Chr T & A dis NEC
C0155835|ICD9CM|HT|476|Chronic laryngitis and laryngotracheitis
C0155836|ICD9CM|AB|476.0|Chronic laryngitis
C0155836|ICD9CM|PT|476.0|Chronic laryngitis
C0155837|ICD9CM|PT|476.1|Chronic laryngotracheitis
C0155837|ICD9CM|AB|476.1|Chr laryngotracheitis
C0155839|ICD9CM|PT|478.9|Other and unspecified diseases of upper respiratory tract
C0155839|ICD9CM|HT|478|Other diseases of upper respiratory tract
C0155839|ICD9CM|HT|470-478.99|OTHER DISEASES OF THE UPPER RESPIRATORY TRACT
C0155839|ICD9CM|AB|478.9|Upper resp dis NEC/NOS
C0155840|ICD9CM|PT|478.0|Hypertrophy of nasal turbinates
C0155840|ICD9CM|AB|478.0|Hypertrph nasal turbinat
C0155841|ICD9CM|PT|478.21|Cellulitis of pharynx or nasopharynx
C0155841|ICD9CM|AB|478.21|Cellulitis of pharynx
C0155842|ICD9CM|AB|478.22|Parapharyngeal abscess
C0155842|ICD9CM|PT|478.22|Parapharyngeal abscess
C0155843|ICD9CM|AB|478.24|Retropharyngeal abscess
C0155843|ICD9CM|PT|478.24|Retropharyngeal abscess
C0155844|ICD9CM|PT|478.25|Edema of pharynx or nasopharynx
C0155844|ICD9CM|AB|478.25|Edema pharynx/nasopharyx
C0155845|ICD9CM|PT|478.26|Cyst of pharynx or nasopharynx
C0155845|ICD9CM|AB|478.26|Cyst pharynx/nasopharynx
C0155847|ICD9CM|PT|478.31|Unilateral paralysis of vocal cords or larynx, partial
C0155847|ICD9CM|AB|478.31|Vocal paral unilat part
C0155848|ICD9CM|PT|478.32|Unilateral paralysis of vocal cords or larynx, complete
C0155848|ICD9CM|AB|478.32|Vocal paral unilat total
C0155849|ICD9CM|PT|478.33|Bilateral paralysis of vocal cords or larynx, partial
C0155849|ICD9CM|AB|478.33|Vocal paral bilat part
C0155850|ICD9CM|PT|478.34|Bilateral paralysis of vocal cords or larynx, complete
C0155850|ICD9CM|AB|478.34|Vocal paral bilat total
C0155851|ICD9CM|PT|478.4|Polyp of vocal cord or larynx
C0155851|ICD9CM|AB|478.4|Vocal cord/larynx polyp
C0155852|ICD9CM|PT|478.5|Other diseases of vocal cords
C0155852|ICD9CM|AB|478.5|Vocal cord disease NEC
C0155853|ICD9CM|PT|478.71|Cellulitis and perichondritis of larynx
C0155853|ICD9CM|AB|478.71|Laryngeal cellulitis
C0155858|ICD9CM|HT|482|Other bacterial pneumonia
C0155860|ICD9CM|PT|482.1|Pneumonia due to Pseudomonas
C0155860|ICD9CM|AB|482.1|Pseudomonal pneumonia
C0155862|ICD9CM|AB|481|Pneumococcal pneumonia
C0155862|ICD9CM|HT|482.3|Pneumonia due to Streptococcus
C0155862|ICD9CM|PT|482.30|Pneumonia due to Streptococcus, unspecified
C0155862|ICD9CM|PT|481|Pneumococcal pneumonia [Streptococcus pneumoniae pneumonia]
C0155862|ICD9CM|AB|482.30|Streptococcal pneumn NOS
C0155863|ICD9CM|HT|484|Pneumonia in infectious diseases classified elsewhere
C0155865|ICD9CM|PT|484.3|Pneumonia in whooping cough
C0155865|ICD9CM|AB|484.3|Pneumonia in whoop cough
C0155866|ICD9CM|AB|022.1|Pulmonary anthrax
C0155866|ICD9CM|PT|022.1|Pulmonary anthrax
C0155866|ICD9CM|AB|484.5|Pneumonia in anthrax
C0155866|ICD9CM|PT|484.5|Pneumonia in anthrax
C0155867|ICD9CM|PT|484.6|Pneumonia in aspergillosis
C0155867|ICD9CM|AB|484.6|Pneum in aspergillosis
C0155868|ICD9CM|PT|484.7|Pneumonia in other systemic mycoses
C0155868|ICD9CM|AB|484.7|Pneum in oth sys mycoses
C0155869|ICD9CM|PT|484.8|Pneumonia in other infectious diseases classified elsewhere
C0155869|ICD9CM|AB|484.8|Pneum in infect dis NEC
C0155870|ICD9CM|HT|480-488.99|PNEUMONIA AND INFLUENZA
C0155870|ICD9CM|AB|487.0|Influenza with pneumonia
C0155870|ICD9CM|PT|487.0|Influenza with pneumonia
C0155871|ICD9CM|PT|487.8|Influenza with other manifestations
C0155871|ICD9CM|AB|487.8|Flu w manifestation NEC
C0155872|ICD9CM|PT|491.0|Simple chronic bronchitis
C0155872|ICD9CM|AB|491.0|Simple chr bronchitis
C0155873|ICD9CM|PT|491.1|Mucopurulent chronic bronchitis
C0155873|ICD9CM|AB|491.1|Mucopurul chr bronchitis
C0155874|ICD9CM|HT|491.2|Obstructive chronic bronchitis
C0155875|ICD9CM|PT|491.20|Obstructive chronic bronchitis without exacerbation
C0155875|ICD9CM|AB|491.20|Obst chr bronc w/o exac
C0155877|ICD9CM|HT|493.0|Extrinsic asthma
C0155878|ICD9CM|AB|493.00|Extrinsic asthma NOS
C0155878|ICD9CM|PT|493.00|Extrinsic asthma, unspecified
C0155879|ICD9CM|PT|493.01|Extrinsic asthma with status asthmaticus
C0155879|ICD9CM|AB|493.01|Ext asthma w status asth
C0155880|ICD9CM|HT|493.1|Intrinsic asthma
C0155881|ICD9CM|AB|493.10|Intrinsic asthma NOS
C0155881|ICD9CM|PT|493.10|Intrinsic asthma, unspecified
C0155882|ICD9CM|PT|493.11|Intrinsic asthma with status asthmaticus
C0155882|ICD9CM|AB|493.11|Int asthma w status asth
C0155883|ICD9CM|HT|493.2|Chronic obstructive asthma
C0155886|ICD9CM|AB|493.90|Asthma NOS
C0155886|ICD9CM|PT|493.90|Asthma, unspecified type, unspecified
C0155888|ICD9CM|AB|495.4|Malt workers' lung
C0155888|ICD9CM|PT|495.4|Malt workers' lung
C0155889|ICD9CM|AB|495.5|Mushroom workers' lung
C0155889|ICD9CM|PT|495.5|Mushroom workers' lung
C0155890|ICD9CM|PT|495.6|Maple bark-strippers' lung
C0155890|ICD9CM|AB|495.6|Mapl bark-stripprs' lung
C0155891|ICD9CM|PT|495.7|"Ventilation" pneumonitis
C0155891|ICD9CM|AB|495.7|"ventilation" pneumonit
C0155892|ICD9CM|PT|495.8|Other specified allergic alveolitis and pneumonitis
C0155892|ICD9CM|AB|495.8|Allerg alveol/pneum NEC
C0155893|ICD9CM|HT|506|Respiratory conditions due to chemical fumes and vapors
C0155894|ICD9CM|PT|506.0|Bronchitis and pneumonitis due to fumes and vapors
C0155894|ICD9CM|AB|506.0|Fum/vapor bronc/pneumon
C0155895|ICD9CM|PT|506.1|Acute pulmonary edema due to fumes and vapors
C0155895|ICD9CM|AB|506.1|Fum/vapor ac pulm edema
C0155896|ICD9CM|PT|506.2|Upper respiratory inflammation due to fumes and vapors
C0155896|ICD9CM|AB|506.2|Fum/vapor up resp inflam
C0155897|ICD9CM|PT|506.3|Other acute and subacute respiratory conditions due to fumes and vapors
C0155897|ICD9CM|AB|506.3|Fum/vap ac resp cond NEC
C0155898|ICD9CM|PT|506.4|Chronic respiratory conditions due to fumes and vapors
C0155898|ICD9CM|AB|506.4|Fum/vapor chr resp cond
C0155899|ICD9CM|HT|507|Pneumonitis due to solids and liquids
C0155900|ICD9CM|PT|507.8|Pneumonitis due to other solids and liquids
C0155900|ICD9CM|AB|507.8|Solid/liq pneumonit NEC
C0155901|ICD9CM|HT|508|Respiratory conditions due to other and unspecified external agents
C0155902|ICD9CM|PT|508.0|Acute pulmonary manifestations due to radiation
C0155902|ICD9CM|AB|508.0|Ac pul manif d/t radiat
C0155903|ICD9CM|PT|508.1|Chronic and other pulmonary manifestations due to radiation
C0155903|ICD9CM|AB|508.1|Chr pul manif d/t radiat
C0155904|ICD9CM|PT|508.8|Respiratory conditions due to other specified external agents
C0155904|ICD9CM|AB|508.8|Resp cond: ext agent NEC
C0155905|ICD9CM|PT|508.9|Respiratory conditions due to unspecified external agent
C0155905|ICD9CM|AB|508.9|Resp cond: ext agent NOS
C0155906|ICD9CM|PT|511.1|Pleurisy with effusion, with mention of a bacterial cause other than tuberculosis
C0155906|ICD9CM|AB|511.1|Bact pleur/effus not TB
C0155907|ICD9CM|PT|512.0|Spontaneous tension pneumothorax
C0155907|ICD9CM|AB|512.0|Spont tens pneumothorax
C0155908|ICD9CM|HT|513|Abscess of lung and mediastinum
C0155909|ICD9CM|AB|513.1|Abscess of mediastinum
C0155909|ICD9CM|PT|513.1|Abscess of mediastinum
C0155910|ICD9CM|PT|514|Pulmonary congestion and hypostasis
C0155910|ICD9CM|AB|514|Pulm congest/hypostasis
C0155912|ICD9CM|PT|516.2|Pulmonary alveolar microlithiasis
C0155912|ICD9CM|AB|516.2|Pulm alveolar microlith
C0155913|ICD9CM|PT|516.8|Other specified alveolar and parietoalveolar pneumonopathies
C0155913|ICD9CM|AB|516.8|Alveol pneumonopathy NEC
C0155914|ICD9CM|PT|516.9|Unspecified alveolar and parietoalveolar pneumonopathy
C0155914|ICD9CM|AB|516.9|Alveol pneumonopathy NOS
C0155915|ICD9CM|HT|517|Lung involvement in conditions classified elsewhere
C0155917|ICD9CM|PT|517.8|Lung involvement in other diseases classified elsewhere
C0155917|ICD9CM|AB|517.8|Lung involv in oth dis
C0155918|ICD9CM|AB|518.2|Compensatory emphysema
C0155918|ICD9CM|PT|518.2|Compensatory emphysema
C0155919|ICD9CM|PT|518.4|Acute edema of lung, unspecified
C0155919|ICD9CM|AB|518.4|Acute lung edema NOS
C0155921|ICD9CM|HT|519.0|Tracheostomy complications
C0155921|ICD9CM|PT|519.00|Tracheostomy complication, unspecified
C0155921|ICD9CM|AB|519.00|Tracheostomy comp NOS
C0155922|ICD9CM|PT|520.9|Unspecified disorder of tooth development and eruption
C0155922|ICD9CM|HT|520|Disorders of tooth development and eruption
C0155922|ICD9CM|AB|520.9|Tooth devel/erup dis NOS
C0155924|ICD9CM|PT|520.8|Other specified disorders of tooth development and eruption
C0155924|ICD9CM|AB|520.8|Tooth devel/erup dis NEC
C0155926|ICD9CM|HT|521|Diseases of hard tissues of teeth
C0155926|ICD9CM|PT|521.9|Unspecified disease of hard tissues of teeth
C0155926|ICD9CM|AB|521.9|Hard tiss dis teeth NOS
C0155930|ICD9CM|AB|521.6|Ankylosis of teeth
C0155930|ICD9CM|PT|521.6|Ankylosis of teeth
C0155933|ICD9CM|HT|522|Diseases of pulp and periapical tissues
C0155934|ICD9CM|PT|522.4|Acute apical periodontitis of pulpal origin
C0155934|ICD9CM|AB|522.4|Ac apical periodontitis
C0155935|ICD9CM|PT|522.9|Other and unspecified diseases of pulp and periapical tissues
C0155935|ICD9CM|AB|522.9|Pulp/periapical dis NEC
C0155936|ICD9CM|HT|523|Gingival and periodontal diseases
C0155936|ICD9CM|PT|523.9|Unspecified gingival and periodontal disease
C0155936|ICD9CM|AB|523.9|Gingiv/periodont dis NOS
C0155937|ICD9CM|HT|523.0|Acute gingivitis
C0155938|ICD9CM|HT|524|Dentofacial anomalies, including malocclusion
C0155939|ICD9CM|HT|524.2|Anomalies of dental arch relationship
C0155939|ICD9CM|AB|524.20|Anomaly dental arch NOS
C0155939|ICD9CM|PT|524.20|Unspecified anomaly of dental arch relationship
C0155940|ICD9CM|PT|524.30|Unspecified anomaly of tooth position
C0155940|ICD9CM|AB|524.30|Tooth position anom NOS
C0155942|ICD9CM|PT|524.61|Temporomandibular joint disorders, adhesions and ankylosis (bony or fibrous)
C0155942|ICD9CM|AB|524.61|Adhesns/ankylosis - TMJ
C0155943|ICD9CM|PT|524.62|Temporomandibular joint disorders, arthralgia of temporomandibular joint
C0155943|ICD9CM|AB|524.62|Arthralgia TMJ
C0155945|ICD9CM|PT|524.69|Other specified temporomandibular joint disorders
C0155945|ICD9CM|AB|524.69|Other specf TMJ disordrs
C0155946|ICD9CM|HT|524.8|Other specified dentofacial anomalies
C0155946|ICD9CM|PT|524.89|Other specified dentofacial anomalies
C0155946|ICD9CM|AB|524.89|Dentofacial anomaly NEC
C0155947|ICD9CM|AB|524.9|Dentofacial anomaly NOS
C0155947|ICD9CM|PT|524.9|Unspecified dentofacial anomalies
C0155948|ICD9CM|HT|525|Other diseases and conditions of the teeth and supporting structures
C0155949|ICD9CM|PT|525.0|Exfoliation of teeth due to systemic causes
C0155949|ICD9CM|AB|525.0|Exfoliation of teeth
C0155951|ICD9CM|HT|525.2|Atrophy of edentulous alveolar ridge
C0155952|ICD9CM|AB|525.3|Retained dental root
C0155952|ICD9CM|PT|525.3|Retained dental root
C0155954|ICD9CM|PT|526.4|Inflammatory conditions of jaw
C0155954|ICD9CM|AB|526.4|Inflammation of jaw
C0155955|ICD9CM|AB|526.81|Exostosis of jaw
C0155955|ICD9CM|PT|526.81|Exostosis of jaw
C0155956|ICD9CM|PT|527.0|Atrophy of salivary gland
C0155956|ICD9CM|AB|527.0|Salivary gland atrophy
C0155957|ICD9CM|PT|527.3|Abscess of salivary gland
C0155957|ICD9CM|AB|527.3|Salivary gland abscess
C0155958|ICD9CM|HT|528|Diseases of the oral soft tissues, excluding lesions specific for gingiva and tongue
C0155959|ICD9CM|PT|528.4|Cysts of oral soft tissues
C0155959|ICD9CM|AB|528.4|Oral soft tissue cyst
C0155961|ICD9CM|HT|528.7|Other disturbances of oral epithelium, including tongue
C0155961|ICD9CM|PT|528.79|Other disturbances of oral epithelium, including tongue
C0155961|ICD9CM|AB|528.79|Dist oral epithelium NEC
C0155962|ICD9CM|HT|529|Diseases and other conditions of the tongue
C0155963|ICD9CM|PT|529.2|Median rhomboid glossitis
C0155963|ICD9CM|AB|529.2|Med rhomboid glossitis
C0155964|ICD9CM|PT|529.4|Atrophy of tongue papillae
C0155964|ICD9CM|AB|529.4|Atrophy tongue papillae
C0155965|ICD9CM|PT|529.8|Other specified conditions of the tongue
C0155965|ICD9CM|AB|529.8|Tongue disorder NEC
C0155966|ICD9CM|PT|530.6|Diverticulum of esophagus, acquired
C0155966|ICD9CM|AB|530.6|Acq esophag diverticulum
C0155967|ICD9CM|HT|531.0|Acute gastric ulcer with hemorrhage
C0155968|ICD9CM|PT|531.00|Acute gastric ulcer with hemorrhage, without mention of obstruction
C0155968|ICD9CM|AB|531.00|Ac stomach ulcer w hem
C0155969|ICD9CM|PT|531.01|Acute gastric ulcer with hemorrhage, with obstruction
C0155969|ICD9CM|AB|531.01|Ac stomac ulc w hem-obst
C0155970|ICD9CM|HT|531.1|Acute gastric ulcer with perforation
C0155971|ICD9CM|PT|531.10|Acute gastric ulcer with perforation, without mention of obstruction
C0155971|ICD9CM|AB|531.10|Ac stomach ulcer w perf
C0155972|ICD9CM|PT|531.11|Acute gastric ulcer with perforation, with obstruction
C0155972|ICD9CM|AB|531.11|Ac stom ulc w perf-obst
C0155973|ICD9CM|HT|531.2|Acute gastric ulcer with hemorrhage and perforation
C0155975|ICD9CM|PT|531.21|Acute gastric ulcer with hemorrhage and perforation, with obstruction
C0155975|ICD9CM|AB|531.21|Ac stom ulc hem/perf-obs
C0155978|ICD9CM|PT|531.31|Acute gastric ulcer without mention of hemorrhage or perforation, with obstruction
C0155978|ICD9CM|AB|531.31|Ac stomach ulc NOS-obstr
C0155979|ICD9CM|HT|531.4|Chronic or unspecified gastric ulcer with hemorrhage
C0155980|ICD9CM|PT|531.40|Chronic or unspecified gastric ulcer with hemorrhage, without mention of obstruction
C0155980|ICD9CM|AB|531.40|Chr stomach ulc w hem
C0155981|ICD9CM|PT|531.41|Chronic or unspecified gastric ulcer with hemorrhage, with obstruction
C0155981|ICD9CM|AB|531.41|Chr stom ulc w hem-obstr
C0155982|ICD9CM|HT|531.5|Chronic or unspecified gastric ulcer with perforation
C0155983|ICD9CM|PT|531.50|Chronic or unspecified gastric ulcer with perforation, without mention of obstruction
C0155983|ICD9CM|AB|531.50|Chr stomach ulcer w perf
C0155984|ICD9CM|PT|531.51|Chronic or unspecified gastric ulcer with perforation, with obstruction
C0155984|ICD9CM|AB|531.51|Chr stom ulc w perf-obst
C0155986|ICD9CM|PT|531.60|Chronic or unspecified gastric ulcer with hemorrhage and perforation, without mention of obstruction
C0155986|ICD9CM|AB|531.60|Chr stomach ulc hem/perf
C0155987|ICD9CM|PT|531.61|Chronic or unspecified gastric ulcer with hemorrhage and perforation, with obstruction
C0155987|ICD9CM|AB|531.61|Chr stom ulc hem/perf-ob
C0155989|ICD9CM|PT|531.70|Chronic gastric ulcer without mention of hemorrhage or perforation, without mention of obstruction
C0155989|ICD9CM|AB|531.70|Chr stomach ulcer NOS
C0155991|ICD9CM|PT|531.91|Gastric ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation, with obstruction
C0155991|ICD9CM|AB|531.91|Stomach ulcer NOS-obstr
C0155992|ICD9CM|HT|532.0|Acute duodenal ulcer with hemorrhage
C0155993|ICD9CM|PT|532.00|Acute duodenal ulcer with hemorrhage, without mention of obstruction
C0155993|ICD9CM|AB|532.00|Ac duodenal ulcer w hem
C0155994|ICD9CM|PT|532.01|Acute duodenal ulcer with hemorrhage, with obstruction
C0155994|ICD9CM|AB|532.01|Ac duoden ulc w hem-obst
C0155995|ICD9CM|HT|532.1|Acute duodenal ulcer with perforation
C0155997|ICD9CM|PT|532.11|Acute duodenal ulcer with perforation, with obstruction
C0155997|ICD9CM|AB|532.11|Ac duoden ulc perf-obstr
C0155998|ICD9CM|HT|532.2|Acute duodenal ulcer with hemorrhage and perforation
C0155999|ICD9CM|PT|532.20|Acute duodenal ulcer with hemorrhage and perforation, without mention of obstruction
C0155999|ICD9CM|AB|532.20|Ac duoden ulc w hem/perf
C0156000|ICD9CM|PT|532.21|Acute duodenal ulcer with hemorrhage and perforation, with obstruction
C0156000|ICD9CM|AB|532.21|Ac duod ulc hem/perf-obs
C0156001|ICD9CM|HT|532.3|Acute duodenal ulcer without mention of hemorrhage or perforation
C0156002|ICD9CM|PT|532.30|Acute duodenal ulcer without mention of hemorrhage or perforation, without mention of obstruction
C0156002|ICD9CM|AB|532.30|Acute duodenal ulcer NOS
C0156003|ICD9CM|PT|532.31|Acute duodenal ulcer without mention of hemorrhage or perforation, with obstruction
C0156003|ICD9CM|AB|532.31|Ac duodenal ulc NOS-obst
C0156004|ICD9CM|HT|532.4|Chronic or unspecified duodenal ulcer with hemorrhage
C0156005|ICD9CM|PT|532.40|Chronic or unspecified duodenal ulcer with hemorrhage, without mention of obstruction
C0156005|ICD9CM|AB|532.40|Chr duoden ulcer w hem
C0156006|ICD9CM|PT|532.41|Chronic or unspecified duodenal ulcer with hemorrhage, with obstruction
C0156006|ICD9CM|AB|532.41|Chr duoden ulc hem-obstr
C0156008|ICD9CM|PT|532.50|Chronic or unspecified duodenal ulcer with perforation, without mention of obstruction
C0156008|ICD9CM|AB|532.50|Chr duoden ulcer w perf
C0156009|ICD9CM|PT|532.51|Chronic or unspecified duodenal ulcer with perforation, with obstruction
C0156009|ICD9CM|AB|532.51|Chr duoden ulc perf-obst
C0156011|ICD9CM|PT|532.60|Chronic or unspecified duodenal ulcer with hemorrhage and perforation, without mention of obstruction
C0156011|ICD9CM|AB|532.60|Chr duoden ulc hem/perf
C0156012|ICD9CM|PT|532.61|Chronic or unspecified duodenal ulcer with hemorrhage and perforation, with obstruction
C0156012|ICD9CM|AB|532.61|Chr duod ulc hem/perf-ob
C0156014|ICD9CM|PT|532.70|Chronic duodenal ulcer without mention of hemorrhage or perforation, without mention of obstruction
C0156014|ICD9CM|AB|532.70|Chr duodenal ulcer NOS
C0156015|ICD9CM|PT|532.71|Chronic duodenal ulcer without mention of hemorrhage or perforation, with obstruction
C0156015|ICD9CM|AB|532.71|Chr duoden ulc NOS-obstr
C0156016|ICD9CM|PT|532.91|Duodenal ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation, with obstruction
C0156016|ICD9CM|AB|532.91|Duodenal ulcer NOS-obstr
C0156019|ICD9CM|PT|533.01|Acute peptic ulcer of unspecified site with hemorrhage, with obstruction
C0156019|ICD9CM|AB|533.01|Ac peptic ulc w hem-obst
C0156022|ICD9CM|PT|533.11|Acute peptic ulcer of unspecified site with perforation, with obstruction
C0156022|ICD9CM|AB|533.11|Ac peptic ulc w perf-obs
C0156024|ICD9CM|PT|533.31|Acute peptic ulcer of unspecified site without mention of hemorrhage and perforation, with obstruction
C0156024|ICD9CM|PT|533.20|Acute peptic ulcer of unspecified site with hemorrhage and perforation, without mention of obstruction
C0156024|ICD9CM|AB|533.31|Ac peptic ulcer NOS-obst
C0156024|ICD9CM|AB|533.20|Ac peptic ulc w hem/perf
C0156025|ICD9CM|PT|533.21|Acute peptic ulcer of unspecified site with hemorrhage and perforation, with obstruction
C0156025|ICD9CM|AB|533.21|Ac pept ulc hem/perf-obs
C0156029|ICD9CM|PT|533.40|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage, without mention of obstruction
C0156029|ICD9CM|AB|533.40|Chr peptic ulcer w hem
C0156030|ICD9CM|PT|533.41|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage, with obstruction
C0156030|ICD9CM|AB|533.41|Chr peptic ulc w hem-obs
C0156032|ICD9CM|PT|533.50|Chronic or unspecified peptic ulcer of unspecified site with perforation, without mention of obstruction
C0156032|ICD9CM|AB|533.50|Chr peptic ulcer w perf
C0156033|ICD9CM|PT|533.51|Chronic or unspecified peptic ulcer of unspecified site with perforation, with obstruction
C0156033|ICD9CM|AB|533.51|Chr peptic ulc perf-obst
C0156035|ICD9CM|PT|533.60|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage and perforation, without mention of obstruction
C0156035|ICD9CM|AB|533.60|Chr pept ulc w hem/perf
C0156036|ICD9CM|PT|533.61|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage and perforation, with obstruction
C0156036|ICD9CM|AB|533.61|Chr pept ulc hem/perf-ob
C0156039|ICD9CM|PT|533.71|Chronic peptic ulcer of unspecified site without mention of hemorrhage or perforation, with obstruction
C0156039|ICD9CM|AB|533.71|Chr peptic ulcer NOS-obs
C0156040|ICD9CM|PT|533.91|Peptic ulcer of unspecified site, unspecified as acute or chronic, without mention of hemorrhage or perforation, with obstruction
C0156040|ICD9CM|AB|533.91|Peptic ulcer NOS-obstruc
C0156042|ICD9CM|HT|534.0|Acute gastrojejunal ulcer with hemorrhage
C0156043|ICD9CM|PT|534.00|Acute gastrojejunal ulcer with hemorrhage, without mention of obstruction
C0156043|ICD9CM|AB|534.00|Ac marginal ulcer w hem
C0156044|ICD9CM|PT|534.01|Acute gastrojejunal ulcer, with hemorrhage, with obstruction
C0156044|ICD9CM|AB|534.01|Ac margin ulc w hem-obst
C0156045|ICD9CM|HT|534.1|Acute gastrojejunal ulcer with perforation
C0156046|ICD9CM|PT|534.10|Acute gastrojejunal ulcer with perforation, without mention of obstruction
C0156046|ICD9CM|AB|534.10|Ac marginal ulcer w perf
C0156047|ICD9CM|PT|534.11|Acute gastrojejunal ulcer with perforation, with obstruction
C0156047|ICD9CM|AB|534.11|Ac margin ulc w perf-obs
C0156048|ICD9CM|HT|534.2|Acute gastrojejunal ulcer with hemorrhage and perforation
C0156049|ICD9CM|PT|534.20|Acute gastrojejunal ulcer with hemorrhage and perforation, without mention of obstruction
C0156049|ICD9CM|AB|534.20|Ac margin ulc w hem/perf
C0156050|ICD9CM|PT|534.21|Acute gastrojejunal ulcer with hemorrhage and perforation, with obstruction
C0156050|ICD9CM|AB|534.21|Ac marg ulc hem/perf-obs
C0156053|ICD9CM|PT|534.31|Acute gastrojejunal ulcer without mention of hemorrhage or perforation, with obstruction
C0156053|ICD9CM|AB|534.31|Ac marginal ulc NOS-obst
C0156054|ICD9CM|HT|534.4|Chronic or unspecified gastrojejunal ulcer with hemorrhage
C0156055|ICD9CM|PT|534.40|Chronic or unspecified gastrojejunal ulcer with hemorrhage, without mention of obstruction
C0156055|ICD9CM|AB|534.40|Chr marginal ulcer w hem
C0156056|ICD9CM|PT|534.41|Chronic or unspecified gastrojejunal ulcer, with hemorrhage, with obstruction
C0156056|ICD9CM|AB|534.41|Chr margin ulc w hem-obs
C0156057|ICD9CM|HT|534.5|Chronic or unspecified gastrojejunal ulcer with perforation
C0156058|ICD9CM|PT|534.50|Chronic or unspecified gastrojejunal ulcer with perforation, without mention of obstruction
C0156058|ICD9CM|AB|534.50|Chr marginal ulc w perf
C0156059|ICD9CM|PT|534.51|Chronic or unspecified gastrojejunal ulcer with perforation, with obstruction
C0156059|ICD9CM|AB|534.51|Chr margin ulc perf-obst
C0156061|ICD9CM|PT|534.60|Chronic or unspecified gastrojejunal ulcer with hemorrhage and perforation, without mention of obstruction
C0156061|ICD9CM|AB|534.60|Chr margin ulc hem/perf
C0156062|ICD9CM|PT|534.61|Chronic or unspecified gastrojejunal ulcer with hemorrhage and perforation, with obstruction
C0156062|ICD9CM|AB|534.61|Chr marg ulc hem/perf-ob
C0156065|ICD9CM|PT|534.71|Chronic gastrojejunal ulcer without mention of hemorrhage or perforation, with obstruction
C0156065|ICD9CM|AB|534.71|Chr marginal ulc NOS-obs
C0156067|ICD9CM|PT|534.90|Gastrojejunal ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation, without mention of obstruction
C0156067|ICD9CM|AB|534.90|Gastrojejunal ulcer NOS
C0156068|ICD9CM|PT|534.91|Gastrojejunal ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation, with obstruction
C0156068|ICD9CM|AB|534.91|Gastrojejun ulc NOS-obst
C0156070|ICD9CM|PT|535.00|Acute gastritis, without mention of hemorrhage
C0156070|ICD9CM|AB|535.00|Acute gastrtis w/o hmrhg
C0156072|ICD9CM|PT|535.10|Atrophic gastritis, without mention of hemorrhage
C0156072|ICD9CM|AB|535.10|Atrph gastrtis w/o hmrhg
C0156073|ICD9CM|PT|535.11|Atrophic gastritis, with hemorrhage
C0156073|ICD9CM|AB|535.11|Atrph gastritis w hmrhg
C0156074|ICD9CM|PT|535.20|Gastric mucosal hypertrophy, without mention of hemorrhage
C0156074|ICD9CM|AB|535.20|Gstr mcsl hyprt w/o hmrg
C0156075|ICD9CM|PT|535.21|Gastric mucosal hypertrophy, with hemorrhage
C0156075|ICD9CM|AB|535.21|Gstr mcsl hyprt w hmrg
C0156076|ICD9CM|HT|535.3|Alcoholic gastritis
C0156077|ICD9CM|PT|535.30|Alcoholic gastritis, without mention of hemorrhage
C0156077|ICD9CM|AB|535.30|Alchl gastrtis w/o hmrhg
C0156078|ICD9CM|PT|535.31|Alcoholic gastritis, with hemorrhage
C0156078|ICD9CM|AB|535.31|Alchl gstritis w hmrhg
C0156079|ICD9CM|PT|535.40|Other specified gastritis, without mention of hemorrhage
C0156079|ICD9CM|AB|535.40|Oth spf gstrt w/o hmrhg
C0156080|ICD9CM|PT|535.41|Other specified gastritis, with hemorrhage
C0156080|ICD9CM|AB|535.41|Oth spf gastrt w hmrhg
C0156081|ICD9CM|PT|535.50|Unspecified gastritis and gastroduodenitis, without mention of hemorrhage
C0156081|ICD9CM|AB|535.50|Gstr/ddnts NOS w/o hmrhg
C0156082|ICD9CM|PT|535.51|Unspecified gastritis and gastroduodenitis, with hemorrhage
C0156082|ICD9CM|AB|535.51|Gstr/ddnts NOS w hmrhg
C0156083|ICD9CM|PT|535.60|Duodenitis, without mention of hemorrhage
C0156083|ICD9CM|AB|535.60|Duodenitis w/o hmrhg
C0156084|ICD9CM|HT|536|Disorders of function of stomach
C0156084|ICD9CM|PT|536.9|Unspecified functional disorder of stomach
C0156084|ICD9CM|AB|536.9|Stomach function dis NOS
C0156086|ICD9CM|HT|537|Other disorders of stomach and duodenum
C0156087|ICD9CM|AB|537.2|Chronic duodenal ileus
C0156087|ICD9CM|PT|537.2|Chronic duodenal ileus
C0156088|ICD9CM|AB|537.5|Gastroptosis
C0156088|ICD9CM|PT|537.5|Gastroptosis
C0156090|ICD9CM|PT|537.82|Angiodysplasia of stomach and duodenum without mention of hemorrhage
C0156090|ICD9CM|AB|537.82|Angio stm/dudn w/o hmrhg
C0156091|ICD9CM|PT|537.83|Angiodysplasia of stomach and duodenum with hemorrhage
C0156091|ICD9CM|AB|537.83|Angio stm/dudn w hmrhg
C0156092|ICD9CM|PT|540.0|Acute appendicitis with generalized peritonitis
C0156092|ICD9CM|AB|540.0|Ac append w peritonitis
C0156093|ICD9CM|PT|540.1|Acute appendicitis with peritoneal abscess
C0156093|ICD9CM|AB|540.1|Abscess of appendix
C0156094|ICD9CM|PT|540.9|Acute appendicitis without mention of peritonitis
C0156094|ICD9CM|AB|540.9|Acute appendicitis NOS
C0156095|ICD9CM|AB|542|Other appendicitis
C0156095|ICD9CM|PT|542|Other appendicitis
C0156098|ICD9CM|PT|543.9|Other and unspecified diseases of appendix
C0156098|ICD9CM|HT|543|Other diseases of appendix
C0156098|ICD9CM|AB|543.9|Diseases of appendix NEC
C0156099|ICD9CM|HT|550.0|Inguinal hernia, with gangrene
C0156100|ICD9CM|PT|550.00|Inguinal hernia, with gangrene, unilateral or unspecified (not specified as recurrent)
C0156100|ICD9CM|AB|550.00|Unilat ing hernia w gang
C0156101|ICD9CM|PT|550.01|Inguinal hernia, with gangrene, unilateral or unspecified, recurrent
C0156101|ICD9CM|AB|550.01|Recur unil ing hern-gang
C0156103|ICD9CM|PT|550.03|Inguinal hernia, with gangrene, bilateral, recurrent
C0156103|ICD9CM|AB|550.03|Recur bil ing hern-gang
C0156104|ICD9CM|HT|550.1|Inguinal hernia, with obstruction, without mention of gangrene
C0156106|ICD9CM|PT|550.11|Inguinal hernia, with obstruction, without mention of gangrene, unilateral or unspecified,recurrent
C0156106|ICD9CM|AB|550.11|Recur unil ing hern-obst
C0156109|ICD9CM|PT|550.90|Inguinal hernia, without mention of obstruction or gangrene, unilateral or unspecified (not specified as recurrent)
C0156109|ICD9CM|AB|550.90|Unilat inguinal hernia
C0156110|ICD9CM|PT|550.91|Inguinal hernia, without mention of obstruction or gangrene, unilateral or unspecified, recurrent
C0156110|ICD9CM|AB|550.91|Recur unilat inguin hern
C0156111|ICD9CM|PT|550.92|Inguinal hernia, without mention of obstruction or gangrene, bilateral (not specified as recurrent)
C0156111|ICD9CM|AB|550.92|Bilat inguinal hernia
C0156112|ICD9CM|PT|550.93|Inguinal hernia, without mention of obstruction or gangrene, bilateral, recurrent
C0156112|ICD9CM|AB|550.93|Recur bilat inguin hern
C0156113|ICD9CM|HT|551|Other hernia of abdominal cavity, with gangrene
C0156114|ICD9CM|HT|551.0|Femoral hernia with gangrene
C0156115|ICD9CM|PT|551.00|Femoral hernia with gangrene, unilateral or unspecified (not specified as recurrent)
C0156115|ICD9CM|AB|551.00|Unil femoral hern w gang
C0156116|ICD9CM|PT|551.01|Femoral hernia with gangrene, unilateral or unspecified, recurrent
C0156116|ICD9CM|AB|551.01|Rec unil fem hern w gang
C0156117|ICD9CM|AB|551.02|Bilat fem hern w gang
C0156117|ICD9CM|PT|551.02|Femoral hernia with gangrene, bilateral (not specified as recurrent)
C0156118|ICD9CM|PT|551.03|Femoral hernia with gangrene, bilateral, recurrent
C0156118|ICD9CM|AB|551.03|Recur bil fem hern-gang
C0156119|ICD9CM|PT|551.1|Umbilical hernia with gangrene
C0156119|ICD9CM|AB|551.1|Umbilical hernia w gangr
C0156120|ICD9CM|HT|551.2|Ventral hernia with gangrene
C0156120|ICD9CM|PT|551.20|Ventral hernia, unspecified, with gangrene
C0156120|ICD9CM|AB|551.20|Gangr ventral hernia NOS
C0156122|ICD9CM|PT|551.21|Incisional ventral hernia, with gangrene
C0156122|ICD9CM|AB|551.21|Gangr incisional hernia
C0156123|ICD9CM|PT|551.29|Other ventral hernia with gangrene
C0156123|ICD9CM|AB|551.29|Gang ventral hernia NEC
C0156124|ICD9CM|PT|551.3|Diaphragmatic hernia with gangrene
C0156124|ICD9CM|AB|551.3|Diaphragm hernia w gangr
C0156125|ICD9CM|PT|551.8|Hernia of other specified sites, with gangrene
C0156125|ICD9CM|AB|551.8|Hernia, site NEC w gangr
C0156127|ICD9CM|HT|552|Other hernia of abdominal cavity, with obstruction, but without mention of gangrene
C0156128|ICD9CM|HT|552.0|Femoral hernia with obstruction
C0156129|ICD9CM|PT|552.00|Femoral hernia with obstruction, unilateral or unspecified (not specified as recurrent)
C0156129|ICD9CM|AB|552.00|Unil femoral hern w obst
C0156130|ICD9CM|PT|552.01|Femoral hernia with obstruction, unilateral or unspecified, recurrent
C0156130|ICD9CM|AB|552.01|Rec unil fem hern w obst
C0156131|ICD9CM|PT|552.02|Femoral hernia with obstruction, bilateral (not specified as recurrent)
C0156131|ICD9CM|AB|552.02|Bil femoral hern w obstr
C0156133|ICD9CM|PT|552.1|Umbilical hernia with obstruction
C0156133|ICD9CM|AB|552.1|Umbilical hernia w obstr
C0156137|ICD9CM|PT|552.29|Other ventral hernia with obstruction
C0156137|ICD9CM|AB|552.29|Obstr ventral hernia NEC
C0156139|ICD9CM|PT|552.8|Hernia of other specified sites, with obstruction
C0156139|ICD9CM|AB|552.8|Hernia, site NEC w obstr
C0156140|ICD9CM|PT|552.9|Hernia of unspecified site, with obstruction
C0156140|ICD9CM|AB|552.9|Hernia, site NOS w obstr
C0156141|ICD9CM|HT|553|Other hernia of abdominal cavity without mention of obstruction or gangrene
C0156142|ICD9CM|PT|553.01|Femoral hernia without mention of obstruction or gangrene, unilateral or unspecified, recurrent
C0156142|ICD9CM|AB|553.01|Recur unil femoral hern
C0156144|ICD9CM|PT|553.03|Femoral hernia without mention of obstruction or gangrene, bilateral,recurrent
C0156144|ICD9CM|AB|553.03|Recur bilat femoral hern
C0156145|ICD9CM|PT|553.21|Incisional hernia without mention of obstruction or gangrene
C0156145|ICD9CM|AB|553.21|Incisional hernia
C0156146|ICD9CM|PT|555.0|Regional enteritis of small intestine
C0156146|ICD9CM|AB|555.0|Reg enteritis, sm intest
C0156147|ICD9CM|PT|555.1|Regional enteritis of large intestine
C0156147|ICD9CM|AB|555.1|Reg enteritis, lg intest
C0156153|ICD9CM|PT|558.1|Gastroenteritis and colitis due to radiation
C0156153|ICD9CM|AB|558.1|Radiation gastroenterit
C0156154|ICD9CM|PT|558.2|Toxic gastroenteritis and colitis
C0156154|ICD9CM|AB|558.2|Toxic gastroenteritis
C0156156|ICD9CM|AB|560.31|Gallstone ileus
C0156156|ICD9CM|PT|560.31|Gallstone ileus
C0156157|ICD9CM|HT|560.8|Other specified intestinal obstruction
C0156157|ICD9CM|PT|560.89|Other specified intestinal obstruction
C0156157|ICD9CM|AB|560.89|Intestinal obstruct NEC
C0156158|ICD9CM|PT|560.81|Intestinal or peritoneal adhesions with obstruction (postoperative) (postinfection)
C0156158|ICD9CM|AB|560.81|Intestinal adhes w obstr
C0156162|ICD9CM|PT|562.00|Diverticulosis of small intestine (without mention of hemorrhage)
C0156162|ICD9CM|AB|562.00|Dvrtclo sml int w/o hmrg
C0156163|ICD9CM|PT|562.01|Diverticulitis of small intestine (without mention of hemorrhage)
C0156163|ICD9CM|AB|562.01|Dvrtcli sml int w/o hmrg
C0156165|ICD9CM|PT|562.03|Diverticulitis of small intestine with hemorrhage
C0156165|ICD9CM|AB|562.03|Dvrtcli sml int w hmrhg
C0156166|ICD9CM|PT|562.10|Diverticulosis of colon (without mention of hemorrhage)
C0156166|ICD9CM|AB|562.10|Dvrtclo colon w/o hmrhg
C0156167|ICD9CM|PT|562.11|Diverticulitis of colon (without mention of hemorrhage)
C0156167|ICD9CM|AB|562.11|Dvrtcli colon w/o hmrhg
C0156168|ICD9CM|PT|562.12|Diverticulosis of colon with hemorrhage
C0156168|ICD9CM|AB|562.12|Dvrtclo colon w hmrhg
C0156171|ICD9CM|PT|564.3|Vomiting following gastrointestinal surgery
C0156171|ICD9CM|AB|564.3|Vomiting post-gi surgery
C0156172|ICD9CM|PT|564.4|Other postoperative functional disorders
C0156172|ICD9CM|AB|564.4|Postop GI funct dis NEC
C0156173|ICD9CM|AB|564.5|Functional diarrhea
C0156173|ICD9CM|PT|564.5|Functional diarrhea
C0156175|ICD9CM|HT|565|Anal fissure and fistula
C0156177|ICD9CM|PT|567.0|Peritonitis in infectious diseases classified elsewhere
C0156177|ICD9CM|AB|567.0|Peritonitis in infec dis
C0156178|ICD9CM|AB|567.1|Pneumococcal peritonitis
C0156178|ICD9CM|PT|567.1|Pneumococcal peritonitis
C0156179|ICD9CM|HT|567.2|Other suppurative peritonitis
C0156179|ICD9CM|PT|567.29|Other suppurative peritonitis
C0156179|ICD9CM|AB|567.29|Suppurat peritonitis NEC
C0156180|ICD9CM|HT|568|Other disorders of peritoneum
C0156182|ICD9CM|HT|569|Other disorders of intestine
C0156183|ICD9CM|PT|569.2|Stenosis of rectum and anus
C0156183|ICD9CM|AB|569.2|Rectal & anal stenosis
C0156185|ICD9CM|PT|569.5|Abscess of intestine
C0156185|ICD9CM|AB|569.5|Intestinal abscess
C0156186|ICD9CM|HT|569.6|Colostomy and enterostomy complications
C0156186|ICD9CM|PT|569.60|Colostomy and enterostomy complication, unspecified
C0156186|ICD9CM|AB|569.60|Colstomy/enter comp NOS
C0156188|ICD9CM|PT|569.85|Angiodysplasia of intestine with hemorrhage
C0156188|ICD9CM|AB|569.85|Angio intes w hmrhg
C0156189|ICD9CM|HT|571|Chronic liver disease and cirrhosis
C0156191|ICD9CM|HT|572|Liver abscess and sequelae of chronic liver disease
C0156192|ICD9CM|AB|572.1|Portal pyemia
C0156192|ICD9CM|PT|572.1|Portal pyemia
C0156193|ICD9CM|PT|572.8|Other sequelae of chronic liver disease
C0156193|ICD9CM|AB|572.8|Oth sequela, chr liv dis
C0156194|ICD9CM|HT|573|Other disorders of liver
C0156195|ICD9CM|PT|573.0|Chronic passive congestion of liver
C0156195|ICD9CM|AB|573.0|Chr passiv congest liver
C0156196|ICD9CM|PT|573.1|Hepatitis in viral diseases classified elsewhere
C0156196|ICD9CM|AB|573.1|Hepatitis in viral dis
C0156197|ICD9CM|PT|573.2|Hepatitis in other infectious diseases classified elsewhere
C0156197|ICD9CM|AB|573.2|Hepatitis in oth inf dis
C0156199|ICD9CM|HT|574.0|Calculus of gallbladder with acute cholecystitis
C0156201|ICD9CM|PT|574.01|Calculus of gallbladder with acute cholecystitis, with obstruction
C0156201|ICD9CM|AB|574.01|Cholelith/ac gb inf-obst
C0156202|ICD9CM|HT|574.1|Calculus of gallbladder with other cholecystitis
C0156203|ICD9CM|PT|574.10|Calculus of gallbladder with other cholecystitis, without mention of obstruction
C0156203|ICD9CM|AB|574.10|Cholelith w cholecys NEC
C0156204|ICD9CM|PT|574.11|Calculus of gallbladder with other cholecystitis, with obstruction
C0156204|ICD9CM|AB|574.11|Cholelith/gb inf NEC-obs
C0156205|ICD9CM|PT|574.21|Calculus of gallbladder without mention of cholecystitis, with obstruction
C0156205|ICD9CM|AB|574.21|Cholelithias NOS w obstr
C0156206|ICD9CM|HT|574.3|Calculus of bile duct with acute cholecystitis
C0156207|ICD9CM|PT|574.30|Calculus of bile duct with acute cholecystitis, without mention of obstruction
C0156207|ICD9CM|AB|574.30|Choledocholith/ac gb inf
C0156208|ICD9CM|PT|574.31|Calculus of bile duct with acute cholecystitis, with obstruction
C0156208|ICD9CM|AB|574.31|Choledochlith/ac gb-obst
C0156209|ICD9CM|HT|574.4|Calculus of bile duct with other cholecystitis
C0156210|ICD9CM|PT|574.40|Calculus of bile duct with other cholecystitis, without mention of obstruction
C0156210|ICD9CM|AB|574.40|Choledochlith/gb inf NEC
C0156211|ICD9CM|PT|574.41|Calculus of bile duct with other cholecystitis, with obstruction
C0156211|ICD9CM|AB|574.41|Choledochlith/gb NEC-obs
C0156212|ICD9CM|PT|574.50|Calculus of bile duct without mention of cholecystitis, without mention of obstruction
C0156212|ICD9CM|AB|574.50|Choledocholithiasis NOS
C0156213|ICD9CM|HT|575|Other disorders of gallbladder
C0156214|ICD9CM|PT|575.2|Obstruction of gallbladder
C0156214|ICD9CM|AB|575.2|Obstruction gallbladder
C0156215|ICD9CM|PT|575.4|Perforation of gallbladder
C0156215|ICD9CM|AB|575.4|Perforation gallbladder
C0156216|ICD9CM|AB|575.5|Fistula of gallbladder
C0156216|ICD9CM|PT|575.5|Fistula of gallbladder
C0156217|ICD9CM|HT|576|Other disorders of biliary tract
C0156218|ICD9CM|AB|576.3|Perforation of bile duct
C0156218|ICD9CM|PT|576.3|Perforation of bile duct
C0156221|ICD9CM|HT|580|Acute glomerulonephritis
C0156223|ICD9CM|PT|580.4|Acute glomerulonephritis with lesion of rapidly progressive glomerulonephritis
C0156223|ICD9CM|AB|580.4|Ac rapidly progr nephrit
C0156224|ICD9CM|HT|580.8|Acute glomerulonephritis with other specified pathological lesion in kidney
C0156224|ICD9CM|PT|580.89|Acute glomerulonephritis with other specified pathological lesion in kidney
C0156224|ICD9CM|AB|580.89|Acute nephritis NEC
C0156225|ICD9CM|PT|580.81|Acute glomerulonephritis in diseases classified elsewhere
C0156225|ICD9CM|AB|580.81|Ac nephritis in oth dis
C0156226|ICD9CM|PT|580.9|Acute glomerulonephritis with unspecified pathological lesion in kidney
C0156226|ICD9CM|AB|580.9|Acute nephritis NOS
C0156227|ICD9CM|PT|581.0|Nephrotic syndrome with lesion of proliferative glomerulonephritis
C0156227|ICD9CM|AB|581.0|Nephrotic syn, prolifer
C0156228|ICD9CM|PT|581.1|Nephrotic syndrome with lesion of membranous glomerulonephritis
C0156228|ICD9CM|AB|581.1|Epimembranous nephritis
C0156229|ICD9CM|PT|581.2|Nephrotic syndrome with lesion of membranoproliferative glomerulonephritis
C0156229|ICD9CM|AB|581.2|Membranoprolif nephrosis
C0156230|ICD9CM|PT|581.81|Nephrotic syndrome in diseases classified elsewhere
C0156230|ICD9CM|AB|581.81|Nephrotic syn in oth dis
C0156231|ICD9CM|PT|582.0|Chronic glomerulonephritis with lesion of proliferative glomerulonephritis
C0156231|ICD9CM|AB|582.0|Chr proliferat nephritis
C0156233|ICD9CM|HT|582.8|Chronic glomerulonephritis with other specified pathological lesion in kidney
C0156233|ICD9CM|PT|582.89|Chronic glomerulonephritis with other specified pathological lesion in kidney
C0156233|ICD9CM|AB|582.89|Chronic nephritis NEC
C0156234|ICD9CM|PT|582.81|Chronic glomerulonephritis in diseases classified elsewhere
C0156234|ICD9CM|AB|582.81|Chr nephritis in oth dis
C0156235|ICD9CM|PT|582.9|Chronic glomerulonephritis with unspecified pathological lesion in kidney
C0156235|ICD9CM|AB|582.9|Chronic nephritis NOS
C0156236|ICD9CM|PT|583.0|Nephritis and nephropathy, not specified as acute or chronic, with lesion of proliferative glomerulonephritis
C0156236|ICD9CM|AB|583.0|Proliferat nephritis NOS
C0156237|ICD9CM|PT|583.4|Nephritis and nephropathy, not specified as acute or chronic, with lesion of rapidly progressive glomerulonephritis
C0156237|ICD9CM|AB|583.4|Rapidly prog nephrit NOS
C0156238|ICD9CM|PT|583.6|Nephritis and nephropathy, not specified as acute or chronic, with lesion of renal cortical necrosis
C0156238|ICD9CM|AB|583.6|Renal cort necrosis NOS
C0156239|ICD9CM|PT|583.7|Nephritis and nephropathy, not specified as acute or chronic, with lesion of renal medullary necrosis
C0156239|ICD9CM|AB|583.7|Nephr NOS/medull necros
C0156245|ICD9CM|AB|589.0|Unilateral small kidney
C0156245|ICD9CM|PT|589.0|Unilateral small kidney
C0156246|ICD9CM|AB|589.1|Bilateral small kidneys
C0156246|ICD9CM|PT|589.1|Bilateral small kidneys
C0156247|ICD9CM|AB|589.9|Small kidney NOS
C0156247|ICD9CM|HT|589|Small kidney of unknown cause
C0156247|ICD9CM|PT|589.9|Small kidney, unspecified
C0156249|ICD9CM|PT|590.00|Chronic pyelonephritis without lesion of renal medullary necrosis
C0156249|ICD9CM|AB|590.00|Chr pyelonephritis NOS
C0156250|ICD9CM|PT|590.01|Chronic pyelonephritis with lesion of renal medullary necrosis
C0156250|ICD9CM|AB|590.01|Chr pyeloneph w med necr
C0156251|ICD9CM|PT|590.10|Acute pyelonephritis without lesion of renal medullary necrosis
C0156251|ICD9CM|AB|590.10|Ac pyelonephritis NOS
C0156252|ICD9CM|PT|590.11|Acute pyelonephritis with lesion of renal medullary necrosis
C0156252|ICD9CM|AB|590.11|Ac pyelonephr w med necr
C0156253|ICD9CM|PT|590.2|Renal and perinephric abscess
C0156253|ICD9CM|AB|590.2|Renal/perirenal abscess
C0156254|ICD9CM|AB|590.3|Pyeloureteritis cystica
C0156254|ICD9CM|PT|590.3|Pyeloureteritis cystica
C0156255|ICD9CM|HT|590.8|Other pyelonephritis or pyonephrosis, not specified as acute or chronic
C0156256|ICD9CM|PT|590.81|Pyelitis or pyelonephritis in diseases classified elsewhere
C0156256|ICD9CM|AB|590.81|Pyelonephrit in oth dis
C0156257|ICD9CM|HT|592|Calculus of kidney and ureter
C0156258|ICD9CM|HT|593|Other disorders of kidney and ureter
C0156259|ICD9CM|AB|593.1|Hypertrophy of kidney
C0156259|ICD9CM|PT|593.1|Hypertrophy of kidney
C0156261|ICD9CM|PT|593.3|Stricture or kinking of ureter
C0156261|ICD9CM|AB|593.3|Stricture of ureter
C0156263|ICD9CM|AB|593.82|Ureteral fistula
C0156263|ICD9CM|PT|593.82|Ureteral fistula
C0156264|ICD9CM|HT|594|Calculus of lower urinary tract
C0156264|ICD9CM|PT|594.9|Calculus of lower urinary tract, unspecified
C0156264|ICD9CM|AB|594.9|Lower urin calcul NOS
C0156265|ICD9CM|PT|594.0|Calculus in diverticulum of bladder
C0156265|ICD9CM|AB|594.0|Blad diverticulum calcul
C0156266|ICD9CM|PT|594.8|Other lower urinary tract calculus
C0156266|ICD9CM|AB|594.8|Lower urin calcul NEC
C0156268|ICD9CM|PT|595.2|Other chronic cystitis
C0156268|ICD9CM|AB|595.2|Chronic cystitis NEC
C0156269|ICD9CM|PT|595.4|Cystitis in diseases classified elsewhere
C0156269|ICD9CM|AB|595.4|Cystitis in oth dis
C0156270|ICD9CM|AB|595.82|Irradiation cystitis
C0156270|ICD9CM|PT|595.82|Irradiation cystitis
C0156271|ICD9CM|HT|596|Other disorders of bladder
C0156272|ICD9CM|AB|596.1|Intestinovesical fistula
C0156272|ICD9CM|PT|596.1|Intestinovesical fistula
C0156273|ICD9CM|AB|596.3|Diverticulum of bladder
C0156273|ICD9CM|PT|596.3|Diverticulum of bladder
C0156274|ICD9CM|PT|596.59|Other functional disorder of bladder
C0156274|ICD9CM|HT|596.5|Other functional disorders of bladder
C0156274|ICD9CM|AB|596.59|Oth func dsdr bladder
C0156275|ICD9CM|PT|596.6|Rupture of bladder, nontraumatic
C0156275|ICD9CM|AB|596.6|Bladder rupt, nontraum
C0156276|ICD9CM|PT|596.7|Hemorrhage into bladder wall
C0156276|ICD9CM|AB|596.7|Bladder wall hemorrhage
C0156277|ICD9CM|HT|597|Urethritis, not sexually transmitted, and urethral syndrome
C0156278|ICD9CM|AB|597.0|Urethral abscess
C0156278|ICD9CM|PT|597.0|Urethral abscess
C0156279|ICD9CM|AB|597.81|Urethral syndrome NOS
C0156279|ICD9CM|PT|597.81|Urethral syndrome NOS
C0156282|ICD9CM|PT|598.01|Urethral stricture due to infective diseases classified elsewhere
C0156282|ICD9CM|AB|598.01|Ureth strict:oth infect
C0156284|ICD9CM|PT|598.2|Postoperative urethral stricture
C0156284|ICD9CM|AB|598.2|Postop urethral strictur
C0156286|ICD9CM|AB|599.4|Urethral false passage
C0156286|ICD9CM|PT|599.4|Urethral false passage
C0156287|ICD9CM|PT|599.5|Prolapsed urethral mucosa
C0156287|ICD9CM|AB|599.5|Prolapse urethral mucosa
C0156288|ICD9CM|HT|599.8|Other specified disorders of urethra and urinary tract
C0156290|ICD9CM|AB|601.2|Abscess of prostate
C0156290|ICD9CM|PT|601.2|Abscess of prostate
C0156291|ICD9CM|AB|601.3|Prostatocystitis
C0156291|ICD9CM|PT|601.3|Prostatocystitis
C0156294|ICD9CM|HT|602|Other disorders of prostate
C0156295|ICD9CM|PT|602.1|Congestion or hemorrhage of prostate
C0156295|ICD9CM|AB|602.1|Prostatic congest/hemorr
C0156296|ICD9CM|AB|602.2|Atrophy of prostate
C0156296|ICD9CM|PT|602.2|Atrophy of prostate
C0156297|ICD9CM|PT|602.8|Other specified disorders of prostate
C0156297|ICD9CM|AB|602.8|Prostatic disorders NEC
C0156299|ICD9CM|AB|603.0|Encysted hydrocele
C0156299|ICD9CM|PT|603.0|Encysted hydrocele
C0156300|ICD9CM|AB|603.1|Infected hydrocele
C0156300|ICD9CM|PT|603.1|Infected hydrocele
C0156301|ICD9CM|PT|604.0|Orchitis, epididymitis, and epididymo-orchitis, with abscess
C0156301|ICD9CM|AB|604.0|Orchitis with abscess
C0156302|ICD9CM|HT|604.9|Other orchitis, epididymitis, and epididymo-orchitis, without mention of abscess
C0156302|ICD9CM|PT|604.99|Other orchitis, epididymitis, and epididymo-orchitis, without mention of abscess
C0156302|ICD9CM|AB|604.99|Orchitis/epididymit NEC
C0156303|ICD9CM|PT|604.91|Orchitis and epididymitis in diseases classified elsewhere
C0156303|ICD9CM|AB|604.91|Orchitis in oth disease
C0156306|ICD9CM|PT|607.2|Other inflammatory disorders of penis
C0156306|ICD9CM|AB|607.2|Inflam dis, penis NEC
C0156307|ICD9CM|PT|607.82|Vascular disorders of penis
C0156307|ICD9CM|AB|607.82|Vascular disorder, penis
C0156308|ICD9CM|AB|607.83|Edema of penis
C0156308|ICD9CM|PT|607.83|Edema of penis
C0156309|ICD9CM|PT|607.84|Impotence of organic origin
C0156309|ICD9CM|AB|607.84|Impotence, organic orign
C0156311|ICD9CM|HT|608|Other disorders of male genital organs
C0156312|ICD9CM|AB|608.3|Atrophy of testis
C0156312|ICD9CM|PT|608.3|Atrophy of testis
C0156313|ICD9CM|PT|608.4|Other inflammatory disorders of male genital organs
C0156313|ICD9CM|AB|608.4|Male gen inflam dis NEC
C0156314|ICD9CM|PT|608.81|Disorders of male genital organs in diseases classified elsewhere
C0156314|ICD9CM|AB|608.81|Male gen dis in oth dis
C0156315|ICD9CM|PT|608.84|Chylocele of tunica vaginalis
C0156315|ICD9CM|AB|608.84|Chylocele, tunic vaginal
C0156316|ICD9CM|PT|608.85|Stricture of male genital organs
C0156316|ICD9CM|AB|608.85|Stricture, male gen orgn
C0156317|ICD9CM|PT|608.86|Edema of male genital organs
C0156317|ICD9CM|AB|608.86|Edema, male genital orgn
C0156318|ICD9CM|AB|610.3|Fibrosclerosis of breast
C0156318|ICD9CM|PT|610.3|Fibrosclerosis of breast
C0156319|ICD9CM|PT|610.8|Other specified benign mammary dysplasias
C0156319|ICD9CM|AB|610.8|Benign mamm dysplas NEC
C0156320|ICD9CM|HT|611|Other disorders of breast
C0156321|ICD9CM|AB|611.3|Fat necrosis of breast
C0156321|ICD9CM|PT|611.3|Fat necrosis of breast
C0156323|ICD9CM|HT|611.7|Signs and symptoms in breast
C0156324|ICD9CM|PT|611.79|Other signs and symptoms in breast
C0156324|ICD9CM|AB|611.79|Symptoms in breast NEC
C0156325|ICD9CM|PT|611.89|Other specified disorders of breast
C0156325|ICD9CM|HT|611.8|Other specified disorders of breast
C0156325|ICD9CM|AB|611.89|Disorders breast NEC
C0156326|ICD9CM|HT|614|Inflammatory disease of ovary, fallopian tube, pelvic cellular tissue, and peritoneum
C0156327|ICD9CM|PT|614.0|Acute salpingitis and oophoritis
C0156327|ICD9CM|AB|614.0|Ac salpingo-oophoritis
C0156328|ICD9CM|PT|614.1|Chronic salpingitis and oophoritis
C0156328|ICD9CM|AB|614.1|Chr salpingo-oophoritis
C0156329|ICD9CM|PT|614.3|Acute parametritis and pelvic cellulitis
C0156329|ICD9CM|AB|614.3|Acute parametritis
C0156332|ICD9CM|PT|614.7|Other chronic pelvic peritonitis, female
C0156332|ICD9CM|AB|614.7|Chr pelv periton NEC-fem
C0156333|ICD9CM|HT|615|Inflammatory diseases of uterus, except cervix
C0156334|ICD9CM|PT|615.0|Acute inflammatory diseases of uterus, except cervix
C0156334|ICD9CM|AB|615.0|Ac uterine inflammation
C0156335|ICD9CM|PT|615.1|Chronic inflammatory diseases of uterus, except cervix
C0156335|ICD9CM|AB|615.1|Chr uterine inflammation
C0156337|ICD9CM|PT|616.11|Vaginitis and vulvovaginitis in diseases classified elsewhere
C0156337|ICD9CM|AB|616.11|Vaginitis in oth disease
C0156338|ICD9CM|PT|616.4|Other abscess of vulva
C0156338|ICD9CM|AB|616.4|Abscess of vulva NEC
C0156339|ICD9CM|HT|616.5|Ulceration of vulva
C0156339|ICD9CM|AB|616.50|Ulceration of vulva NOS
C0156339|ICD9CM|PT|616.50|Ulceration of vulva, unspecified
C0156340|ICD9CM|PT|616.51|Ulceration of vulva in diseases classified elsewhere
C0156340|ICD9CM|AB|616.51|Vulvar ulcer in oth dis
C0156341|ICD9CM|HT|616.8|Other specified inflammatory diseases of cervix, vagina, and vulva
C0156342|ICD9CM|PT|616.9|Unspecified inflammatory disease of cervix, vagina, and vulva
C0156342|ICD9CM|HT|616|Inflammatory disease of cervix, vagina, and vulva
C0156342|ICD9CM|AB|616.9|Female gen inflam NOS
C0156344|ICD9CM|PT|617.1|Endometriosis of ovary
C0156344|ICD9CM|AB|617.1|Ovarian endometriosis
C0156345|ICD9CM|PT|617.3|Endometriosis of pelvic peritoneum
C0156345|ICD9CM|AB|617.3|Pelv perit endometriosis
C0156346|ICD9CM|PT|617.4|Endometriosis of rectovaginal septum and vagina
C0156346|ICD9CM|AB|617.4|Vaginal endometriosis
C0156347|ICD9CM|PT|617.5|Endometriosis of intestine
C0156347|ICD9CM|AB|617.5|Intestinal endometriosis
C0156348|ICD9CM|PT|617.6|Endometriosis in scar of skin
C0156348|ICD9CM|AB|617.6|Endometriosis in scar
C0156349|ICD9CM|HT|618|Genital prolapse
C0156350|ICD9CM|HT|618.0|Prolapse of vaginal walls without mention of uterine prolapse
C0156351|ICD9CM|PT|618.2|Uterovaginal prolapse, incomplete
C0156351|ICD9CM|AB|618.2|Uterovag prolaps-incompl
C0156353|ICD9CM|PT|618.4|Uterovaginal prolapse, unspecified
C0156353|ICD9CM|AB|618.4|Utervaginal prolapse NOS
C0156354|ICD9CM|PT|618.5|Prolapse of vaginal vault after hysterectomy
C0156354|ICD9CM|AB|618.5|Postop vaginal prolapse
C0156355|ICD9CM|PT|618.7|Old laceration of muscles of pelvic floor
C0156355|ICD9CM|AB|618.7|Old lacer pelvic muscle
C0156356|ICD9CM|PT|618.9|Unspecified genital prolapse
C0156356|ICD9CM|AB|618.9|Genital prolapse NOS
C0156357|ICD9CM|HT|619|Fistula involving female genital tract
C0156358|ICD9CM|PT|619.2|Genital tract-skin fistula, female
C0156358|ICD9CM|AB|619.2|Genital-skin fistul, fem
C0156361|ICD9CM|PT|620.1|Corpus luteum cyst or hematoma
C0156361|ICD9CM|AB|620.1|Corpus luteum cyst
C0156362|ICD9CM|PT|620.3|Acquired atrophy of ovary and fallopian tube
C0156362|ICD9CM|AB|620.3|Acq atrophy ovary & tube
C0156364|ICD9CM|PT|620.5|Torsion of ovary, ovarian pedicle, or fallopian tube
C0156364|ICD9CM|AB|620.5|Torsion of ovary or tube
C0156365|ICD9CM|PT|620.7|Hematoma of broad ligament
C0156365|ICD9CM|AB|620.7|Broad ligament hematoma
C0156366|ICD9CM|PT|620.8|Other noninflammatory disorders of ovary, fallopian tube, and broad ligament
C0156366|ICD9CM|AB|620.8|Noninfl dis ova/adnx NEC
C0156367|ICD9CM|PT|620.9|Unspecified noninflammatory disorder of ovary, fallopian tube, and broad ligament
C0156367|ICD9CM|HT|620|Noninflammatory disorders of ovary, fallopian tube, and broad ligament
C0156367|ICD9CM|AB|620.9|Noninfl dis ova/adnx NOS
C0156369|ICD9CM|AB|621.0|Polyp of corpus uteri
C0156369|ICD9CM|PT|621.0|Polyp of corpus uteri
C0156370|ICD9CM|PT|621.1|Chronic subinvolution of uterus
C0156370|ICD9CM|AB|621.1|Chr uterine subinvolutn
C0156371|ICD9CM|AB|621.2|Hypertrophy of uterus
C0156371|ICD9CM|PT|621.2|Hypertrophy of uterus
C0156373|ICD9CM|AB|621.6|Malposition of uterus
C0156373|ICD9CM|PT|621.6|Malposition of uterus
C0156374|ICD9CM|PT|621.7|Chronic inversion of uterus
C0156374|ICD9CM|AB|621.7|Chr inversion of uterus
C0156377|ICD9CM|HT|622|Noninflammatory disorders of cervix
C0156377|ICD9CM|PT|622.9|Unspecified noninflammatory disorder of cervix
C0156377|ICD9CM|AB|622.9|Noninflam dis cervix NOS
C0156379|ICD9CM|AB|622.3|Old laceration of cervix
C0156379|ICD9CM|PT|622.3|Old laceration of cervix
C0156380|ICD9CM|PT|622.4|Stricture and stenosis of cervix
C0156380|ICD9CM|AB|622.4|Stricture of cervix
C0156383|ICD9CM|HT|623|Noninflammatory disorders of vagina
C0156383|ICD9CM|PT|623.9|Unspecified noninflammatory disorder of vagina
C0156383|ICD9CM|AB|623.9|Noninflam dis vagina NOS
C0156384|ICD9CM|AB|623.0|Dysplasia of vagina
C0156384|ICD9CM|PT|623.0|Dysplasia of vagina
C0156385|ICD9CM|AB|623.1|Leukoplakia of vagina
C0156385|ICD9CM|PT|623.1|Leukoplakia of vagina
C0156386|ICD9CM|PT|623.2|Stricture or atresia of vagina
C0156386|ICD9CM|AB|623.2|Stricture of vagina
C0156387|ICD9CM|AB|623.3|Tight hymenal ring
C0156387|ICD9CM|PT|623.3|Tight hymenal ring
C0156388|ICD9CM|AB|623.4|Old vaginal laceration
C0156388|ICD9CM|PT|623.4|Old vaginal laceration
C0156389|ICD9CM|AB|623.6|Vaginal hematoma
C0156389|ICD9CM|PT|623.6|Vaginal hematoma
C0156390|ICD9CM|AB|623.7|Polyp of vagina
C0156390|ICD9CM|PT|623.7|Polyp of vagina
C0156393|ICD9CM|AB|624.1|Atrophy of vulva
C0156393|ICD9CM|PT|624.1|Atrophy of vulva
C0156394|ICD9CM|AB|624.2|Hypertrophy of clitoris
C0156394|ICD9CM|PT|624.2|Hypertrophy of clitoris
C0156397|ICD9CM|AB|624.5|Hematoma of vulva
C0156397|ICD9CM|PT|624.5|Hematoma of vulva
C0156398|ICD9CM|AB|624.6|Polyp of labia and vulva
C0156398|ICD9CM|PT|624.6|Polyp of labia and vulva
C0156399|ICD9CM|PT|624.8|Other specified noninflammatory disorders of vulva and perineum
C0156399|ICD9CM|AB|624.8|Noninflam dis vulva NEC
C0156400|ICD9CM|PT|624.9|Unspecified noninflammatory disorder of vulva and perineum
C0156400|ICD9CM|HT|624|Noninflammatory disorders of vulva and perineum
C0156400|ICD9CM|AB|624.9|Noninflam dis vulva NOS
C0156401|ICD9CM|HT|625|Pain and other symptoms associated with female genital organs
C0156402|ICD9CM|PT|625.8|Other specified symptoms associated with female genital organs
C0156402|ICD9CM|AB|625.8|Fem genital symptoms NEC
C0156403|ICD9CM|AB|626.3|Pubertal menorrhagia
C0156403|ICD9CM|PT|626.3|Puberty bleeding
C0156404|ICD9CM|AB|626.4|Irregular menstruation
C0156404|ICD9CM|PT|626.4|Irregular menstrual cycle
C0156405|ICD9CM|AB|626.5|Ovulation bleeding
C0156405|ICD9CM|PT|626.5|Ovulation bleeding
C0156406|ICD9CM|AB|626.7|Postcoital bleeding
C0156406|ICD9CM|PT|626.7|Postcoital bleeding
C0156407|ICD9CM|HT|627|Menopausal and postmenopausal disorders
C0156407|ICD9CM|PT|627.9|Unspecified menopausal and postmenopausal disorder
C0156407|ICD9CM|AB|627.9|Menopausal disorder NOS
C0156408|ICD9CM|PT|627.0|Premenopausal menorrhagia
C0156408|ICD9CM|AB|627.0|Premenopause menorrhagia
C0156409|ICD9CM|PT|627.3|Postmenopausal atrophic vaginitis
C0156409|ICD9CM|AB|627.3|Atrophic vaginitis
C0156411|ICD9CM|PT|627.8|Other specified menopausal and postmenopausal disorders
C0156411|ICD9CM|AB|627.8|Menopausal disorder NEC
C0156414|ICD9CM|PT|628.1|Infertility, female, of pituitary-hypothalamic origin
C0156414|ICD9CM|AB|628.1|Infertil-pituitary orig
C0156415|ICD9CM|PT|628.2|Infertility, female, of tubal origin
C0156415|ICD9CM|AB|628.2|Infertility-tubal origin
C0156416|ICD9CM|PT|628.3|Infertility, female, of uterine origin
C0156416|ICD9CM|AB|628.3|Infertility-uterine orig
C0156417|ICD9CM|PT|628.4|Infertility, female, of cervical or vaginal origin
C0156417|ICD9CM|AB|628.4|Infertil-cervical orig
C0156418|ICD9CM|HT|629|Other disorders of female genital organs
C0156420|ICD9CM|PT|629.1|Hydrocele, canal of nuck
C0156420|ICD9CM|AB|629.1|Hydrocele canal nuck-fem
C0156421|ICD9CM|HT|629.8|Other specified disorders of female genital organs
C0156421|ICD9CM|PT|629.89|Other specified disorders of female genital organs
C0156421|ICD9CM|AB|629.89|Female genital disor NEC
C0156422|ICD9CM|PT|631.8|Other abnormal products of conception
C0156422|ICD9CM|HT|631|Other abnormal product of conception
C0156422|ICD9CM|AB|631.8|Oth abn prod conception
C0156424|ICD9CM|PT|634.00|Spontaneous abortion, complicated by genital tract and pelvic infection, unspecified
C0156424|ICD9CM|HT|634.0|Spontaneous abortion complicated by genital tract and pelvic infection
C0156424|ICD9CM|AB|634.00|Spon abor w pel inf-unsp
C0156425|ICD9CM|PT|634.01|Spontaneous abortion, complicated by genital tract and pelvic infection, incomplete
C0156425|ICD9CM|AB|634.01|Spon abor w pelv inf-inc
C0156426|ICD9CM|PT|634.02|Spontaneous abortion, complicated by genital tract and pelvic infection, complete
C0156426|ICD9CM|AB|634.02|Spon abor w pel inf-comp
C0156427|ICD9CM|HT|634.1|Spontaneous abortion complicated by delayed or excessive hemorrhage
C0156428|ICD9CM|PT|634.10|Spontaneous abortion, complicated by delayed or excessive hemorrhage, unspecified
C0156428|ICD9CM|AB|634.10|Spon abort w hemorr-unsp
C0156429|ICD9CM|PT|634.11|Spontaneous abortion, complicated by delayed or excessive hemorrhage, incomplete
C0156429|ICD9CM|AB|634.11|Spon abort w hemorr-inc
C0156430|ICD9CM|PT|634.12|Spontaneous abortion, complicated by delayed or excessive hemorrhage, complete
C0156430|ICD9CM|AB|634.12|Spon abort w hemorr-comp
C0156433|ICD9CM|PT|634.21|Spontaneous abortion, complicated by damage to pelvic organs or tissues, incomplete
C0156433|ICD9CM|AB|634.21|Spon ab w pelv damag-inc
C0156434|ICD9CM|PT|634.22|Spontaneous abortion, complicated by damage to pelvic organs or tissues, complete
C0156434|ICD9CM|AB|634.22|Spon ab w pel damag-comp
C0156435|ICD9CM|HT|634.3|Spontaneous abortion complicated by renal failure
C0156436|ICD9CM|PT|634.30|Spontaneous abortion, complicated by renal failure, unspecified
C0156436|ICD9CM|AB|634.30|Spon ab w ren fail-unsp
C0156439|ICD9CM|HT|634.4|Spontaneous abortion complicated by metabolic disorder
C0156439|ICD9CM|PT|634.40|Spontaneous abortion, complicated by metabolic disorder, unspecified
C0156439|ICD9CM|AB|634.40|Spon ab w metab dis-unsp
C0156442|ICD9CM|PT|634.42|Spontaneous abortion, complicated by metabolic disorder, complete
C0156442|ICD9CM|AB|634.42|Spon ab w metab dis-comp
C0156443|ICD9CM|HT|634.5|Spontaneous abortion complicated by shock
C0156444|ICD9CM|PT|634.50|Spontaneous abortion, complicated by shock, unspecified
C0156444|ICD9CM|AB|634.50|Spon abort w shock-unsp
C0156445|ICD9CM|PT|634.51|Spontaneous abortion, complicated by shock, incomplete
C0156445|ICD9CM|AB|634.51|Spon abort w shock-inc
C0156447|ICD9CM|HT|634.6|Spontaneous abortion complicated by embolism
C0156448|ICD9CM|PT|634.60|Spontaneous abortion, complicated by embolism, unspecified
C0156448|ICD9CM|AB|634.60|Spon abort w embol-unsp
C0156452|ICD9CM|PT|634.70|Spontaneous abortion, with other specified complications, unspecified
C0156452|ICD9CM|HT|634.7|Spontaneous abortion with other specified complications
C0156452|ICD9CM|AB|634.70|Spon ab w compl NEC-unsp
C0156453|ICD9CM|PT|634.71|Spontaneous abortion, with other specified complications, incomplete
C0156453|ICD9CM|AB|634.71|Spon ab w compl NEC-inc
C0156454|ICD9CM|PT|634.72|Spontaneous abortion, with other specified complications, complete
C0156454|ICD9CM|AB|634.72|Spon ab w compl NEC-comp
C0156456|ICD9CM|HT|634.8|Spontaneous abortion with unspecified complication
C0156456|ICD9CM|PT|634.80|Spontaneous abortion, with unspecified complication, unspecified
C0156456|ICD9CM|AB|634.80|Spon ab w compl NOS-unsp
C0156457|ICD9CM|PT|634.81|Spontaneous abortion, with unspecified complication, incomplete
C0156457|ICD9CM|AB|634.81|Spon ab w compl NOS-inc
C0156458|ICD9CM|PT|634.82|Spontaneous abortion, with unspecified complication, complete
C0156458|ICD9CM|AB|634.82|Spon ab w compl NOS-comp
C0156459|ICD9CM|PT|634.90|Spontaneous abortion, without mention of complication, unspecified
C0156459|ICD9CM|HT|634.9|Spontaneous abortion without mention of complication
C0156459|ICD9CM|AB|634.90|Spon abort uncompl-unsp
C0156461|ICD9CM|PT|634.92|Spontaneous abortion, without mention of complication, complete
C0156461|ICD9CM|AB|634.92|Spon abort uncompl-comp
C0156464|ICD9CM|PT|635.00|Legally induced abortion, complicated by genital tract and pelvic infection, unspecified
C0156464|ICD9CM|HT|635.0|Legally induced abortion complicated by genital tract and pelvic infection
C0156464|ICD9CM|AB|635.00|Leg abor w pelv inf-unsp
C0156465|ICD9CM|PT|635.01|Legally induced abortion, complicated by genital tract and pelvic infection, incomplete
C0156465|ICD9CM|AB|635.01|Leg abor w pelv inf-inc
C0156466|ICD9CM|PT|635.02|Legally induced abortion, complicated by genital tract and pelvic infection, complete
C0156466|ICD9CM|AB|635.02|Leg abor w pelv inf-comp
C0156469|ICD9CM|PT|635.11|Legally induced abortion, complicated by delayed or excessive hemorrhage, incomplete
C0156469|ICD9CM|AB|635.11|Legal abort w hemorr-inc
C0156470|ICD9CM|PT|635.12|Legally induced abortion, complicated by delayed or excessive hemorrhage, complete
C0156470|ICD9CM|AB|635.12|Legal abor w hemorr-comp
C0156472|ICD9CM|HT|635.2|Legally induced abortion complicated by damage to pelvic organs or tissues
C0156472|ICD9CM|PT|635.20|Legally induced abortion, complicated by damage to pelvic organs or tissues, unspecified
C0156472|ICD9CM|AB|635.20|Leg ab w pelv damag-unsp
C0156473|ICD9CM|PT|635.21|Legally induced abortion, complicated by damage to pelvic organs or tissues, incomplete
C0156473|ICD9CM|AB|635.21|Leg ab w pelv damag-inc
C0156474|ICD9CM|PT|635.22|Legally induced abortion, complicated by damage to pelvic organs or tissues, complete
C0156474|ICD9CM|AB|635.22|Leg ab w pelv damag-comp
C0156477|ICD9CM|PT|635.31|Legally induced abortion, complicated by renal failure, incomplete
C0156477|ICD9CM|AB|635.31|Leg abor w ren fail-inc
C0156478|ICD9CM|PT|635.32|Legally induced abortion, complicated by renal failure, complete
C0156478|ICD9CM|AB|635.32|Leg abor w ren fail-comp
C0156481|ICD9CM|PT|635.41|Legally induced abortion, complicated by metabolic disorder, incomplete
C0156481|ICD9CM|AB|635.41|Leg ab w metab dis-inc
C0156482|ICD9CM|PT|635.42|Legally induced abortion, complicated by metabolic disorder, complete
C0156482|ICD9CM|AB|635.42|Leg ab w metab dis-comp
C0156485|ICD9CM|PT|635.51|Legally induced abortion, complicated by shock, incomplete
C0156485|ICD9CM|AB|635.51|Legal abort w shock-inc
C0156486|ICD9CM|PT|635.52|Legally induced abortion, complicated by shock, complete
C0156486|ICD9CM|AB|635.52|Legal abort w shock-comp
C0156489|ICD9CM|PT|635.61|Legally induced abortion, complicated by embolism, incomplete
C0156489|ICD9CM|AB|635.61|Legal abort w embol-inc
C0156490|ICD9CM|PT|635.62|Legally induced abortion, complicated by embolism, complete
C0156490|ICD9CM|AB|635.62|Legal abort w embol-comp
C0156492|ICD9CM|PT|635.70|Legally induced abortion, with other specified complications, unspecified
C0156492|ICD9CM|HT|635.7|Legally induced abortion with other specified complications
C0156492|ICD9CM|AB|635.70|Leg ab w compl NEC-unsp
C0156493|ICD9CM|PT|635.71|Legally induced abortion, with other specified complications, incomplete
C0156493|ICD9CM|AB|635.71|Leg ab w compl NEC-inc
C0156494|ICD9CM|PT|635.72|Legally induced abortion, with other specified complications, complete
C0156494|ICD9CM|AB|635.72|Leg ab w compl NEC-comp
C0156499|ICD9CM|PT|635.90|Legally induced abortion, without mention of complication, unspecified
C0156499|ICD9CM|HT|635.9|Legally induced abortion without mention of complication
C0156499|ICD9CM|AB|635.90|Legal abort uncompl-unsp
C0156504|ICD9CM|PT|636.00|Illegally induced abortion, complicated by genital tract and pelvic infection, unspecified
C0156504|ICD9CM|HT|636.0|Illegally induced abortion complicated by genital tract and pelvic infection
C0156504|ICD9CM|AB|636.00|Illeg ab w pelv inf-unsp
C0156505|ICD9CM|PT|636.01|Illegally induced abortion, complicated by genital tract and pelvic infection, incomplete
C0156505|ICD9CM|AB|636.01|Illeg ab w pelv inf-inc
C0156506|ICD9CM|PT|636.02|Illegally induced abortion, complicated by genital tract and pelvic infection, complete
C0156506|ICD9CM|AB|636.02|Illeg ab w pelv inf-comp
C0156509|ICD9CM|PT|636.11|Illegally induced abortion, complicated by delayed or excessive hemorrhage, incomplete
C0156509|ICD9CM|AB|636.11|Illeg ab w hemorr-inc
C0156510|ICD9CM|PT|636.12|Illegally induced abortion, complicated by delayed or excessive hemorrhage, complete
C0156510|ICD9CM|AB|636.12|Illeg ab w hemorr-comp
C0156513|ICD9CM|PT|636.21|Illegally induced abortion, complicated by damage to pelvic organs or tissues, incomplete
C0156513|ICD9CM|AB|636.21|Illeg ab w pel damag-inc
C0156514|ICD9CM|PT|636.22|Illegally induced abortion, complicated by damage to pelvic organs or tissues, complete
C0156514|ICD9CM|AB|636.22|Illeg ab w pel damg-comp
C0156517|ICD9CM|PT|636.31|Illegally induced abortion, complicated by renal failure, incomplete
C0156517|ICD9CM|AB|636.31|Illeg ab w ren fail-inc
C0156518|ICD9CM|PT|636.32|Illegally induced abortion, complicated by renal failure, complete
C0156518|ICD9CM|AB|636.32|Illeg ab w ren fail-comp
C0156521|ICD9CM|PT|636.41|Illegally induced abortion, complicated by metabolic disorder, incomplete
C0156521|ICD9CM|AB|636.41|Illeg ab w metab dis-inc
C0156522|ICD9CM|PT|636.42|Illegally induced abortion, complicated by metabolic disorder, complete
C0156522|ICD9CM|AB|636.42|Illeg ab w met dis-comp
C0156525|ICD9CM|PT|636.51|Illegally induced abortion, complicated by shock, incomplete
C0156525|ICD9CM|AB|636.51|Illeg abort w shock-inc
C0156526|ICD9CM|PT|636.52|Illegally induced abortion, complicated by shock, complete
C0156526|ICD9CM|AB|636.52|Illeg abort w shock-comp
C0156529|ICD9CM|PT|636.61|Illegally induced abortion, complicated by embolism, incomplete
C0156529|ICD9CM|AB|636.61|Illeg ab w embolism-inc
C0156530|ICD9CM|PT|636.62|Illegally induced abortion, complicated by embolism, complete
C0156530|ICD9CM|AB|636.62|Illeg ab w embolism-comp
C0156532|ICD9CM|PT|636.70|Illegally induced abortion, with other specified complications, unspecified
C0156532|ICD9CM|HT|636.7|Illegally induced abortion with other specified complications
C0156532|ICD9CM|AB|636.70|Illg ab w compl NEC-unsp
C0156533|ICD9CM|PT|636.71|Illegally induced abortion, with other specified complications, incomplete
C0156533|ICD9CM|AB|636.71|Illeg ab w compl NEC-inc
C0156534|ICD9CM|PT|636.72|Illegally induced abortion, with other specified complications, complete
C0156534|ICD9CM|AB|636.72|Illg ab w compl NEC-comp
C0156537|ICD9CM|PT|636.81|Illegally induced abortion, with unspecified complication, incomplete
C0156537|ICD9CM|AB|636.81|Illeg ab w compl NOS-inc
C0156538|ICD9CM|PT|636.82|Illegally induced abortion, with unspecified complication, complete
C0156538|ICD9CM|AB|636.82|Illg ab w compl NOS-comp
C0156541|ICD9CM|PT|636.91|Illegally induced abortion, without mention of complication, incomplete
C0156541|ICD9CM|AB|636.91|Illeg abort uncompl-inc
C0156542|ICD9CM|PT|636.92|Illegally induced abortion, without mention of complication, complete
C0156542|ICD9CM|AB|636.92|Illeg abort uncompl-comp
C0156543|ICD9CM|HT|637|Unspecified abortion
C0156545|ICD9CM|PT|637.00|Unspecified abortion, complicated by genital tract and pelvic infection, unspecified
C0156545|ICD9CM|HT|637.0|Unspecified abortion complicated by genital tract and pelvic infection
C0156545|ICD9CM|AB|637.00|Abort NOS w pel inf-unsp
C0156546|ICD9CM|PT|637.01|Unspecified abortion, complicated by genital tract and pelvic infection, incomplete
C0156546|ICD9CM|AB|637.01|Abort NOS w pel inf-inc
C0156547|ICD9CM|PT|637.02|Unspecified abortion, complicated by genital tract and pelvic infection, complete
C0156547|ICD9CM|AB|637.02|Abort NOS w pel inf-comp
C0156548|ICD9CM|HT|637.1|Unspecified abortion complicated by delayed or excessive hemorrhage
C0156548|ICD9CM|PT|637.10|Unspecified abortion, complicated by delayed or excessive hemorrhage, unspecified
C0156548|ICD9CM|AB|637.10|Abort NOS w hemorr-unsp
C0156550|ICD9CM|PT|637.11|Unspecified abortion, complicated by delayed or excessive hemorrhage, incomplete
C0156550|ICD9CM|AB|637.11|Abort NOS w hemorr-inc
C0156551|ICD9CM|PT|637.12|Unspecified abortion, complicated by delayed or excessive hemorrhage, complete
C0156551|ICD9CM|AB|637.12|Abort NOS w hemorr-comp
C0156554|ICD9CM|PT|637.21|Unspecified abortion, complicated by damage to pelvic organs or tissues, incomplete
C0156554|ICD9CM|AB|637.21|Ab NOS w pelv damag-inc
C0156555|ICD9CM|PT|637.22|Unspecified abortion, complicated by damage to pelvic organs or tissues, complete
C0156555|ICD9CM|AB|637.22|Ab NOS w pelv damag-comp
C0156556|ICD9CM|HT|637.3|Unspecified abortion complicated by renal failure
C0156556|ICD9CM|PT|637.30|Unspecified abortion, complicated by renal failure, unspecified
C0156556|ICD9CM|AB|637.30|Ab NOS w renal fail-unsp
C0156558|ICD9CM|PT|637.31|Unspecified abortion, complicated by renal failure, incomplete
C0156558|ICD9CM|AB|637.31|Ab NOS w renal fail-inc
C0156559|ICD9CM|PT|637.32|Unspecified abortion, complicated by renal failure, complete
C0156559|ICD9CM|AB|637.32|Ab NOS w renal fail-comp
C0156560|ICD9CM|HT|637.4|Unspecified abortion complicated by metabolic disorder
C0156561|ICD9CM|PT|637.40|Unspecified abortion, complicated by metabolic disorder, unspecified
C0156561|ICD9CM|AB|637.40|Ab NOS w metab dis-unsp
C0156562|ICD9CM|PT|637.41|Unspecified abortion, complicated by metabolic disorder, incomplete
C0156562|ICD9CM|AB|637.41|Ab NOS w metab dis-inc
C0156563|ICD9CM|PT|637.42|Unspecified abortion, complicated by metabolic disorder, complete
C0156563|ICD9CM|AB|637.42|Ab NOS w metab dis-comp
C0156564|ICD9CM|HT|637.5|Unspecified abortion complicated by shock
C0156564|ICD9CM|PT|637.50|Unspecified abortion, complicated by shock, unspecified
C0156564|ICD9CM|AB|637.50|Abort NOS w shock-unsp
C0156566|ICD9CM|PT|637.51|Unspecified abortion, complicated by shock, incomplete
C0156566|ICD9CM|AB|637.51|Abort NOS w shock-inc
C0156567|ICD9CM|PT|637.52|Unspecified abortion, complicated by shock, complete
C0156567|ICD9CM|AB|637.52|Abort NOS w shock-comp
C0156568|ICD9CM|HT|637.6|Unspecified abortion complicated by embolism
C0156568|ICD9CM|PT|637.60|Unspecified abortion, complicated by embolism, unspecified
C0156568|ICD9CM|AB|637.60|Ab NOS w embolism-unsp
C0156570|ICD9CM|PT|637.61|Unspecified abortion, complicated by embolism, incomplete
C0156570|ICD9CM|AB|637.61|Ab NOS w embolism-inc
C0156571|ICD9CM|PT|637.62|Unspecified abortion, complicated by embolism, complete
C0156571|ICD9CM|AB|637.62|Ab NOS w embolism-comp
C0156572|ICD9CM|HT|637.7|Unspecified abortion with other specified complications
C0156573|ICD9CM|PT|637.70|Unspecified abortion, with other specified complications, unspecified
C0156573|ICD9CM|AB|637.70|Ab NOS w compl NEC-unsp
C0156574|ICD9CM|PT|637.71|Unspecified abortion, with other specified complications, incomplete
C0156574|ICD9CM|AB|637.71|Ab NOS w compl NEC-inc
C0156575|ICD9CM|PT|637.72|Unspecified abortion, with other specified complications, complete
C0156575|ICD9CM|AB|637.72|Ab NOS w compl NEC-comp
C0156578|ICD9CM|PT|637.81|Unspecified abortion, with unspecified complication, incomplete
C0156578|ICD9CM|AB|637.81|Ab NOS w compl NOS-inc
C0156579|ICD9CM|PT|637.82|Unspecified abortion, with unspecified complication, complete
C0156579|ICD9CM|AB|637.82|Ab NOS w compl NOS-comp
C0156580|ICD9CM|PT|637.90|Unspecified abortion, without mention of complication, unspecified
C0156580|ICD9CM|HT|637.9|Unspecified abortion without mention of complication
C0156580|ICD9CM|AB|637.90|Ab NOS uncomplicat-unsp
C0156581|ICD9CM|PT|637.91|Unspecified abortion, without mention of complication, incomplete
C0156581|ICD9CM|AB|637.91|Ab NOS uncomplicat-inc
C0156582|ICD9CM|PT|637.92|Unspecified abortion, without mention of complication, complete
C0156582|ICD9CM|AB|637.92|Ab NOS uncomplicat-comp
C0156584|ICD9CM|PT|638.0|Failed attempted abortion complicated by genital tract and pelvic infection
C0156584|ICD9CM|AB|638.0|Attem abort w pelvic inf
C0156585|ICD9CM|PT|638.1|Failed attempted abortion complicated by delayed or excessive hemorrhage
C0156585|ICD9CM|AB|638.1|Attem abort w hemorrhage
C0156587|ICD9CM|PT|638.3|Failed attempted abortion complicated by renal failure
C0156587|ICD9CM|AB|638.3|Attem abort w renal fail
C0156588|ICD9CM|PT|638.4|Failed attempted abortion complicated by metabolic disorder
C0156588|ICD9CM|AB|638.4|Attem abor w metabol dis
C0156589|ICD9CM|PT|638.5|Failed attempted abortion complicated by shock
C0156589|ICD9CM|AB|638.5|Attem abortion w shock
C0156590|ICD9CM|PT|638.6|Failed attempted abortion complicated by embolism
C0156590|ICD9CM|AB|638.6|Attemp abort w embolism
C0156591|ICD9CM|PT|638.7|Failed attempted abortion with other specified complications
C0156591|ICD9CM|AB|638.7|Attemp abort w compl NEC
C0156592|ICD9CM|PT|638.8|Failed attempted abortion with unspecified complication
C0156592|ICD9CM|AB|638.8|Attemp abort w compl NOS
C0156602|ICD9CM|PT|639.8|Other specified complications following abortion or ectopic and molar pregnancy
C0156602|ICD9CM|AB|639.8|Postabortion compl NEC
C0156604|ICD9CM|HT|640|Hemorrhage in early pregnancy
C0156604|ICD9CM|HT|640.9|Unspecified hemorrhage in early pregnancy
C0156605|ICD9CM|PT|640.00|Threatened abortion, unspecified as to episode of care or not applicable
C0156605|ICD9CM|AB|640.00|Threatened abort-unspec
C0156606|ICD9CM|PT|640.01|Threatened abortion, delivered, with or without mention of antepartum condition
C0156606|ICD9CM|AB|640.01|Threatened abort-deliver
C0156608|ICD9CM|HT|640.8|Other specified hemorrhage in early pregnancy
C0156609|ICD9CM|PT|640.80|Other specified hemorrhage in early pregnancy, unspecified as to episode of care or not applicable
C0156609|ICD9CM|AB|640.80|Hem early preg NEC-unsp
C0156610|ICD9CM|PT|640.81|Other specified hemorrhage in early pregnancy, delivered, with or without mention of antepartum condition
C0156610|ICD9CM|AB|640.81|Hem early preg NEC-deliv
C0156613|ICD9CM|PT|640.90|Unspecified hemorrhage in early pregnancy, unspecified as to episode of care or not applicable
C0156613|ICD9CM|AB|640.90|Hemorr early preg-unspec
C0156614|ICD9CM|PT|640.91|Unspecified hemorrhage in early pregnancy, delivered, with or without mention of antepartum condition
C0156614|ICD9CM|AB|640.91|Hem early preg-delivered
C0156616|ICD9CM|HT|641|Antepartum hemorrhage, abruptio placentae, and placenta previa
C0156617|ICD9CM|HT|641.0|Placenta previa without hemorrhage
C0156618|ICD9CM|PT|641.00|Placenta previa without hemorrhage, unspecified as to episode of care or not applicable
C0156618|ICD9CM|AB|641.00|Placenta previa-unspec
C0156619|ICD9CM|PT|641.01|Placenta previa without hemorrhage, delivered, with or without mention of antepartum condition
C0156619|ICD9CM|AB|641.01|Placenta previa-deliver
C0156620|ICD9CM|PT|641.03|Placenta previa without hemorrhage, antepartum condition or complication
C0156620|ICD9CM|AB|641.03|Placenta previa-antepart
C0156621|ICD9CM|HT|641.1|Hemorrhage from placenta previa
C0156621|ICD9CM|PT|641.10|Hemorrhage from placenta previa, unspecified as to episode of care or not applicable
C0156621|ICD9CM|AB|641.10|Placenta prev hem-unspec
C0156623|ICD9CM|PT|641.11|Hemorrhage from placenta previa, delivered, with or without mention of antepartum condition
C0156623|ICD9CM|AB|641.11|Placenta prev hem-deliv
C0156624|ICD9CM|PT|641.13|Hemorrhage from placenta previa, antepartum condition or complication
C0156624|ICD9CM|AB|641.13|Placen prev hem-antepart
C0156626|ICD9CM|PT|641.21|Premature separation of placenta, delivered, with or without mention of antepartum condition
C0156626|ICD9CM|AB|641.21|Prem separ placen-deliv
C0156627|ICD9CM|PT|641.23|Premature separation of placenta, antepartum condition or complication
C0156627|ICD9CM|AB|641.23|Prem separ plac-antepart
C0156629|ICD9CM|PT|641.30|Antepartum hemorrhage associated with coagulation defects, unspecified as to episode of care or not applicable
C0156629|ICD9CM|AB|641.30|Coag def hemorr-unspec
C0156630|ICD9CM|PT|641.31|Antepartum hemorrhage associated with coagulation defects, delivered, with or without mention of antepartum condition
C0156630|ICD9CM|AB|641.31|Coag def hemorr-deliver
C0156631|ICD9CM|HT|641.3|Antepartum hemorrhage associated with coagulation defects
C0156631|ICD9CM|PT|641.33|Antepartum hemorrhage associated with coagulation defects, antepartum condition or complication
C0156631|ICD9CM|AB|641.33|Coag def hemorr-antepart
C0156633|ICD9CM|PT|641.80|Other antepartum hemorrhage, unspecified as to episode of care or not applicable
C0156633|ICD9CM|AB|641.80|Antepart hem NEC-unspec
C0156634|ICD9CM|PT|641.81|Other antepartum hemorrhage, delivered, with or without mention of antepartum condition
C0156634|ICD9CM|AB|641.81|Antepartum hem NEC-deliv
C0156635|ICD9CM|HT|641.8|Other antepartum hemorrhage
C0156635|ICD9CM|PT|641.83|Other antepartum hemorrhage, antepartum condition or complication
C0156635|ICD9CM|AB|641.83|Antepart hem NEC-antepar
C0156637|ICD9CM|PT|641.90|Unspecified antepartum hemorrhage, unspecified as to episode of care or not applicable
C0156637|ICD9CM|AB|641.90|Antepart hem NOS-unspec
C0156638|ICD9CM|PT|641.91|Unspecified antepartum hemorrhage, delivered, with or without mention of antepartum condition
C0156638|ICD9CM|AB|641.91|Antepartum hem NOS-deliv
C0156642|ICD9CM|PT|642.00|Benign essential hypertension complicating pregnancy, childbirth, and the puerperium, unspecified as to episode of care or not applicable
C0156642|ICD9CM|AB|642.00|Essen hyperten preg-unsp
C0156643|ICD9CM|PT|642.01|Benign essential hypertension complicating pregnancy, childbirth, and the puerperium, delivered, with or without mention of antepartum condition
C0156643|ICD9CM|AB|642.01|Essen hyperten-delivered
C0156644|ICD9CM|PT|642.02|Benign essential hypertension, complicating pregnancy, childbirth, and the puerperium, delivered, with mention of postpartum complication
C0156644|ICD9CM|AB|642.02|Essen hyperten-del w p/p
C0156645|ICD9CM|PT|642.03|Benign essential hypertension complicating pregnancy, childbirth, and the puerperium, antepartum condition or complication
C0156645|ICD9CM|AB|642.03|Essen hyperten-antepart
C0156646|ICD9CM|PT|642.04|Benign essential hypertension complicating pregnancy, childbirth, and the puerperium, postpartum condition or complication
C0156646|ICD9CM|AB|642.04|Essen hyperten-postpart
C0156647|ICD9CM|HT|642.1|Hypertension secondary to renal disease, complicating pregnancy, childbirth, and the puerperium
C0156648|ICD9CM|PT|642.10|Hypertension secondary to renal disease, complicating pregnancy, childbirth, and the puerperium, unspecified as to episode of care or not applicable
C0156648|ICD9CM|AB|642.10|Renal hyperten preg-unsp
C0156649|ICD9CM|PT|642.11|Hypertension secondary to renal disease, complicating pregnancy, childbirth, and the puerperium, delivered, with or without mention of antepartum condition
C0156649|ICD9CM|AB|642.11|Renal hyperten pg-deliv
C0156650|ICD9CM|PT|642.12|Hypertension secondary to renal disease, complicating pregnancy, childbirth, and the puerperium, delivered, with mention of postpartum complication
C0156650|ICD9CM|AB|642.12|Renal hyperten-del p/p
C0156651|ICD9CM|PT|642.13|Hypertension secondary to renal disease, complicating pregnancy, childbirth, and the puerperium, antepartum condition or complication
C0156651|ICD9CM|AB|642.13|Renal hyperten-antepart
C0156652|ICD9CM|PT|642.14|Hypertension secondary to renal disease, complicating pregnancy, childbirth, and the puerperium, postpartum condition or complication
C0156652|ICD9CM|AB|642.14|Renal hyperten-postpart
C0156653|ICD9CM|HT|642.2|Other pre-existing hypertension complicating pregnancy, childbirth, and the puerperium
C0156654|ICD9CM|PT|642.20|Other pre-existing hypertension complicating pregnancy, childbirth, and the puerperium, unspecified as to episode of care or not applicable
C0156654|ICD9CM|AB|642.20|Old hyperten preg-unspec
C0156655|ICD9CM|PT|642.21|Other pre-existing hypertension, complicating pregnancy, childbirth, and the puerperium, delivered, with or without mention of antepartum condition
C0156655|ICD9CM|AB|642.21|Old hyperten NEC-deliver
C0156656|ICD9CM|PT|642.22|Other pre-existing hypertension, complicating pregnancy, childbirth, and the puerperium, delivered, with mention of postpartum complication
C0156656|ICD9CM|AB|642.22|Old hyperten-deliv w p/p
C0156657|ICD9CM|PT|642.23|Other pre-existing hypertension, complicating pregnancy, childbirth, and the puerperium, antepartum condition or complication
C0156657|ICD9CM|AB|642.23|Old hyperten NEC-antepar
C0156658|ICD9CM|PT|642.24|Other pre-existing hypertension,complicating pregnancy, childbirth, and the puerperium, , postpartum condition or complication
C0156658|ICD9CM|AB|642.24|Old hyperten NEC-postpar
C0156659|ICD9CM|PT|642.30|Transient hypertension of pregnancy, unspecified as to episode of care or not applicable
C0156659|ICD9CM|AB|642.30|Trans hyperten preg-unsp
C0156660|ICD9CM|PT|642.31|Transient hypertension of pregnancy, delivered , with or without mention of antepartum condition
C0156660|ICD9CM|AB|642.31|Trans hyperten-delivered
C0156661|ICD9CM|PT|642.32|Transient hypertension of pregnancy, delivered, with mention of postpartum complication
C0156661|ICD9CM|AB|642.32|Trans hyperten-del w p/p
C0156662|ICD9CM|PT|642.33|Transient hypertension of pregnancy, antepartum condition or complication
C0156662|ICD9CM|AB|642.33|Trans hyperten-antepart
C0156663|ICD9CM|PT|642.34|Transient hypertension of pregnancy, postpartum condition or complication
C0156663|ICD9CM|AB|642.34|Trans hyperten-postpart
C0156664|ICD9CM|PT|642.40|Mild or unspecified pre-eclampsia, unspecified as to episode of care or not applicable
C0156664|ICD9CM|AB|642.40|Mild/NOS preeclamp-unsp
C0156665|ICD9CM|PT|642.41|Mild or unspecified pre-eclampsia, delivered, with or without mention of antepartum condition
C0156665|ICD9CM|AB|642.41|Mild/NOS preeclamp-deliv
C0156666|ICD9CM|PT|642.42|Mild or unspecified pre-eclampsia, delivered, with mention of postpartum complication
C0156666|ICD9CM|AB|642.42|Mild preeclamp-del w p/p
C0156667|ICD9CM|PT|642.43|Mild or unspecified pre-eclampsia, antepartum condition or complication
C0156667|ICD9CM|AB|642.43|Mild/NOS preeclamp-antep
C0156668|ICD9CM|PT|642.44|Mild or unspecified pre-eclampsia, postpartum condition or complication
C0156668|ICD9CM|AB|642.44|Mild/NOS preeclamp-p/p
C0156669|ICD9CM|PT|642.50|Severe pre-eclampsia, unspecified as to episode of care or not applicable
C0156669|ICD9CM|AB|642.50|Severe preeclamp-unspec
C0156670|ICD9CM|PT|642.51|Severe pre-eclampsia, delivered, with or without mention of antepartum condition
C0156670|ICD9CM|AB|642.51|Severe preeclamp-deliver
C0156671|ICD9CM|PT|642.52|Severe pre-eclampsia, delivered, with mention of postpartum complication
C0156671|ICD9CM|AB|642.52|Sev preeclamp-del w p/p
C0156672|ICD9CM|PT|642.53|Severe pre-eclampsia, antepartum condition or complication
C0156672|ICD9CM|AB|642.53|Sev preeclamp-antepartum
C0156673|ICD9CM|PT|642.54|Severe pre-eclampsia, postpartum condition or complication
C0156673|ICD9CM|AB|642.54|Sev preeclamp-postpartum
C0156674|ICD9CM|PT|642.60|Eclampsia, unspecified as to episode of care or not applicable
C0156674|ICD9CM|AB|642.60|Eclampsia-unspecified
C0156675|ICD9CM|PT|642.61|Eclampsia, delivered, with or without mention of antepartum condition
C0156675|ICD9CM|AB|642.61|Eclampsia-delivered
C0156676|ICD9CM|PT|642.62|Eclampsia, delivered, with mention of postpartum complication
C0156676|ICD9CM|AB|642.62|Eclampsia-deliv w p/p
C0156677|ICD9CM|AB|642.63|Eclampsia-antepartum
C0156677|ICD9CM|PT|642.63|Eclampsia, antepartum condition or complication
C0156678|ICD9CM|AB|642.64|Eclampsia-postpartum
C0156678|ICD9CM|PT|642.64|Eclampsia, postpartum condition or complication
C0156679|ICD9CM|HT|642.7|Pre-eclampsia or eclampsia superimposed on pre-existing hypertension
C0156680|ICD9CM|PT|642.70|Pre-eclampsia or eclampsia superimposed on pre-existing hypertension, unspecified as to episode of care or not applicable
C0156680|ICD9CM|AB|642.70|Tox w old hyperten-unsp
C0156681|ICD9CM|PT|642.71|Pre-eclampsia or eclampsia superimposed on pre-existing hypertension, delivered, with or without mention of antepartum condition
C0156681|ICD9CM|AB|642.71|Tox w old hyperten-deliv
C0156682|ICD9CM|PT|642.72|Pre-eclampsia or eclampsia superimposed on pre-existing hypertension, delivered, with mention of postpartum complication
C0156682|ICD9CM|AB|642.72|Tox w old hyp-del w p/p
C0156683|ICD9CM|PT|642.73|Pre-eclampsia or eclampsia superimposed on pre-existing hypertension, antepartum condition or complication
C0156683|ICD9CM|AB|642.73|Tox w old hyper-antepart
C0156684|ICD9CM|PT|642.74|Pre-eclampsia or eclampsia superimposed on pre-existing hypertension, postpartum condition or complication
C0156684|ICD9CM|AB|642.74|Tox w old hyper-postpart
C0156686|ICD9CM|PT|642.90|Unspecified hypertension complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C0156686|ICD9CM|AB|642.90|Hyperten preg NOS-unspec
C0156687|ICD9CM|PT|642.91|Unspecified hypertension complicating pregnancy, childbirth, or the puerperium, delivered, with or without mention of antepartum condition
C0156687|ICD9CM|AB|642.91|Hypertens NOS-delivered
C0156688|ICD9CM|PT|642.92|Unspecified hypertension complicating pregnancy, childbirth, or the puerperium, delivered, with mention of postpartum complication
C0156688|ICD9CM|AB|642.92|Hypertens NOS-del w p/p
C0156689|ICD9CM|PT|642.93|Unspecified hypertension complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C0156689|ICD9CM|AB|642.93|Hypertens NOS-antepartum
C0156690|ICD9CM|PT|642.94|Unspecified hypertension complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication
C0156690|ICD9CM|AB|642.94|Hypertens NOS-postpartum
C0156692|ICD9CM|PT|643.00|Mild hyperemesis gravidarum, unspecified as to episode of care or not applicable
C0156692|ICD9CM|AB|643.00|Mild hyperem grav-unspec
C0156693|ICD9CM|PT|643.01|Mild hyperemesis gravidarum, delivered, with or without mention of antepartum condition
C0156693|ICD9CM|AB|643.01|Mild hyperem grav-deliv
C0156694|ICD9CM|PT|643.03|Mild hyperemesis gravidarum, antepartum condition or complication
C0156694|ICD9CM|AB|643.03|Mild hyperemesis-antepar
C0156696|ICD9CM|PT|643.10|Hyperemesis gravidarum with metabolic disturbance, unspecified as to episode of care or not applicable
C0156696|ICD9CM|AB|643.10|Hyperem w metab dis-unsp
C0156697|ICD9CM|PT|643.11|Hyperemesis gravidarum with metabolic disturbance, delivered, with or without mention of antepartum condition
C0156697|ICD9CM|AB|643.11|Hyperem w metab dis-del
C0156698|ICD9CM|PT|643.13|Hyperemesis gravidarum with metabolic disturbance, antepartum condition or complication
C0156698|ICD9CM|AB|643.13|Hyperem w metab-antepart
C0156699|ICD9CM|HT|643.2|Late vomiting of pregnancy
C0156700|ICD9CM|PT|643.20|Late vomiting of pregnancy, unspecified as to episode of care or not applicable
C0156700|ICD9CM|AB|643.20|Late vomit of preg-unsp
C0156701|ICD9CM|PT|643.21|Late vomiting of pregnancy, delivered, with or without mention of antepartum condition
C0156701|ICD9CM|AB|643.21|Late vomit of preg-deliv
C0156702|ICD9CM|PT|643.23|Late vomiting of pregnancy, antepartum condition or complication
C0156702|ICD9CM|AB|643.23|Late vomit preg-antepart
C0156703|ICD9CM|HT|643.8|Other vomiting complicating pregnancy
C0156704|ICD9CM|PT|643.80|Other vomiting complicating pregnancy, unspecified as to episode of care or not applicable
C0156704|ICD9CM|AB|643.80|Vomit compl preg-unspec
C0156705|ICD9CM|PT|643.81|Other vomiting complicating pregnancy, delivered, with or without mention of antepartum condition
C0156705|ICD9CM|AB|643.81|Vomit compl preg-deliver
C0156706|ICD9CM|PT|643.83|Other vomiting complicating pregnancy, antepartum condition or complication
C0156706|ICD9CM|AB|643.83|Vomit compl preg-antepar
C0156708|ICD9CM|PT|643.90|Unspecified vomiting of pregnancy, unspecified as to episode of care or not applicable
C0156708|ICD9CM|AB|643.90|Vomit of preg NOS-unspec
C0156709|ICD9CM|PT|643.91|Unspecified vomiting of pregnancy, delivered, with or without mention of antepartum condition
C0156709|ICD9CM|AB|643.91|Vomit of preg NOS-deliv
C0156710|ICD9CM|PT|643.93|Unspecified vomiting of pregnancy, antepartum condition or complication
C0156710|ICD9CM|AB|643.93|Vomit of pg NOS-antepart
C0156711|ICD9CM|HT|644|Early or threatened labor
C0156713|ICD9CM|PT|644.00|Threatened premature labor, unspecified as to episode of care or not applicable
C0156713|ICD9CM|AB|644.00|Threat prem labor-unspec
C0156714|ICD9CM|PT|644.03|Threatened premature labor, antepartum condition or complication
C0156714|ICD9CM|AB|644.03|Thrt prem labor-antepart
C0156716|ICD9CM|PT|644.10|Other threatened labor, unspecified as to episode of care or not applicable
C0156716|ICD9CM|AB|644.10|Threat labor NEC-unspec
C0156717|ICD9CM|PT|644.13|Other threatened labor, antepartum condition or complication
C0156717|ICD9CM|AB|644.13|Threat labor NEC-antepar
C0156718|ICD9CM|PT|644.20|Early onset of delivery, unspecified as to episode of care or not applicable
C0156718|ICD9CM|AB|644.20|Early onset deliv-unspec
C0156719|ICD9CM|PT|644.21|Early onset of delivery, delivered, with or without mention of antepartum condition
C0156719|ICD9CM|AB|644.21|Early onset delivery-del
C0156724|ICD9CM|HT|646.0|Papyraceous fetus
C0156725|ICD9CM|PT|646.00|Papyraceous fetus, unspecified as to episode of care or not applicable
C0156725|ICD9CM|AB|646.00|Papyraceous fetus-unspec
C0156726|ICD9CM|PT|646.01|Papyraceous fetus, delivered, with or without mention of antepartum condition
C0156726|ICD9CM|AB|646.01|Papyraceous fetus-deliv
C0156727|ICD9CM|PT|646.03|Papyraceous fetus, antepartum condition or complication
C0156727|ICD9CM|AB|646.03|Papyraceous fet-antepar
C0156728|ICD9CM|HT|646.1|Edema or excessive weight gain in pregnancy, without mention of hypertension
C0156729|ICD9CM|PT|646.10|Edema or excessive weight gain in pregnancy, without mention of hypertension, unspecified as to episode of care or not applicable
C0156729|ICD9CM|AB|646.10|Edema in preg-unspec
C0156730|ICD9CM|PT|646.11|Edema or excessive weight gain in pregnancy, without mention of hypertension, delivered, with or without mention of antepartum complication
C0156730|ICD9CM|AB|646.11|Edema in preg-delivered
C0156733|ICD9CM|PT|646.14|Edema or excessive weight gain in pregnancy, without mention of hypertension, postpartum condition or complication
C0156733|ICD9CM|AB|646.14|Edema in preg-postpartum
C0156736|ICD9CM|PT|646.21|Unspecified renal disease in pregnancy, without mention of hypertension, delivered, with or without mention of antepartum condition
C0156736|ICD9CM|AB|646.21|Renal dis NOS-delivered
C0156737|ICD9CM|PT|646.22|Unspecified renal disease in pregnancy, without mention of hypertension, delivered, with mention of postpartum complication
C0156737|ICD9CM|AB|646.22|Renal dis NOS-del w p/p
C0156738|ICD9CM|PT|646.23|Unspecified renal disease in pregnancy, without mention of hypertension, antepartum condition or complication
C0156738|ICD9CM|PT|646.20|Unspecified renal disease in pregnancy, without mention of hypertension, unspecified as to episode of care or not applicable
C0156738|ICD9CM|AB|646.23|Renal dis NOS-antepartum
C0156738|ICD9CM|AB|646.20|Renal dis preg NOS-unsp
C0156739|ICD9CM|PT|646.24|Unspecified renal disease in pregnancy, without mention of hypertension, postpartum condition or complication
C0156739|ICD9CM|AB|646.24|Renal dis NOS-postpartum
C0156741|ICD9CM|PT|646.30|Recurrent pregnancy loss, unspecified as to episode of care or not applicable
C0156741|ICD9CM|AB|646.30|Recur preg loss-unspec
C0156742|ICD9CM|PT|646.31|Recurrent pregnancy loss, delivered, with or without mention of antepartum condition
C0156742|ICD9CM|AB|646.31|Recurnt preg loss-deliv
C0156743|ICD9CM|PT|646.33|Recurrent pregnancy loss, antepartum condition or complication
C0156743|ICD9CM|AB|646.33|Recurnt preg loss-antep
C0156745|ICD9CM|PT|646.40|Peripheral neuritis in pregnancy, unspecified as to episode of care or not applicable
C0156745|ICD9CM|AB|646.40|Neuritis of preg-unspec
C0156746|ICD9CM|PT|646.41|Peripheral neuritis in pregnancy, delivered, with or without mention of antepartum condition
C0156746|ICD9CM|AB|646.41|Neuritis-delivered
C0156747|ICD9CM|PT|646.42|Peripheral neuritis in pregnancy, delivered, with mention of postpartum complication
C0156747|ICD9CM|AB|646.42|Neuritis-delivered w p/p
C0156749|ICD9CM|PT|646.44|Peripheral neuritis in pregnancy, postpartum condition or complication
C0156749|ICD9CM|AB|646.44|Neuritis of preg-postpar
C0156750|ICD9CM|HT|646.5|Asymptomatic bacteriuria in pregnancy
C0156750|ICD9CM|PT|646.53|Asymptomatic bacteriuria in pregnancy, antepartum condition or complication
C0156750|ICD9CM|PT|646.50|Asymptomatic bacteriuria in pregnancy, unspecified as to episode of care or not applicable
C0156750|ICD9CM|AB|646.53|Asy bacteriuria-antepart
C0156750|ICD9CM|AB|646.50|Bacteriuria preg-unspec
C0156752|ICD9CM|PT|646.51|Asymptomatic bacteriuria in pregnancy, delivered, with or without mention of antepartum condition
C0156752|ICD9CM|AB|646.51|Asym bacteriuria-deliver
C0156753|ICD9CM|PT|646.52|Asymptomatic bacteriuria in pregnancy, delivered, with mention of postpartum complication
C0156753|ICD9CM|AB|646.52|Asy bacteruria-del w p/p
C0156755|ICD9CM|PT|646.54|Asymptomatic bacteriuria in pregnancy, postpartum condition or complication
C0156755|ICD9CM|AB|646.54|Asy bacteriuria-postpart
C0156756|ICD9CM|HT|646.6|Infections of genitourinary tract in pregnancy
C0156756|ICD9CM|PT|646.60|Infections of genitourinary tract in pregnancy, unspecified as to episode of care or not applicable
C0156756|ICD9CM|PT|646.63|Infections of genitourinary tract in pregnancy, antepartum condition or complication
C0156756|ICD9CM|AB|646.63|Gu infection-antepartum
C0156756|ICD9CM|AB|646.60|Gu infect in preg-unspec
C0156758|ICD9CM|PT|646.61|Infections of genitourinary tract in pregnancy, delivered, with or without mention of antepartum condition
C0156758|ICD9CM|AB|646.61|Gu infection-delivered
C0156759|ICD9CM|PT|646.62|Infections of genitourinary tract in pregnancy, delivered, with mention of postpartum complication
C0156759|ICD9CM|AB|646.62|Gu infection-deliv w p/p
C0156761|ICD9CM|PT|646.64|Infections of genitourinary tract in pregnancy, postpartum condition or complication
C0156761|ICD9CM|AB|646.64|Gu infection-postpartum
C0156762|ICD9CM|PT|646.70|Liver and biliary tract disorders in pregnancy, unspecified as to episode of care or not applicable
C0156762|ICD9CM|PT|646.73|Liver and biliary tract disorders in pregnancy, antepartum condition or complication
C0156762|ICD9CM|AB|646.70|Liver/bil trct disr-unsp
C0156762|ICD9CM|AB|646.73|Liver/bil trct disr-ante
C0156767|ICD9CM|PT|646.81|Other specified complications of pregnancy, delivered, with or without mention of antepartum condition
C0156767|ICD9CM|AB|646.81|Preg compl NEC-delivered
C0156768|ICD9CM|PT|646.82|Other specified complications of pregnancy, delivered, with mention of postpartum complication
C0156768|ICD9CM|AB|646.82|Preg compl NEC-del w p/p
C0156769|ICD9CM|PT|646.83|Other specified complications of pregnancy, antepartum condition or complication
C0156769|ICD9CM|HT|646.8|Other specified complications of pregnancy
C0156769|ICD9CM|PT|646.80|Other specified complications of pregnancy, unspecified as to episode of care or not applicable
C0156769|ICD9CM|AB|646.83|Preg compl NEC-antepart
C0156769|ICD9CM|AB|646.80|Preg compl NEC-unspec
C0156770|ICD9CM|PT|646.84|Other specified complications of pregnancy, postpartum condition or complication
C0156770|ICD9CM|AB|646.84|Preg compl NEC-postpart
C0156771|ICD9CM|PT|646.90|Unspecified complication of pregnancy, unspecified as to episode of care or not applicable
C0156771|ICD9CM|AB|646.90|Preg compl NOS-unspec
C0156772|ICD9CM|PT|646.91|Unspecified complication of pregnancy, delivered, with or without mention of antepartum condition
C0156772|ICD9CM|AB|646.91|Preg compl NOS-delivered
C0156773|ICD9CM|PT|646.93|Unspecified complication of pregnancy, antepartum condition or complication
C0156773|ICD9CM|AB|646.93|Preg compl NOS-antepart
C0156776|ICD9CM|PT|647.00|Syphilis of mother, complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C0156776|ICD9CM|AB|647.00|Syphilis in preg-unspec
C0156777|ICD9CM|PT|647.01|Syphilis of mother, complicating pregnancy, childbirth, or the puerperium, delivered, with or without mention of antepartum condition
C0156777|ICD9CM|AB|647.01|Syphilis-delivered
C0156778|ICD9CM|PT|647.02|Syphilis of mother, complicating pregnancy, childbirth, or the puerperium, delivered, with mention of postpartum complication
C0156778|ICD9CM|AB|647.02|Syphilis-delivered w p/p
C0156780|ICD9CM|AB|647.04|Syphilis-postpartum
C0156780|ICD9CM|PT|647.04|Syphilis of mother, complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication
C0156782|ICD9CM|PT|647.10|Gonorrhea of mother, complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C0156782|ICD9CM|AB|647.10|Gonorrhea in preg-unspec
C0156783|ICD9CM|PT|647.11|Gonorrhea of mother, complicating pregnancy, childbirth, or the puerperium, delivered, with or without mention of antepartum condition
C0156783|ICD9CM|AB|647.11|Gonorrhea-delivered
C0156784|ICD9CM|PT|647.12|Gonorrhea of mother, complicating pregnancy, childbirth, or the puerperium, delivered, with mention of postpartum complication
C0156784|ICD9CM|AB|647.12|Gonorrhea-deliver w p/p
C0156788|ICD9CM|PT|647.20|Other venereal diseases of mother, complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C0156788|ICD9CM|AB|647.20|Other VD in preg-unspec
C0156794|ICD9CM|PT|647.30|Tuberculosis of mother, complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C0156794|ICD9CM|AB|647.30|TB in preg-unspecified
C0156795|ICD9CM|PT|647.31|Tuberculosis of mother, complicating pregnancy, childbirth, or the puerperium, delivered, with or without mention of antepartum condition
C0156795|ICD9CM|AB|647.31|Tuberculosis-delivered
C0156796|ICD9CM|PT|647.32|Tuberculosis of mother, complicating pregnancy, childbirth, or the puerperium, delivered, with mention of postpartum complication
C0156796|ICD9CM|AB|647.32|Tuberculosis-deliv w p/p
C0156797|ICD9CM|AB|647.33|Tuberculosis-antepartum
C0156797|ICD9CM|PT|647.33|Tuberculosis of mother, complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C0156798|ICD9CM|AB|647.34|Tuberculosis-postpartum
C0156798|ICD9CM|PT|647.34|Tuberculosis of mother, complicating pregnancy, childbirth, or the puerperium,postpartum condition or complication
C0156799|ICD9CM|HT|647.4|Malaria complicating pregnancy, childbirth, or the puerperium
C0156800|ICD9CM|PT|647.40|Malaria in the mother, unspecified as to episode of care or not applicable
C0156800|ICD9CM|AB|647.40|Malaria in preg-unspec
C0156801|ICD9CM|PT|647.41|Malaria in the mother, delivered, with or without mention of antepartum condition
C0156801|ICD9CM|AB|647.41|Malaria-delivered
C0156802|ICD9CM|PT|647.42|Malaria in the mother, delivered, with mention of postpartum complication
C0156802|ICD9CM|AB|647.42|Malaria-delivered w p/p
C0156804|ICD9CM|AB|647.44|Malaria-postpartum
C0156804|ICD9CM|PT|647.44|Malaria in the mother, postpartum condition or complication
C0156805|ICD9CM|HT|647.5|Rubella complicating pregnancy, childbirth, or the puerperium
C0156807|ICD9CM|PT|647.51|Rubella in the mother, delivered, with or without mention of antepartum condition
C0156807|ICD9CM|AB|647.51|Rubella-delivered
C0156808|ICD9CM|PT|647.52|Rubella in the mother, delivered, with mention of postpartum complication
C0156808|ICD9CM|AB|647.52|Rubella-delivered w p/p
C0156809|ICD9CM|AB|647.53|Rubella-antepartum
C0156809|ICD9CM|PT|647.53|Rubella in the mother, antepartum condition or complication
C0156810|ICD9CM|AB|647.54|Rubella-postpartum
C0156810|ICD9CM|PT|647.54|Rubella in the mother, postpartum condition or complication
C0156812|ICD9CM|PT|647.60|Other viral diseases in the mother, unspecified as to episode of care or not applicable
C0156812|ICD9CM|AB|647.60|Oth virus in preg-unspec
C0156813|ICD9CM|PT|647.61|Other viral diseases in the mother, delivered, with or without mention of antepartum condition
C0156813|ICD9CM|AB|647.61|Oth viral dis-delivered
C0156814|ICD9CM|PT|647.62|Other viral diseases in the mother, delivered, with mention of postpartum complication
C0156814|ICD9CM|AB|647.62|Oth viral dis-del w p/p
C0156815|ICD9CM|PT|647.63|Other viral diseases in the mother, antepartum condition or complication
C0156815|ICD9CM|AB|647.63|Oth viral dis-antepartum
C0156816|ICD9CM|PT|647.64|Other viral diseases in the mother, postpartum condition or complication
C0156816|ICD9CM|AB|647.64|Oth viral dis-postpartum
C0156818|ICD9CM|PT|647.80|Other specified infectious and parasitic diseases of mother, unspecified as to episode of care or not applicable
C0156818|ICD9CM|AB|647.80|Inf dis in preg NEC-unsp
C0156819|ICD9CM|PT|647.81|Other specified infectious and parasitic diseases of mother, delivered, with or without mention of antepartum condition
C0156819|ICD9CM|AB|647.81|Infect dis NEC-delivered
C0156820|ICD9CM|PT|647.82|Other specified infectious and parasitic diseases of mother, delivered, with mention of postpartum complication
C0156820|ICD9CM|AB|647.82|Infect dis NEC-del w p/p
C0156821|ICD9CM|PT|647.83|Other specified infectious and parasitic diseases of mother, antepartum condition or complication
C0156821|ICD9CM|AB|647.83|Infect dis NEC-antepart
C0156822|ICD9CM|PT|647.84|Other specified infectious and parasitic diseases of mother, postpartum condition or complication
C0156822|ICD9CM|AB|647.84|Infect dis NEC-postpart
C0156823|ICD9CM|HT|647.9|Unspecified infection or infestation complicating pregnancy, childbirth, or the puerperium
C0156824|ICD9CM|PT|647.90|Unspecified infection or infestation of mother, unspecified as to episode of care or not applicable
C0156824|ICD9CM|AB|647.90|Infect in preg NOS-unsp
C0156825|ICD9CM|PT|647.91|Unspecified infection or infestation of mother, delivered, with or without mention of antepartum condition
C0156825|ICD9CM|AB|647.91|Infect NOS-delivered
C0156826|ICD9CM|PT|647.92|Unspecified infection or infestation of mother, delivered, with mention of postpartum complication
C0156826|ICD9CM|AB|647.92|Infect NOS-deliver w p/p
C0156827|ICD9CM|PT|647.93|Unspecified infection or infestation of mother, antepartum condition or complication
C0156827|ICD9CM|AB|647.93|Infect NOS-antepartum
C0156828|ICD9CM|PT|647.94|Unspecified infection or infestation of mother, postpartum condition or complication
C0156828|ICD9CM|AB|647.94|Infect NOS-postpartum
C0156837|ICD9CM|PT|648.10|Thyroid dysfunction of mother, unspecified as to episode of care or not applicable
C0156837|ICD9CM|AB|648.10|Thyroid dysfun preg-unsp
C0156838|ICD9CM|PT|648.11|Thyroid dysfunction of mother, delivered, with or without mention of antepartum condition
C0156838|ICD9CM|AB|648.11|Thyroid dysfunc-deliver
C0156839|ICD9CM|PT|648.12|Thyroid dysfunction of mother, delivered, with mention of postpartum complication
C0156839|ICD9CM|AB|648.12|Thyroid dysfun-del w p/p
C0156841|ICD9CM|PT|648.14|Thyroid dysfunction of mother, postpartum condition or complication
C0156841|ICD9CM|AB|648.14|Thyroid dysfunc-postpart
C0156844|ICD9CM|PT|648.21|Anemia of mother, delivered, with or without mention of antepartum condition
C0156844|ICD9CM|AB|648.21|Anemia-delivered
C0156845|ICD9CM|PT|648.22|Anemia of mother, delivered, with mention of postpartum complication
C0156845|ICD9CM|AB|648.22|Anemia-delivered w p/p
C0156847|ICD9CM|AB|648.24|Anemia-postpartum
C0156847|ICD9CM|PT|648.24|Anemia of mother, postpartum condition or complication
C0156850|ICD9CM|PT|648.31|Drug dependence of mother, delivered, with or without mention of antepartum condition
C0156850|ICD9CM|AB|648.31|Drug dependence-deliver
C0156851|ICD9CM|PT|648.32|Drug dependence of mother, delivered, with mention of postpartum complication
C0156851|ICD9CM|AB|648.32|Drug dependen-del w p/p
C0156852|ICD9CM|PT|648.33|Drug dependence of mother, antepartum condition or complication
C0156852|ICD9CM|AB|648.33|Drug dependence-antepart
C0156853|ICD9CM|PT|648.34|Drug dependence of mother, postpartum condition or complication
C0156853|ICD9CM|AB|648.34|Drug dependence-postpart
C0156854|ICD9CM|HT|648.4|Mental disorders complicating pregnancy, childbirth, or the puerperium
C0156855|ICD9CM|PT|648.40|Mental disorders of mother, unspecified as to episode of care or not applicable
C0156855|ICD9CM|AB|648.40|Mental dis preg-unspec
C0156856|ICD9CM|PT|648.41|Mental disorders of mother, delivered, with or without mention of antepartum condition
C0156856|ICD9CM|AB|648.41|Mental disorder-deliver
C0156857|ICD9CM|PT|648.42|Mental disorders of mother, delivered, with mention of postpartum complication
C0156857|ICD9CM|AB|648.42|Mental dis-deliv w p/p
C0156858|ICD9CM|PT|648.43|Mental disorders of mother, antepartum condition or complication
C0156858|ICD9CM|AB|648.43|Mental disorder-antepart
C0156859|ICD9CM|PT|648.44|Mental disorders of mother, postpartum condition or complication
C0156859|ICD9CM|AB|648.44|Mental disorder-postpart
C0156860|ICD9CM|HT|648.5|Congenital cardiovascular disorders complicating pregnancy, childbirth, or the puerperium
C0156861|ICD9CM|PT|648.50|Congenital cardiovascular disorders of mother, unspecified as to episode of care or not applicable
C0156861|ICD9CM|AB|648.50|Congen CV dis preg-unsp
C0156862|ICD9CM|PT|648.51|Congenital cardiovascular disorders of mother, delivered, with or without mention of antepartum condition
C0156862|ICD9CM|AB|648.51|Congen CV dis-delivered
C0156863|ICD9CM|PT|648.52|Congenital cardiovascular disorders of mother, delivered, with mention of postpartum complication
C0156863|ICD9CM|AB|648.52|Congen CV dis-del w p/p
C0156864|ICD9CM|PT|648.53|Congenital cardiovascular disorders of mother, antepartum condition or complication
C0156864|ICD9CM|AB|648.53|Congen CV dis-antepartum
C0156865|ICD9CM|PT|648.54|Congenital cardiovascular disorders of mother, postpartum condition or complication
C0156865|ICD9CM|AB|648.54|Congen CV dis-postpartum
C0156866|ICD9CM|HT|648.6|Other cardiovascular diseases complicating pregnancy, childbirth, or the puerperium
C0156867|ICD9CM|PT|648.60|Other cardiovascular diseases of mother, unspecified as to episode of care or not applicable
C0156867|ICD9CM|AB|648.60|CV dis NEC preg-unspec
C0156868|ICD9CM|PT|648.61|Other cardiovascular diseases of mother, delivered, with or without mention of antepartum condition
C0156868|ICD9CM|AB|648.61|CV dis NEC preg-deliver
C0156869|ICD9CM|PT|648.62|Other cardiovascular diseases of mother, delivered, with mention of postpartum complication
C0156869|ICD9CM|AB|648.62|CV dis NEC-deliver w p/p
C0156870|ICD9CM|PT|648.63|Other cardiovascular diseases of mother, antepartum condition or complication
C0156870|ICD9CM|AB|648.63|CV dis NEC-antepartum
C0156871|ICD9CM|PT|648.64|Other cardiovascular diseases of mother, postpartum condition or complication
C0156871|ICD9CM|AB|648.64|CV dis NEC-postpartum
C0156872|ICD9CM|HT|648.7|Bone and joint disorders of back, pelvis, and lower limbs of mother, complicating pregnancy, childbirth, or the puerperium
C0156873|ICD9CM|PT|648.70|Bone and joint disorders of back, pelvis, and lower limbs of mother, unspecified as to episode of care or not applicable
C0156873|ICD9CM|AB|648.70|Bone disord in preg-unsp
C0156874|ICD9CM|PT|648.71|Bone and joint disorders of back, pelvis, and lower limbs of mother, delivered, with or without mention of antepartum condition
C0156874|ICD9CM|AB|648.71|Bone disorder-delivered
C0156875|ICD9CM|PT|648.72|Bone and joint disorders of back, pelvis, and lower limbs of mother, delivered, with mention of postpartum complication
C0156875|ICD9CM|AB|648.72|Bone disorder-del w p/p
C0156876|ICD9CM|PT|648.73|Bone and joint disorders of back, pelvis, and lower limbs of mother, antepartum condition or complication
C0156876|ICD9CM|AB|648.73|Bone disorder-antepartum
C0156877|ICD9CM|PT|648.74|Bone and joint disorders of back, pelvis, and lower limbs of mother, postpartum condition or complication
C0156877|ICD9CM|AB|648.74|Bone disorder-postpartum
C0156878|ICD9CM|HT|648.8|Abnormal glucose tolerance of mother, complicating pregnancy, childbirth, or the puerperium
C0156879|ICD9CM|PT|648.80|Abnormal glucose tolerance of mother, unspecified as to episode of care or not applicable
C0156879|ICD9CM|AB|648.80|Abn glucose in preg-unsp
C0156880|ICD9CM|PT|648.81|Abnormal glucose tolerance of mother, delivered, with or without mention of antepartum condition
C0156880|ICD9CM|AB|648.81|Abn glucose toler-deliv
C0156881|ICD9CM|PT|648.82|Abnormal glucose tolerance of mother, delivered, with mention of postpartum complication
C0156881|ICD9CM|AB|648.82|Abn glucose-deliv w p/p
C0156882|ICD9CM|PT|648.83|Abnormal glucose tolerance of mother, antepartum condition or complication
C0156882|ICD9CM|AB|648.83|Abn glucose-antepartum
C0156883|ICD9CM|PT|648.84|Abnormal glucose tolerance of mother, postpartum condition or complication
C0156883|ICD9CM|AB|648.84|Abn glucose-postpartum
C0156884|ICD9CM|HT|648.9|Other current conditions complicating pregnancy, childbirth, or the puerperium
C0156885|ICD9CM|PT|648.90|Other current conditions classifiable elsewhere of mother, unspecified as to episode of care or not applicable
C0156885|ICD9CM|AB|648.90|Oth curr cond preg-unsp
C0156886|ICD9CM|PT|648.91|Other current conditions classifiable elsewhere of mother, delivered, with or without mention of antepartum condition
C0156886|ICD9CM|AB|648.91|Oth curr cond-delivered
C0156887|ICD9CM|PT|648.92|Other current conditions classifiable elsewhere of mother, delivered, with mention of postpartum complication
C0156887|ICD9CM|AB|648.92|Oth curr cond-del w p/p
C0156888|ICD9CM|PT|648.93|Other current conditions classifiable elsewhere of mother, antepartum condition or complication
C0156888|ICD9CM|AB|648.93|Oth curr cond-antepartum
C0156889|ICD9CM|PT|648.94|Other current conditions classifiable elsewhere of mother, postpartum condition or complication
C0156889|ICD9CM|AB|648.94|Oth curr cond-postpartum
C0156892|ICD9CM|PT|651.00|Twin pregnancy, unspecified as to episode of care or not applicable
C0156892|ICD9CM|AB|651.00|Twin pregnancy-unspec
C0156893|ICD9CM|AB|651.01|Twin pregnancy-delivered
C0156893|ICD9CM|PT|651.01|Twin pregnancy, delivered, with or without mention of antepartum condition
C0156894|ICD9CM|PT|651.03|Twin pregnancy, antepartum condition or complication
C0156894|ICD9CM|AB|651.03|Twin pregnancy-antepart
C0156895|ICD9CM|PT|651.10|Triplet pregnancy, unspecified as to episode of care or not applicable
C0156895|ICD9CM|AB|651.10|Triplet pregnancy-unspec
C0156896|ICD9CM|PT|651.11|Triplet pregnancy, delivered, with or without mention of antepartum condition
C0156896|ICD9CM|AB|651.11|Triplet pregnancy-deliv
C0156897|ICD9CM|PT|651.13|Triplet pregnancy, antepartum condition or complication
C0156897|ICD9CM|AB|651.13|Triplet preg-antepartum
C0156898|ICD9CM|PT|651.20|Quadruplet pregnancy, unspecified as to episode of care or not applicable
C0156898|ICD9CM|AB|651.20|Quadruplet preg-unspec
C0156899|ICD9CM|PT|651.21|Quadruplet pregnancy, delivered, with or without mention of antepartum condition
C0156899|ICD9CM|AB|651.21|Quadruplet preg-deliver
C0156900|ICD9CM|PT|651.23|Quadruplet pregnancy, antepartum condition or complication
C0156900|ICD9CM|AB|651.23|Quadruplet preg-antepart
C0156901|ICD9CM|HT|651.3|Twin pregnancy with fetal loss and retention of one fetus
C0156902|ICD9CM|PT|651.30|Twin pregnancy with fetal loss and retention of one fetus, unspecified as to episode of care or not applicable
C0156902|ICD9CM|AB|651.30|Twins w fetal loss-unsp
C0156903|ICD9CM|PT|651.31|Twin pregnancy with fetal loss and retention of one fetus, delivered, with or without mention of antepartum condition
C0156903|ICD9CM|AB|651.31|Twins w fetal loss-del
C0156904|ICD9CM|PT|651.33|Twin pregnancy with fetal loss and retention of one fetus, antepartum condition or complication
C0156904|ICD9CM|AB|651.33|Twins w fetal loss-ante
C0156905|ICD9CM|HT|651.4|Triplet pregnancy with fetal loss and retention of one or more fetus (es)
C0156906|ICD9CM|PT|651.40|Triplet pregnancy with fetal loss and retention of one or more fetus(es), unspecified as to episode of care or not applicable
C0156906|ICD9CM|AB|651.40|Triplets w fet loss-unsp
C0156907|ICD9CM|PT|651.41|Triplet pregnancy with fetal loss and retention of one or more fetus(es), delivered, with or without mention of antepartum condition
C0156907|ICD9CM|AB|651.41|Triplets w fet loss-del
C0156908|ICD9CM|PT|651.43|Triplet pregnancy with fetal loss and retention of one or more fetus(es), antepartum condition or complication
C0156908|ICD9CM|AB|651.43|Triplets w fet loss-ante
C0156909|ICD9CM|HT|651.5|Quadruplet pregnancy with fetal loss and retention of one or more fetus(es)
C0156910|ICD9CM|PT|651.50|Quadruplet pregnancy with fetal loss and retention of one or more fetus(es), unspecified as to episode of care or not applicable
C0156910|ICD9CM|AB|651.50|Quads w fetal loss-unsp
C0156911|ICD9CM|PT|651.51|Quadruplet pregnancy with fetal loss and retention of one or more fetus(es), delivered, with or without mention of antepartum condition
C0156911|ICD9CM|AB|651.51|Quads w fetal loss-del
C0156912|ICD9CM|PT|651.53|Quadruplet pregnancy with fetal loss and retention of one or more fetus(es), antepartum condition or complication
C0156912|ICD9CM|AB|651.53|Quads w fetal loss-ante
C0156913|ICD9CM|HT|651.6|Other multiple pregnancy with fetal loss and retention of one or more fetus(es)
C0156914|ICD9CM|PT|651.60|Other multiple pregnancy with fetal loss and retention of one or more fetus(es), unspecified as to episode of care or not applicable
C0156914|ICD9CM|AB|651.60|Mult ges w fet loss-unsp
C0156915|ICD9CM|PT|651.61|Other multiple pregnancy with fetal loss and retention of one or more fetus(es), delivered, with or without mention of antepartum condition
C0156915|ICD9CM|AB|651.61|Mult ges w fet loss-del
C0156916|ICD9CM|PT|651.63|Other multiple pregnancy with fetal loss and retention of one or more fetus(es), antepartum condition or complication
C0156916|ICD9CM|AB|651.63|Mult ges w fet loss-ante
C0156917|ICD9CM|HT|651.8|Other specified multiple gestation
C0156918|ICD9CM|PT|651.80|Other specified multiple gestation, unspecified as to episode of care or not applicable
C0156918|ICD9CM|AB|651.80|Multi gestat NEC-unspec
C0156919|ICD9CM|PT|651.81|Other specified multiple gestation, delivered, with or without mention of antepartum condition
C0156919|ICD9CM|AB|651.81|Multi gestat NEC-deliver
C0156920|ICD9CM|PT|651.83|Other specified multiple gestation, antepartum condition or complication
C0156920|ICD9CM|AB|651.83|Multi gest NEC-antepart
C0156922|ICD9CM|PT|651.91|Unspecified multiple gestation, delivered, with or without mention of antepartum condition
C0156922|ICD9CM|AB|651.91|Mult gestation NOS-deliv
C0156923|ICD9CM|PT|651.93|Unspecified multiple gestation, antepartum condition or complication
C0156923|ICD9CM|AB|651.93|Multi gest NOS-antepart
C0156924|ICD9CM|HT|652|Malposition and malpresentation of fetus
C0156924|ICD9CM|HT|652.9|Unspecified malposition or malpresentation of fetus
C0156926|ICD9CM|PT|652.00|Unstable lie, unspecified as to episode of care or not applicable
C0156926|ICD9CM|AB|652.00|Unstable lie-unspecified
C0156927|ICD9CM|AB|652.01|Unstable lie-delivered
C0156927|ICD9CM|PT|652.01|Unstable lie, delivered, with or without mention of antepartum condition
C0156928|ICD9CM|PT|652.03|Unstable lie, antepartum condition or complication
C0156928|ICD9CM|AB|652.03|Unstable lie-antepartum
C0156929|ICD9CM|HT|652.1|Breech or other malpresentation successfully converted to cephalic presentation
C0156930|ICD9CM|PT|652.10|Breech or other malpresentation successfully converted to cephalic presentation, unspecified as to episode of care or not applicable
C0156930|ICD9CM|AB|652.10|Cephalic vers NOS-unspec
C0156931|ICD9CM|PT|652.11|Breech or other malpresentation successfully converted to cephalic presentation, delivered, with or without mention of antepartum condition
C0156931|ICD9CM|AB|652.11|Cephalic vers NOS-deliv
C0156932|ICD9CM|PT|652.13|Breech or other malpresentation successfully converted to cephalic presentation, antepartum condition or complication
C0156932|ICD9CM|AB|652.13|Cephal vers NOS-antepart
C0156933|ICD9CM|PT|652.20|Breech presentation without mention of version, unspecified as to episode of care or not applicable
C0156933|ICD9CM|AB|652.20|Breech presentat-unspec
C0156934|ICD9CM|PT|652.21|Breech presentation without mention of version, delivered, with or without mention of antepartum condition
C0156934|ICD9CM|AB|652.21|Breech presentat-deliver
C0156935|ICD9CM|PT|652.23|Breech presentation without mention of version, antepartum condition or complication
C0156935|ICD9CM|AB|652.23|Breech present-antepart
C0156936|ICD9CM|HT|652.3|Transverse or oblique presentation of fetus
C0156940|ICD9CM|HT|652.4|Face or brow presentation of fetus
C0156941|ICD9CM|PT|652.40|Face or brow presentation, unspecified as to episode of care or not applicable
C0156941|ICD9CM|AB|652.40|Face/brow present-unspec
C0156942|ICD9CM|PT|652.41|Face or brow presentation, delivered, with or without mention of antepartum condition
C0156942|ICD9CM|AB|652.41|Face/brow present-deliv
C0156943|ICD9CM|PT|652.43|Face or brow presentation, antepartum condition or complication
C0156943|ICD9CM|AB|652.43|Face/brow pres-antepart
C0156945|ICD9CM|PT|652.50|High head at term, unspecified as to episode of care or not applicable
C0156945|ICD9CM|AB|652.50|High head at term-unspec
C0156946|ICD9CM|PT|652.51|High head at term, delivered, with or without mention of antepartum condition
C0156946|ICD9CM|AB|652.51|High head at term-deliv
C0156947|ICD9CM|PT|652.53|High head at term, antepartum condition or complication
C0156947|ICD9CM|AB|652.53|High head term-antepart
C0156948|ICD9CM|HT|652.6|Multiple gestation with malpresentation of one fetus or more
C0156949|ICD9CM|PT|652.60|Multiple gestation with malpresentation of one fetus or more, unspecified as to episode of care or not applicable
C0156949|ICD9CM|AB|652.60|Mult gest malpresen-unsp
C0156950|ICD9CM|PT|652.61|Multiple gestation with malpresentation of one fetus or more, delivered, with or without mention of antepartum condition
C0156950|ICD9CM|AB|652.61|Mult gest malpres-deliv
C0156951|ICD9CM|PT|652.63|Multiple gestation with malpresentation of one fetus or more, antepartum condtion or complication
C0156951|ICD9CM|AB|652.63|Mult ges malpres-antepar
C0156953|ICD9CM|PT|652.70|Prolapsed arm of fetus, unspecified as to episode of care or not applicable
C0156953|ICD9CM|AB|652.70|Prolapsed arm-unspec
C0156954|ICD9CM|AB|652.71|Prolapsed arm-delivered
C0156954|ICD9CM|PT|652.71|Prolapsed arm of fetus, delivered, with or without mention of antepartum condition
C0156955|ICD9CM|AB|652.73|Prolapsed arm-antepart
C0156955|ICD9CM|PT|652.73|Prolapsed arm of fetus, antepartum condition or complication
C0156956|ICD9CM|HT|652.8|Other specified malposition or malpresentation of fetus
C0156957|ICD9CM|PT|652.80|Other specified malposition or malpresentation, unspecified as to episode of care or not applicable
C0156957|ICD9CM|AB|652.80|Malposition NEC-unspec
C0156958|ICD9CM|PT|652.81|Other specified malposition or malpresentation, delivered, with or without mention of antepartum condition
C0156958|ICD9CM|AB|652.81|Malposition NEC-deliver
C0156959|ICD9CM|PT|652.83|Other specified malposition or malpresentation, antepartum condition or complication
C0156959|ICD9CM|AB|652.83|Malposition NEC-antepart
C0156961|ICD9CM|PT|652.90|Unspecified malposition or malpresentation, unspecified as to episode of care or not applicable
C0156961|ICD9CM|AB|652.90|Malposition NOS-unspec
C0156962|ICD9CM|PT|652.91|Unspecified malposition or malpresentation, delivered, with or without mention of antepartum condition
C0156962|ICD9CM|AB|652.91|Malposition NOS-deliver
C0156963|ICD9CM|PT|652.93|Unspecified malposition or malpresentation, antepartum condition or complication
C0156963|ICD9CM|AB|652.93|Malposition NOS-antepart
C0156964|ICD9CM|HT|653|Disproportion in pregnancy, labor, and delivery
C0156966|ICD9CM|PT|653.00|Major abnormality of bony pelvis, not further specified, unspecified as to episode of care or not applicable
C0156966|ICD9CM|AB|653.00|Pelvic deform NOS-unspec
C0156967|ICD9CM|PT|653.01|Major abnormality of bony pelvis, not further specified, delivered, with or without mention of antepartum condition
C0156967|ICD9CM|AB|653.01|Pelvic deform NOS-deliv
C0156968|ICD9CM|PT|653.03|Major abnormality of bony pelvis, not further specified, antepartum condition or complication
C0156968|ICD9CM|AB|653.03|Pelv deform NOS-antepart
C0156969|ICD9CM|HT|653.1|Generally contracted pelvis in pregnancy, labor, and delivery
C0156970|ICD9CM|PT|653.10|Generally contracted pelvis, unspecified as to episode of care or not applicable
C0156970|ICD9CM|AB|653.10|Contract pelv NOS-unspec
C0156971|ICD9CM|PT|653.11|Generally contracted pelvis, delivered, with or without mention of antepartum condition
C0156971|ICD9CM|AB|653.11|Contract pelv NOS-deliv
C0156972|ICD9CM|PT|653.13|Generally contracted pelvis, antepartum condition or complication
C0156972|ICD9CM|AB|653.13|Contrac pelv NOS-antepar
C0156973|ICD9CM|HT|653.2|Inlet contraction of pelvis in pregnancy, labor, and delivery
C0156974|ICD9CM|PT|653.20|Inlet contraction of pelvis, unspecified as to episode of care or not applicable
C0156974|ICD9CM|AB|653.20|Inlet contraction-unspec
C0156975|ICD9CM|PT|653.21|Inlet contraction of pelvis, delivered, with or without mention of antepartum condition
C0156975|ICD9CM|AB|653.21|Inlet contraction-deliv
C0156976|ICD9CM|PT|653.23|Inlet contraction of pelvis, antepartum condition or complication
C0156976|ICD9CM|AB|653.23|Inlet contract-antepart
C0156977|ICD9CM|HT|653.3|Outlet contraction of pelvis in pregnancy, labor, and delivery
C0156978|ICD9CM|PT|653.30|Outlet contraction of pelvis, unspecified as to episode of care or not applicable
C0156978|ICD9CM|AB|653.30|Outlet contraction-unsp
C0156979|ICD9CM|PT|653.31|Outlet contraction of pelvis, delivered, with or without mention of antepartum condition
C0156979|ICD9CM|AB|653.31|Outlet contraction-deliv
C0156980|ICD9CM|PT|653.33|Outlet contraction of pelvis, antepartum condition or complication
C0156980|ICD9CM|AB|653.33|Outlet contract-antepart
C0156982|ICD9CM|PT|653.41|Fetopelvic disproportion, delivered, with or without mention of antepartum condition
C0156982|ICD9CM|AB|653.41|Fetopelv dispropor-deliv
C0156984|ICD9CM|HT|653.5|Unusually large fetus causing disproportion
C0156985|ICD9CM|PT|653.50|Unusually large fetus causing disproportion, unspecified as to episode of care or not applicable
C0156985|ICD9CM|AB|653.50|Fetal disprop NOS-unspec
C0156986|ICD9CM|PT|653.51|Unusually large fetus causing disproportion, delivered, with or without mention of antepartum condition
C0156986|ICD9CM|AB|653.51|Fetal disprop NOS-deliv
C0156987|ICD9CM|PT|653.53|Unusually large fetus causing disproportion, antepartum condition or complication
C0156987|ICD9CM|AB|653.53|Fetal dispro NOS-antepar
C0156989|ICD9CM|PT|653.60|Hydrocephalic fetus causing disproportion, unspecified as to episode of care or not applicable
C0156989|ICD9CM|AB|653.60|Hydrocephal fetus-unspec
C0156990|ICD9CM|PT|653.61|Hydrocephalic fetus causing disproportion, delivered, with or without mention of antepartum condition
C0156990|ICD9CM|AB|653.61|Hydroceph fetus-deliver
C0156991|ICD9CM|PT|653.63|Hydrocephalic fetus causing disproportion, antepartum condition or complication
C0156991|ICD9CM|AB|653.63|Hydroceph fetus-antepart
C0156993|ICD9CM|PT|653.70|Other fetal abnormality causing disproportion, unspecified as to episode of care or not applicable
C0156993|ICD9CM|AB|653.70|Oth abn fet disprop-unsp
C0156994|ICD9CM|PT|653.71|Other fetal abnormality causing disproportion, delivered, with or without mention of antepartum condition
C0156994|ICD9CM|AB|653.71|Oth abn fet dispro-deliv
C0156995|ICD9CM|PT|653.73|Other fetal abnormality causing disproportion, antepartum condition or complication
C0156995|ICD9CM|AB|653.73|Oth abn fet dispro-antep
C0156996|ICD9CM|HT|653.8|Disproportion of other origin in pregnancy, labor, and delivery
C0156997|ICD9CM|PT|653.80|Disproportion of other origin, unspecified as to episode of care or not applicable
C0156997|ICD9CM|AB|653.80|Disproportion NEC-unspec
C0156998|ICD9CM|PT|653.81|Disproportion of other origin, delivered, with or without mention of antepartum condition
C0156998|ICD9CM|AB|653.81|Disproportion NEC-deliv
C0156999|ICD9CM|PT|653.83|Disproportion of other origin, antepartum condition or complication
C0156999|ICD9CM|AB|653.83|Dispropor NEC-antepartum
C0157000|ICD9CM|HT|653.9|Unspecified disproportion in pregnancy, labor, and delivery
C0157001|ICD9CM|PT|653.90|Unspecified disproportion, unspecified as to episode of care or not applicable
C0157001|ICD9CM|AB|653.90|Disproportion NOS-unspec
C0157002|ICD9CM|PT|653.91|Unspecified disproportion, delivered, with or without mention of antepartum condition
C0157002|ICD9CM|AB|653.91|Disproportion NOS-deliv
C0157003|ICD9CM|PT|653.93|Unspecified disproportion, antepartum condition or complication
C0157003|ICD9CM|AB|653.93|Dispropor NOS-antepartum
C0157004|ICD9CM|HT|654|Abnormality of organs and soft tissues of pelvis complicating pregnancy, childbirth, or the puerperium
C0157005|ICD9CM|HT|654.0|Congenital abnormalities of uterus complicating pregnancy, childbirth, or the puerperium
C0157006|ICD9CM|PT|654.00|Congenital abnormalities of uterus, unspecified as to episode of care or not applicable
C0157006|ICD9CM|AB|654.00|Cong abn uter preg-unsp
C0157007|ICD9CM|PT|654.01|Congenital abnormalities of uterus, delivered, with or without mention of antepartum condition
C0157007|ICD9CM|AB|654.01|Congen abn uterus-deliv
C0157008|ICD9CM|PT|654.02|Congenital abnormalities of uterus, delivered, with mention of postpartum complication
C0157008|ICD9CM|AB|654.02|Cong abn uter-del w p/p
C0157009|ICD9CM|PT|654.03|Congenital abnormalities of uterus, antepartum condition or complication
C0157009|ICD9CM|AB|654.03|Congen abn uter-antepart
C0157010|ICD9CM|PT|654.04|Congenital abnormalities of uterus, postpartum condition or complication
C0157010|ICD9CM|AB|654.04|Congen abn uter-postpart
C0157011|ICD9CM|HT|654.1|Tumors of body of uterus complicating pregnancy, childbirth, or the puerperium
C0157012|ICD9CM|PT|654.10|Tumors of body of uterus, unspecified as to episode of care or not applicable
C0157012|ICD9CM|AB|654.10|Uter tumor in preg-unsp
C0157013|ICD9CM|PT|654.11|Tumors of body of uterus, delivered, with or without mention of antepartum condition
C0157013|ICD9CM|AB|654.11|Uterine tumor-delivered
C0157014|ICD9CM|PT|654.12|Tumors of body of uterus, delivered, with mention of postpartum complication
C0157014|ICD9CM|AB|654.12|Uterine tumor-del w p/p
C0157015|ICD9CM|PT|654.13|Tumors of body of uterus, antepartum condition or complication
C0157015|ICD9CM|AB|654.13|Uterine tumor-antepartum
C0157016|ICD9CM|PT|654.14|Tumors of body of uterus, postpartum condition or complication
C0157016|ICD9CM|AB|654.14|Uterine tumor-postpartum
C0157018|ICD9CM|PT|654.20|Previous cesarean delivery, unspecified as to episode of care or not applicable
C0157018|ICD9CM|AB|654.20|Prev c-delivery unspec
C0157020|ICD9CM|PT|654.23|Previous cesarean delivery, antepartum condition or complication
C0157020|ICD9CM|AB|654.23|Prev c-delivery-antepart
C0157022|ICD9CM|PT|654.30|Retroverted and incarcerated gravid uterus, unspecified as to episode of care or not applicable
C0157022|ICD9CM|AB|654.30|Retrovert uterus-unspec
C0157023|ICD9CM|PT|654.31|Retroverted and incarcerated gravid uterus, delivered, with mention of antepartum condition
C0157023|ICD9CM|AB|654.31|Retrovert uterus-deliver
C0157024|ICD9CM|PT|654.32|Retroverted and incarcerated gravid uterus, delivered, with mention of postpartum complication
C0157024|ICD9CM|AB|654.32|Retrovert uter-del w p/p
C0157025|ICD9CM|AB|654.33|Retrovert uter-antepart
C0157025|ICD9CM|PT|654.33|Retroverted and incarcerated gravid uterus, antepartum condition or complication
C0157026|ICD9CM|AB|654.34|Retrovert uter-postpart
C0157026|ICD9CM|PT|654.34|Retroverted and incarcerated gravid uterus, postpartum condition or complication
C0157028|ICD9CM|PT|654.40|Other abnormalities in shape or position of gravid uterus and of neighboring structures, unspecified as to episode of care or not applicable
C0157028|ICD9CM|AB|654.40|Abn grav uterus NEC-unsp
C0157029|ICD9CM|PT|654.41|Other abnormalities in shape or position of gravid uterus and of neighboring structures, delivered, with or without mention of antepartum condition
C0157029|ICD9CM|AB|654.41|Abn uterus NEC-delivered
C0157030|ICD9CM|PT|654.42|Other abnormalities in shape or position of gravid uterus and of neighboring structures, delivered, with mention of postpartum complication
C0157030|ICD9CM|AB|654.42|Abn uterus NEC-del w p/p
C0157031|ICD9CM|PT|654.43|Other abnormalities in shape or position of gravid uterus and of neighboring structures, antepartum condition or complication
C0157031|ICD9CM|AB|654.43|Abn uterus NEC-antepart
C0157032|ICD9CM|PT|654.44|Other abnormalities in shape or position of gravid uterus and of neighboring structures, postpartum condition or complication
C0157032|ICD9CM|AB|654.44|Abn uterus NEC-postpart
C0157033|ICD9CM|HT|654.5|Cervical incompetence complicating pregnancy, childbirth, or the puerperium
C0157034|ICD9CM|PT|654.50|Cervical incompetence, unspecified as to episode of care or not applicable
C0157034|ICD9CM|AB|654.50|Cerv incompet preg-unsp
C0157035|ICD9CM|PT|654.51|Cervical incompetence, delivered, with or without mention of antepartum condition
C0157035|ICD9CM|AB|654.51|Cervical incompet-deliv
C0157036|ICD9CM|PT|654.52|Cervical incompetence, delivered, with mention of postpartum complication
C0157036|ICD9CM|AB|654.52|Cerv incompet-del w p/p
C0157037|ICD9CM|PT|654.53|Cervical incompetence, antepartum condition or complication
C0157037|ICD9CM|AB|654.53|Cerv incompet-antepartum
C0157038|ICD9CM|PT|654.54|Cervical incompetence, postpartum condition or complication
C0157038|ICD9CM|AB|654.54|Cerv incompet-postpartum
C0157039|ICD9CM|HT|654.6|Other congenital or acquired abnormality of cervix complicating pregnancy, childbirth, or the puerperium
C0157040|ICD9CM|PT|654.60|Other congenital or acquired abnormality of cervix, unspecified as to episode of care or not applicable
C0157040|ICD9CM|AB|654.60|Abn cervix NEC preg-unsp
C0157041|ICD9CM|PT|654.61|Other congenital or acquired abnormality of cervix, delivered, with or without mention of antepartum condition
C0157041|ICD9CM|AB|654.61|Abn cervix NEC-delivered
C0157042|ICD9CM|PT|654.62|Other congenital or acquired abnormality of cervix, delivered, with mention of postpartum complication
C0157042|ICD9CM|AB|654.62|Abn cervix NEC-del w p/p
C0157043|ICD9CM|PT|654.63|Other congenital or acquired abnormality of cervix, antepartum condition or complication
C0157043|ICD9CM|AB|654.63|Abn cervix NEC-antepart
C0157044|ICD9CM|PT|654.64|Other congenital or acquired abnormality of cervix, postpartum condition or complication
C0157044|ICD9CM|AB|654.64|Abn cervix NEC-postpart
C0157045|ICD9CM|HT|654.7|Congenital or acquired abnormality of vagina complicating pregnancy, childbirth, or the puerperium
C0157046|ICD9CM|PT|654.70|Congenital or acquired abnormality of vagina, unspecified as to episode of care or not applicable
C0157046|ICD9CM|AB|654.70|Abn vagina in preg-unsp
C0157047|ICD9CM|PT|654.71|Congenital or acquired abnormality of vagina, delivered, with or without mention of antepartum condition
C0157047|ICD9CM|AB|654.71|Abnorm vagina-delivered
C0157048|ICD9CM|PT|654.72|Congenital or acquired abnormality of vagina, delivered, with mention of postpartum complication
C0157048|ICD9CM|AB|654.72|Abnorm vagina-del w p/p
C0157049|ICD9CM|PT|654.73|Congenital or acquired abnormality of vagina, antepartum condition or complication
C0157049|ICD9CM|AB|654.73|Abnorm vagina-antepartum
C0157050|ICD9CM|PT|654.74|Congenital or acquired abnormality of vagina, postpartum condition or complication
C0157050|ICD9CM|AB|654.74|Abnorm vagina-postpartum
C0157051|ICD9CM|HT|654.8|Congenital or acquired abnormality of vulva complicating pregnancy, childbirth, or the puerperium
C0157052|ICD9CM|PT|654.80|Congenital or acquired abnormality of vulva, unspecified as to episode of care or not applicable
C0157052|ICD9CM|AB|654.80|Abn vulva in preg-unspec
C0157053|ICD9CM|PT|654.81|Congenital or acquired abnormality of vulva, delivered, with or without mention of antepartum condition
C0157053|ICD9CM|AB|654.81|Abnormal vulva-delivered
C0157054|ICD9CM|PT|654.82|Congenital or acquired abnormality of vulva, delivered, with mention of postpartum complication
C0157054|ICD9CM|AB|654.82|Abnormal vulva-del w p/p
C0157055|ICD9CM|PT|654.83|Congenital or acquired abnormality of vulva, antepartum condition or complication
C0157055|ICD9CM|AB|654.83|Abnormal vulva-antepart
C0157056|ICD9CM|PT|654.84|Congenital or acquired abnormality of vulva, postpartum condition or complication
C0157056|ICD9CM|AB|654.84|Abnormal vulva-postpart
C0157057|ICD9CM|HT|654.9|Other and unspecified abnormality of organs and soft tissues of pelvis complicating pregnancy, childbirth, and the puerperium
C0157058|ICD9CM|PT|654.90|Other and unspecified abnormality of organs and soft tissues of pelvis, unspecified as to episode of care or not applicable
C0157058|ICD9CM|AB|654.90|Abn pel NEC in preg-unsp
C0157059|ICD9CM|PT|654.91|Other and unspecified abnormality of organs and soft tissues of pelvis, delivered, with or without mention of antepartum condition
C0157059|ICD9CM|AB|654.91|Abn pelv org NEC-deliver
C0157060|ICD9CM|PT|654.92|Other and unspecified abnormality of organs and soft tissues of pelvis, delivered, with mention of postpartum complication
C0157060|ICD9CM|AB|654.92|Abn pelv NEC-deliv w p/p
C0157061|ICD9CM|PT|654.93|Other and unspecified abnormality of organs and soft tissues of pelvis, antepartum condition or complication
C0157061|ICD9CM|AB|654.93|Abn pelv org NEC-antepar
C0157062|ICD9CM|PT|654.94|Other and unspecified abnormality of organs and soft tissues of pelvis, postpartum condition or complication
C0157062|ICD9CM|AB|654.94|Abn pelv org NEC-postpar
C0157063|ICD9CM|HT|655|Known or suspected fetal abnormality affecting management of mother
C0157063|ICD9CM|HT|655.9|Unspecified, known or suspected fetal abnormality affecting management of mother
C0157064|ICD9CM|HT|655.0|Central nervous system malformation in fetus affecting management of mother
C0157065|ICD9CM|PT|655.00|Central nervous system malformation in fetus, unspecified as to episode of care or not applicable
C0157065|ICD9CM|AB|655.00|Fetal cns malform-unspec
C0157066|ICD9CM|PT|655.01|Central nervous system malformation in fetus, delivered, with or without mention of antepartum condition
C0157066|ICD9CM|AB|655.01|Fetal cns malform-deliv
C0157067|ICD9CM|PT|655.03|Central nervous system malformation in fetus, antepartum condition or complication
C0157067|ICD9CM|AB|655.03|Fetal cns malfor-antepar
C0157068|ICD9CM|HT|655.1|Chromosomal abnormality in fetus affecting management of mother
C0157069|ICD9CM|PT|655.10|Chromosomal abnormality in fetus, affecting management of mother, unspecified as to episode of care or not applicable
C0157069|ICD9CM|AB|655.10|Fetal chromos abn-unspec
C0157070|ICD9CM|PT|655.11|Chromosomal abnormality in fetus, affecting management of mother, delivered, with or without mention of antepartum condition
C0157070|ICD9CM|AB|655.11|Fetal chromoso abn-deliv
C0157071|ICD9CM|PT|655.13|Chromosomal abnormality in fetus, affecting management of mother, antepartum condition or complication
C0157071|ICD9CM|AB|655.13|Fet chromo abn-antepart
C0157072|ICD9CM|HT|655.2|Hereditary disease in family possibly affecting fetus, affecting management of mother
C0157073|ICD9CM|PT|655.20|Hereditary disease in family possibly affecting fetus, affecting management of mother, unspecified as to episode of care or not applicable
C0157073|ICD9CM|AB|655.20|Famil heredit dis-unspec
C0157074|ICD9CM|PT|655.21|Hereditary disease in family possibly affecting fetus, affecting management of mother, delivered, with or without mention of antepartum condition
C0157074|ICD9CM|AB|655.21|Famil heredit dis-deliv
C0157075|ICD9CM|PT|655.23|Hereditary disease in family possibly affecting fetus, affecting management of mother, antepartum condition or complication
C0157075|ICD9CM|AB|655.23|Famil hered dis-antepart
C0157076|ICD9CM|HT|655.3|Suspected damage to fetus from viral disease in the mother, affecting management of mother
C0157077|ICD9CM|PT|655.30|Suspected damage to fetus from viral disease in the mother, affecting management of mother, unspecified as to episode of care or not applicable
C0157077|ICD9CM|AB|655.30|Fet damg d/t virus-unsp
C0157078|ICD9CM|PT|655.31|Suspected damage to fetus from viral disease in the mother, affecting management of mother, delivered, with or without mention of antepartum condition
C0157078|ICD9CM|AB|655.31|Fet damg d/t virus-deliv
C0157079|ICD9CM|PT|655.33|Suspected damage to fetus from viral disease in the mother, affecting management of mother, antepartum condition or complication
C0157079|ICD9CM|AB|655.33|Fet damg d/t virus-antep
C0157080|ICD9CM|HT|655.4|Suspected damage to fetus from other disease in the mother, affecting management of mother
C0157081|ICD9CM|PT|655.40|Suspected damage to fetus from other disease in the mother, affecting management of mother, unspecified as to episode of care or not applicable
C0157081|ICD9CM|AB|655.40|Fet damg d/t dis-unspec
C0157082|ICD9CM|PT|655.41|Suspected damage to fetus from other disease in the mother, affecting management of mother, delivered, with or without mention of antepartum condition
C0157082|ICD9CM|AB|655.41|Fet damg d/t dis-deliver
C0157083|ICD9CM|PT|655.43|Suspected damage to fetus from other disease in the mother, affecting management of mother, antepartum condition or complication
C0157083|ICD9CM|AB|655.43|Fet damg d/t dis-antepar
C0157084|ICD9CM|HT|655.5|Suspected damage to fetus from drugs, affecting management of mother
C0157085|ICD9CM|PT|655.50|Suspected damage to fetus from drugs, affecting management of mother, unspecified as to episode of care or not applicable
C0157085|ICD9CM|AB|655.50|Fetal damg d/t drug-unsp
C0157086|ICD9CM|PT|655.51|Suspected damage to fetus from drugs, affecting management of mother, delivered, with or without mention of antepartum condition
C0157086|ICD9CM|AB|655.51|Fet damag d/t drug-deliv
C0157087|ICD9CM|PT|655.53|Suspected damage to fetus from drugs, affecting management of mother, antepartum condition or complication
C0157087|ICD9CM|AB|655.53|Fet damg d/t drug-antepa
C0157088|ICD9CM|HT|655.6|Suspected damage to fetus from radiation, affecting management of mother
C0157089|ICD9CM|PT|655.60|Suspected damage to fetus from radiation, affecting management of mother, unspecified as to episode of care or not applicable
C0157089|ICD9CM|AB|655.60|Radiat fetal damag-unsp
C0157090|ICD9CM|PT|655.61|Suspected damage to fetus from radiation, affecting management of mother, delivered,
C0157090|ICD9CM|AB|655.61|Radiat fetal damag-deliv
C0157091|ICD9CM|PT|655.63|Suspected damage to fetus from radiation, affecting management of mother, antepartum condition or complication
C0157091|ICD9CM|AB|655.63|Radiat fet damag-antepar
C0157093|ICD9CM|PT|655.80|Other known or suspected fetal abnormality, not elsewhere classified, affecting management of mother, unspecified as to episode of care or not applicable
C0157093|ICD9CM|AB|655.80|Fetal abnorm NEC-unspec
C0157094|ICD9CM|PT|655.81|Other known or suspected fetal abnormality, not elsewhere classified, affecting management of mother, delivered, with or without mention of antepartum condition
C0157094|ICD9CM|AB|655.81|Fetal abnorm NEC-deliver
C0157095|ICD9CM|PT|655.83|Other known or suspected fetal abnormality, not elsewhere classified, affecting management of mother, antepartum condition or complication
C0157095|ICD9CM|AB|655.83|Fetal abnorm NEC-antepar
C0157097|ICD9CM|PT|655.90|Unspecified suspected fetal abnormality, affecting management of mother, unspecified as to episode of care or not applicable
C0157097|ICD9CM|AB|655.90|Fetal abnorm NOS-unspec
C0157098|ICD9CM|PT|655.91|Unspecified suspected fetal abnormality, affecting management of mother, delivered, with or without mention of antepartum condition
C0157098|ICD9CM|AB|655.91|Fetal abnorm NOS-deliver
C0157099|ICD9CM|PT|655.93|Unspecified suspected fetal abnormality, affecting management of mother, antepartum condition or complication
C0157099|ICD9CM|AB|655.93|Fetal abnorm NOS-antepar
C0157101|ICD9CM|HT|656.0|Fetal-maternal hemorrhage affecting management of mother
C0157103|ICD9CM|PT|656.01|Fetal-maternal hemorrhage, delivered, with or without mention of antepartum condition
C0157103|ICD9CM|AB|656.01|Fetal-maternal hem-deliv
C0157104|ICD9CM|PT|656.03|Fetal-maternal hemorrhage, antepartum condition or complication
C0157104|ICD9CM|AB|656.03|Fetal-matern hem-antepar
C0157105|ICD9CM|PT|656.10|Rhesus isoimmunization, unspecified as to episode of care or not applicable
C0157105|ICD9CM|AB|656.10|Rh isoimmunization-unsp
C0157106|ICD9CM|PT|656.11|Rhesus isoimmunization, delivered, with or without mention of antepartum condition
C0157106|ICD9CM|AB|656.11|Rh isoimmunizat-deliver
C0157107|ICD9CM|PT|656.13|Rhesus isoimmunization, antepartum condition or complication
C0157107|ICD9CM|AB|656.13|Rh isoimmunizat-antepart
C0157108|ICD9CM|HT|656.2|Isoimmunization from other and unspecified blood-group incompatibility affecting management of mother
C0157109|ICD9CM|PT|656.20|Isoimmunization from other and unspecified blood-group incompatibility, unspecified as to episode of care or not applicable
C0157109|ICD9CM|AB|656.20|Abo isoimmunization-unsp
C0157110|ICD9CM|PT|656.21|Isoimmunization from other and unspecified blood-group incompatibility, delivered, with or without mention of antepartum condition
C0157110|ICD9CM|AB|656.21|Abo isoimmunizat-deliver
C0157111|ICD9CM|PT|656.23|Isoimmunization from other and unspecified blood-group incompatibility, antepartum condition or complication
C0157111|ICD9CM|AB|656.23|Abo isoimmunizat-antepar
C0157112|ICD9CM|PT|656.30|Fetal distress, affecting management of mother, unspecified as to episode of care or not applicable
C0157112|ICD9CM|AB|656.30|Fetal distress-unspec
C0157113|ICD9CM|PT|656.31|Fetal distress, affecting management of mother, delivered, with or without mention of antepartum condition
C0157113|ICD9CM|AB|656.31|Fetal distress-delivered
C0157114|ICD9CM|PT|656.33|Fetal distress, affecting management of mother, antepartum condition or complication
C0157114|ICD9CM|AB|656.33|Fetal distress-antepart
C0157116|ICD9CM|PT|656.40|Intrauterine death, affecting management of mother, unspecified as to episode of care or not applicable
C0157116|ICD9CM|AB|656.40|Intrauterine death-unsp
C0157117|ICD9CM|PT|656.41|Intrauterine death, affecting management of mother, delivered, with or without mention of antepartum condition
C0157117|ICD9CM|AB|656.41|Intrauter death-deliver
C0157118|ICD9CM|PT|656.43|Intrauterine death, affecting management of mother, antepartum condition or complication
C0157118|ICD9CM|AB|656.43|Intrauter death-antepart
C0157119|ICD9CM|HT|656.5|Poor fetal growth affecting management of mother
C0157120|ICD9CM|PT|656.50|Poor fetal growth, affecting management of mother, unspecified as to episode of care or not applicable
C0157120|ICD9CM|AB|656.50|Poor fetal growth-unspec
C0157121|ICD9CM|PT|656.51|Poor fetal growth, affecting management of mother, delivered, with or without mention of antepartum condition
C0157121|ICD9CM|AB|656.51|Poor fetal growth-deliv
C0157122|ICD9CM|PT|656.53|Poor fetal growth, affecting management of mother, antepartum condition or complication
C0157122|ICD9CM|AB|656.53|Poor fetal grth-antepart
C0157123|ICD9CM|HT|656.6|Excessive fetal growth affecting management of mother
C0157124|ICD9CM|PT|656.60|Excessive fetal growth, affecting management of mother, unspecified as to episode of care or not applicable
C0157124|ICD9CM|AB|656.60|Excess fetal grth-unspec
C0157125|ICD9CM|PT|656.61|Excessive fetal growth, affecting management of mother, delivered, with or without mention of antepartum condition
C0157125|ICD9CM|AB|656.61|Excess fetal grth-deliv
C0157126|ICD9CM|PT|656.63|Excessive fetal growth, affecting management of mother, antepartum condition or complication
C0157126|ICD9CM|AB|656.63|Excess fet grth-antepart
C0157127|ICD9CM|PT|656.70|Other placental conditions, affecting management of mother, unspecified as to episode of care or not applicable
C0157127|ICD9CM|AB|656.70|Oth placent cond-unspec
C0157128|ICD9CM|PT|656.71|Other placental conditions, affecting management of mother, delivered, with or without mention of antepartum condition
C0157128|ICD9CM|AB|656.71|Oth placent cond-deliver
C0157129|ICD9CM|PT|656.73|Other placental conditions, affecting management of mother, antepartum condition or complication
C0157129|ICD9CM|AB|656.73|Oth placent cond-antepar
C0157130|ICD9CM|HT|656.8|Other specified fetal and placental problems affecting management of mother
C0157131|ICD9CM|PT|656.80|Other specified fetal and placental problems, affecting management of mother, unspecified as to episode of care or not applicable
C0157131|ICD9CM|AB|656.80|Fet/plac prob NEC-unspec
C0157132|ICD9CM|PT|656.81|Other specified fetal and placental problems, affecting management of mother, delivered, with or without mention of antepartum condition
C0157132|ICD9CM|AB|656.81|Fet/plac prob NEC-deliv
C0157133|ICD9CM|PT|656.83|Other specified fetal and placental problems, affecting management of mother, antepartum condition or complication
C0157133|ICD9CM|AB|656.83|Fet/plac prob NEC-antepa
C0157134|ICD9CM|HT|656.9|Unspecified fetal and placental problem affecting management of mother
C0157135|ICD9CM|PT|656.90|Unspecified fetal and placental problem, affecting management of mother, unspecified as to episode of care or not applicable
C0157135|ICD9CM|AB|656.90|Fet/plac prob NOS-unspec
C0157136|ICD9CM|PT|656.91|Unspecified fetal and placental problem, affecting management of mother, delivered, with or without mention of antepartum condition
C0157136|ICD9CM|AB|656.91|Fet/plac prob NOS-deliv
C0157137|ICD9CM|PT|656.93|Unspecified fetal and placental problem, affecting management of mother, antepartum condition or complication
C0157137|ICD9CM|AB|656.93|Fet/plac prob NOS-antepa
C0157141|ICD9CM|PT|658.00|Oligohydramnios, unspecified as to episode of care or not applicable
C0157141|ICD9CM|AB|658.00|Oligohydramnios-unspec
C0157142|ICD9CM|AB|658.01|Oligohydramnios-deliver
C0157142|ICD9CM|PT|658.01|Oligohydramnios, delivered, with or without mention of antepartum condition
C0157143|ICD9CM|AB|658.03|Oligohydramnios-antepar
C0157143|ICD9CM|PT|658.03|Oligohydramnios, antepartum condition or complication
C0157145|ICD9CM|PT|658.10|Premature rupture of membranes, unspecified as to episode of care or not applicable
C0157145|ICD9CM|AB|658.10|Prem rupt membran-unspec
C0157146|ICD9CM|PT|658.11|Premature rupture of membranes, delivered, with or without mention of antepartum condition
C0157146|ICD9CM|AB|658.11|Prem rupt membran-deliv
C0157147|ICD9CM|AB|658.13|Prem rupt memb-antepart
C0157147|ICD9CM|PT|658.13|Premature rupture of membranes, antepartum condition or complication
C0157149|ICD9CM|PT|658.20|Delayed delivery after spontaneous or unspecified rupture of membranes, unspecified as to episode of care or not applicable
C0157149|ICD9CM|AB|658.20|Prolong rupt memb-unspec
C0157150|ICD9CM|PT|658.21|Delayed delivery after spontaneous or unspecified rupture of membranes, delivered, with or without mention of antepartum condition
C0157150|ICD9CM|AB|658.21|Prolong rupt memb-deliv
C0157151|ICD9CM|PT|658.23|Delayed delivery after spontaneous or unspecified rupture of membranes, antepartum condition or complication
C0157151|ICD9CM|AB|658.23|Prolong rup memb-antepar
C0157152|ICD9CM|HT|658.3|Delayed delivery after artificial rupture of membranes
C0157153|ICD9CM|PT|658.30|Delayed delivery after artificial rupture of membranes, unspecified as to episode of care or not applicable
C0157153|ICD9CM|AB|658.30|Artific rupt membr-unsp
C0157154|ICD9CM|PT|658.31|Delayed delivery after artificial rupture of membranes, delivered, with or without mention of antepartum condition
C0157154|ICD9CM|AB|658.31|Artific rupt membr-deliv
C0157155|ICD9CM|PT|658.33|Delayed delivery after artificial rupture of membranes, antepartum condition or complication
C0157155|ICD9CM|AB|658.33|Artif rupt memb-antepart
C0157157|ICD9CM|PT|658.41|Infection of amniotic cavity, delivered, with or without mention of antepartum condition
C0157157|ICD9CM|AB|658.41|Amniotic infection-deliv
C0157158|ICD9CM|AB|658.43|Amniotic infect-antepart
C0157158|ICD9CM|PT|658.43|Infection of amniotic cavity, antepartum condition or complication
C0157159|ICD9CM|PT|658.80|Other problems associated with amniotic cavity and membranes, unspecified as to episode of care or not applicable
C0157159|ICD9CM|AB|658.80|Amniotic prob NEC-unspec
C0157160|ICD9CM|PT|658.81|Other problems associated with amniotic cavity and membranes, delivered, with or without mention of antepartum condition
C0157160|ICD9CM|AB|658.81|Amniotic prob NEC-deliv
C0157161|ICD9CM|PT|658.83|Other problems associated with amniotic cavity and membranes, antepartum
C0157161|ICD9CM|AB|658.83|Amnion prob NEC-antepart
C0157165|ICD9CM|PT|658.93|Unspecified problem associated with amniotic cavity and membranes, antepartum condition or complication
C0157165|ICD9CM|AB|658.93|Amnion prob NOS-antepart
C0157168|ICD9CM|PT|659.00|Failed mechanical induction of labor, unspecified as to episode of care or not applicable
C0157168|ICD9CM|AB|659.00|Fail mechan induct-unsp
C0157169|ICD9CM|PT|659.01|Failed mechanical induction of labor, delivered, with or without mention of antepartum condition
C0157169|ICD9CM|AB|659.01|Fail mech induct-deliver
C0157170|ICD9CM|PT|659.03|Failed mechanical induction of labor, antepartum condition or complication
C0157170|ICD9CM|AB|659.03|Fail mech induct-antepar
C0157172|ICD9CM|PT|659.10|Failed medical or unspecified induction of labor, unspecified as to episode of care or not applicable
C0157172|ICD9CM|AB|659.10|Fail induction NOS-unsp
C0157173|ICD9CM|PT|659.11|Failed medical or unspecified induction of labor, delivered, with or without mention of antepartum condition
C0157173|ICD9CM|AB|659.11|Fail induction NOS-deliv
C0157174|ICD9CM|PT|659.13|Failed medical or unspecified induction of labor, antepartum condition or complication
C0157174|ICD9CM|AB|659.13|Fail induct NOS-antepart
C0157176|ICD9CM|PT|659.20|Maternal pyrexia during labor, unspecified, unspecified as to episode of care or not applicable
C0157176|ICD9CM|AB|659.20|Pyrexia in labor-unspec
C0157177|ICD9CM|PT|659.21|Maternal pyrexia during labor, unspecified, delivered, with or without mention of antepartum condition
C0157177|ICD9CM|AB|659.21|Pyrexia in labor-deliver
C0157178|ICD9CM|PT|659.23|Maternal pyrexia during labor, unspecified, antepartum condition or complication
C0157178|ICD9CM|AB|659.23|Pyrexia in labor-antepar
C0157179|ICD9CM|HT|659.3|Generalized infection during labor
C0157180|ICD9CM|PT|659.30|Generalized infection during labor, unspecified as to episode of care or not applicable
C0157180|ICD9CM|AB|659.30|Septicemia in labor-unsp
C0157181|ICD9CM|PT|659.31|Generalized infection during labor, delivered, with or without mention of antepartum condition
C0157181|ICD9CM|AB|659.31|Septicem in labor-deliv
C0157182|ICD9CM|PT|659.33|Generalized infection during labor, antepartum condition or complication
C0157182|ICD9CM|AB|659.33|Septicem in labor-antepa
C0157183|ICD9CM|HT|659.4|Grand multiparity, with current pregnancy
C0157184|ICD9CM|PT|659.40|Grand multiparity, unspecified as to episode of care or not applicable
C0157184|ICD9CM|AB|659.40|Grand multiparity-unspec
C0157185|ICD9CM|PT|659.41|Grand multiparity, delivered, with or without mention of antepartum condition
C0157185|ICD9CM|AB|659.41|Grand multiparity-deliv
C0157186|ICD9CM|PT|659.43|Grand multiparity, antepartum condition or complication
C0157186|ICD9CM|AB|659.43|Grand multiparity-antepa
C0157187|ICD9CM|HT|659.5|Elderly primigravida
C0157188|ICD9CM|PT|659.50|Elderly primigravida, unspecified as to episode of care or not applicable
C0157188|ICD9CM|AB|659.50|Elderly primigravid-unsp
C0157189|ICD9CM|PT|659.51|Elderly primigravida, delivered, with or without mention of antepartum condition
C0157189|ICD9CM|AB|659.51|Elderly primigravida-del
C0157190|ICD9CM|AB|659.53|Elder primigravid-antepa
C0157190|ICD9CM|PT|659.53|Elderly primigravida, antepartum condition or complication
C0157191|ICD9CM|HT|659.8|Other specified indications for care or intervention related to labor and delivery
C0157192|ICD9CM|PT|659.80|Other specified indications for care or intervention related to labor and delivery, unspecified as to episode of care or not applicable
C0157192|ICD9CM|AB|659.80|Complic labor NEC-unsp
C0157193|ICD9CM|PT|659.81|Other specified indications for care or intervention related to labor and delivery, delivered, with or without mention of antepartum condition
C0157193|ICD9CM|AB|659.81|Complic labor NEC-deliv
C0157194|ICD9CM|PT|659.83|Other specified indications for care or intervention related to labor and delivery, antepartum condition or complication
C0157194|ICD9CM|AB|659.83|Compl labor NEC-antepart
C0157195|ICD9CM|HT|659.9|Unspecified indication for care or intervention related to labor and delivery
C0157196|ICD9CM|PT|659.90|Unspecified indication for care or intervention related to labor and delivery, unspecified as to episode of care or not applicable
C0157196|ICD9CM|AB|659.90|Complic labor NOS-unsp
C0157197|ICD9CM|PT|659.91|Unspecified indication for care or intervention related to labor and delivery, delivered, with or without mention of antepartum condition
C0157197|ICD9CM|AB|659.91|Complic labor NOS-deliv
C0157198|ICD9CM|PT|659.93|Unspecified indication for care or intervention related to labor and delivery, antepartum condition or complication
C0157198|ICD9CM|AB|659.93|Compl labor NOS-antepart
C0157199|ICD9CM|HT|660.0|Obstruction caused by malposition of fetus at onset of labor
C0157200|ICD9CM|PT|660.00|Obstruction caused by malposition of fetus at onset of labor, unspecified as to episode of care or not applicable
C0157200|ICD9CM|AB|660.00|Obstruct/fet malpos-unsp
C0157201|ICD9CM|PT|660.01|Obstruction caused by malposition of fetus at onset of labor, delivered, with or without mention of antepartum condition
C0157201|ICD9CM|AB|660.01|Obstruc/fet malpos-deliv
C0157202|ICD9CM|PT|660.03|Obstruction caused by malposition of fetus at onset of labor, antepartum condition or complication
C0157202|ICD9CM|AB|660.03|Obstruc/fet malpos-antep
C0157203|ICD9CM|HT|660.1|Obstruction by bony pelvis during labor
C0157204|ICD9CM|PT|660.10|Obstruction by bony pelvis during labor, unspecified as to episode of care or not applicable
C0157204|ICD9CM|AB|660.10|Bony pelv obstruc-unspec
C0157205|ICD9CM|PT|660.11|Obstruction by bony pelvis during labor, delivered, with or without mention of antepartum condition
C0157205|ICD9CM|AB|660.11|Bony pelv obstruct-deliv
C0157206|ICD9CM|PT|660.13|Obstruction by bony pelvis during labor, antepartum condition or complication
C0157206|ICD9CM|AB|660.13|Bony pelv obstruc-antepa
C0157207|ICD9CM|HT|660.2|Obstruction by abnormal pelvic soft tissues during labor
C0157208|ICD9CM|PT|660.20|Obstruction by abnormal pelvic soft tissues during labor, unspecified as to episode of care or not applicable
C0157208|ICD9CM|AB|660.20|Abn pelv tiss obstr-unsp
C0157209|ICD9CM|PT|660.21|Obstruction by abnormal pelvic soft tissues during labor, delivered, with or without mention of antepartum condition
C0157209|ICD9CM|AB|660.21|Abn pelv tis obstr-deliv
C0157210|ICD9CM|PT|660.23|Obstruction by abnormal pelvic soft tissues during labor, antepartum condition or complication
C0157210|ICD9CM|AB|660.23|Abn pelv tis obstr-antep
C0157211|ICD9CM|HT|660.3|Deep transverse arrest and persistent occipitoposterior position during labor and delivery
C0157212|ICD9CM|PT|660.30|Deep transverse arrest and persistent occipitoposterior position, unspecified as to episode of care or not applicable
C0157212|ICD9CM|AB|660.30|Persist occipitpost-unsp
C0157213|ICD9CM|PT|660.31|Deep transverse arrest and persistent occipitoposterior position, delivered, with or without mention of antepartum condition
C0157213|ICD9CM|AB|660.31|Persist occiptpost-deliv
C0157214|ICD9CM|PT|660.33|Deep transverse arrest and persistent occipitoposterior position, antepartum condition or complication
C0157214|ICD9CM|AB|660.33|Persist occiptpost-antep
C0157216|ICD9CM|PT|660.40|Shoulder (girdle) dystocia, unspecified as to episode of care or not applicable
C0157216|ICD9CM|AB|660.40|Shoulder dystocia-unspec
C0157218|ICD9CM|PT|660.43|Shoulder (girdle) dystocia, antepartum condition or complication
C0157218|ICD9CM|AB|660.43|Shoulder dystocia-antepa
C0157220|ICD9CM|AB|660.50|Locked twins-unspecified
C0157220|ICD9CM|PT|660.50|Locked twins, unspecified as to episode of care or not applicable
C0157221|ICD9CM|AB|660.51|Locked twins-delivered
C0157221|ICD9CM|PT|660.51|Locked twins, delivered, with or without mention of antepartum condition
C0157222|ICD9CM|AB|660.53|Locked twins-antepartum
C0157222|ICD9CM|PT|660.53|Locked twins, antepartum condition or complication
C0157223|ICD9CM|HT|660.6|Failed trial of labor, unspecified
C0157224|ICD9CM|PT|660.60|Unspecified failed trial of labor, unspecified as to episode of care or not applicable
C0157224|ICD9CM|AB|660.60|Fail trial lab NOS-unsp
C0157225|ICD9CM|PT|660.61|Unspecified failed trial of labor, delivered, with or without mention of antepartum condition
C0157225|ICD9CM|AB|660.61|Fail trial lab NOS-deliv
C0157226|ICD9CM|PT|660.63|Unspecified failed trial of labor, antepartum condition or complication
C0157226|ICD9CM|AB|660.63|Fail trial lab NOS-antep
C0157228|ICD9CM|PT|660.70|Failed forceps or vacuum extractor, unspecified, unspecified as to episode of care or not applicable
C0157228|ICD9CM|AB|660.70|Failed forcep NOS-unspec
C0157229|ICD9CM|PT|660.71|Failed forceps or vacuum extractor, unspecified, delivered, with or without mention of antepartum condition
C0157229|ICD9CM|AB|660.71|Failed forceps NOS-deliv
C0157230|ICD9CM|PT|660.73|Failed forceps or vacuum extractor, unspecified, antepartum condition or complication
C0157230|ICD9CM|AB|660.73|Fail forceps NOS-antepar
C0157231|ICD9CM|HT|660.8|Other causes of obstructed labor
C0157232|ICD9CM|PT|660.80|Other causes of obstructed labor, unspecified as to episode of care or not applicable
C0157232|ICD9CM|AB|660.80|Obstruc labor NEC-unspec
C0157233|ICD9CM|PT|660.81|Other causes of obstructed labor, delivered, with or without mention of antepartum condition
C0157233|ICD9CM|AB|660.81|Obstruct labor NEC-deliv
C0157234|ICD9CM|PT|660.83|Other causes of obstructed labor, antepartum condition or complication
C0157234|ICD9CM|AB|660.83|Obstruc labor NEC-antepa
C0157235|ICD9CM|PT|660.90|Unspecified obstructed labor, unspecified as to episode of care or not applicable
C0157235|ICD9CM|AB|660.90|Obstruc labor NOS-unspec
C0157236|ICD9CM|PT|660.91|Unspecified obstructed labor, delivered, with or without mention of antepartum condition
C0157236|ICD9CM|AB|660.91|Obstruct labor NOS-deliv
C0157237|ICD9CM|PT|660.93|Unspecified obstructed labor, antepartum condition or complication
C0157237|ICD9CM|AB|660.93|Obstruc labor NOS-antepa
C0157239|ICD9CM|PT|661.00|Primary uterine inertia, unspecified as to episode of care or not applicable
C0157239|ICD9CM|AB|661.00|Prim uterine inert-unsp
C0157240|ICD9CM|PT|661.01|Primary uterine inertia, delivered, with or without mention of antepartum condition
C0157240|ICD9CM|AB|661.01|Prim uterine inert-deliv
C0157241|ICD9CM|AB|661.03|Prim uter inert-antepart
C0157241|ICD9CM|PT|661.03|Primary uterine inertia, antepartum condition or complication
C0157242|ICD9CM|PT|661.10|Secondary uterine inertia, unspecified as to episode of care or not applicable
C0157242|ICD9CM|AB|661.10|Sec uterine inert-unspec
C0157243|ICD9CM|PT|661.11|Secondary uterine inertia, delivered, with or without mention of antepartum condition
C0157243|ICD9CM|AB|661.11|Sec uterine inert-deliv
C0157244|ICD9CM|AB|661.13|Sec uterine inert-antepa
C0157244|ICD9CM|PT|661.13|Secondary uterine inertia, antepartum condition or complication
C0157246|ICD9CM|PT|661.21|Other and unspecified uterine inertia, delivered, with or without mention of antepartum condition
C0157246|ICD9CM|AB|661.21|Uterine inert NEC-deliv
C0157247|ICD9CM|PT|661.23|Other and unspecified uterine inertia, antepartum condition or complication
C0157247|ICD9CM|AB|661.23|Uterine inert NEC-antepa
C0157248|ICD9CM|PT|661.30|Precipitate labor, unspecified as to episode of care or not applicable
C0157248|ICD9CM|AB|661.30|Precipitate labor-unspec
C0157249|ICD9CM|PT|661.31|Precipitate labor, delivered, with or without mention of antepartum condition
C0157249|ICD9CM|AB|661.31|Precipitate labor-deliv
C0157250|ICD9CM|AB|661.33|Precipitate labor-antepa
C0157250|ICD9CM|PT|661.33|Precipitate labor, antepartum condition or complication
C0157252|ICD9CM|PT|661.40|Hypertonic, incoordinate, or prolonged uterine contractions, unspecified as to episode of care or not applicable
C0157252|ICD9CM|AB|661.40|Uter dystocia NOS-unspec
C0157253|ICD9CM|PT|661.41|Hypertonic, incoordinate, or prolonged uterine contractions, delivered, with or without mention of antepartum condition
C0157253|ICD9CM|AB|661.41|Uter dystocia NOS-deliv
C0157254|ICD9CM|PT|661.43|Hypertonic, incoordinate, or prolonged uterine contractions, antepartum condition or complication
C0157254|ICD9CM|AB|661.43|Uter dystocia NOS-antepa
C0157256|ICD9CM|AB|661.90|Abnormal labor NOS-unsp
C0157256|ICD9CM|PT|661.90|Unspecified abnormality of labor, unspecified as to episode of care or not applicable
C0157258|ICD9CM|PT|661.93|Unspecified abnormality of labor, antepartum condition or complication
C0157258|ICD9CM|AB|661.93|Abnorm labor NOS-antepar
C0157259|ICD9CM|HT|662.0|Prolonged first stage of labor
C0157260|ICD9CM|PT|662.00|Prolonged first stage of labor, unspecified as to episode of care or not applicable
C0157260|ICD9CM|AB|662.00|Prolonged 1st stage-unsp
C0157261|ICD9CM|PT|662.01|Prolonged first stage of labor, delivered, with or without mention of antepartum condition
C0157261|ICD9CM|AB|662.01|Prolong 1st stage-deliv
C0157262|ICD9CM|AB|662.03|Prolong 1st stage-antepa
C0157262|ICD9CM|PT|662.03|Prolonged first stage of labor, antepartum condition or complication
C0157263|ICD9CM|PT|662.10|Unspecified prolonged labor, unspecified as to episode of care or not applicable
C0157263|ICD9CM|AB|662.10|Prolonged labor NOS-unsp
C0157264|ICD9CM|PT|662.11|Unspecified prolonged labor, delivered, with or without mention of antepartum condition
C0157264|ICD9CM|AB|662.11|Prolong labor NOS-deliv
C0157265|ICD9CM|PT|662.13|Unspecified prolonged labor, antepartum condition or complication
C0157265|ICD9CM|AB|662.13|Prolong labor NOS-antepa
C0157266|ICD9CM|HT|662.2|Prolonged second stage of labor
C0157267|ICD9CM|PT|662.20|Prolonged second stage of labor, unspecified as to episode of care or not applicable
C0157267|ICD9CM|AB|662.20|Prolonged 2nd stage-unsp
C0157268|ICD9CM|PT|662.21|Prolonged second stage of labor, delivered, with or without mention of antepartum condition
C0157268|ICD9CM|AB|662.21|Prolong 2nd stage-deliv
C0157269|ICD9CM|AB|662.23|Prolong 2nd stage-antepa
C0157269|ICD9CM|PT|662.23|Prolonged second stage of labor, antepartum condition or complication
C0157270|ICD9CM|HT|662.3|Delayed delivery of second twin, triplet, etc.
C0157270|ICD9CM|PT|662.33|Delayed delivery of second twin, triplet, etc., antepartum condition or complication
C0157270|ICD9CM|AB|662.33|Delay del 2 twin-antepar
C0157271|ICD9CM|PT|662.30|Delayed delivery of second twin, triplet, etc., unspecified as to episode of care or not applicable
C0157271|ICD9CM|AB|662.30|Delay del 2nd twin-unsp
C0157272|ICD9CM|PT|662.31|Delayed delivery of second twin, triplet, etc., delivered, with or without mention of antepartum condition
C0157272|ICD9CM|AB|662.31|Delay del 2nd twin-deliv
C0157275|ICD9CM|HT|663.0|Prolapse of cord complicating labor and delivery
C0157275|ICD9CM|PT|663.00|Prolapse of cord complicating labor and delivery, unspecified as to episode of care or not applicable
C0157275|ICD9CM|AB|663.00|Cord prolapse-unspec
C0157277|ICD9CM|AB|663.01|Cord prolapse-delivered
C0157277|ICD9CM|PT|663.01|Prolapse of cord complicating labor and delivery, delivered, with or without mention of antepartum condition
C0157278|ICD9CM|PT|663.03|Prolapse of cord complicating labor and delivery, antepartum condition or complication
C0157278|ICD9CM|AB|663.03|Cord prolapse-antepartum
C0157280|ICD9CM|PT|663.10|Cord around neck with compression, complicating labor and delivery, unspecified as to episode of care or not applicable
C0157280|ICD9CM|AB|663.10|Cord around neck-unspec
C0157281|ICD9CM|PT|663.11|Cord around neck, with compression, complicating labor and delivery, delivered, with or without mention of antepartum condition
C0157281|ICD9CM|AB|663.11|Cord around neck-deliver
C0157282|ICD9CM|PT|663.13|Cord around neck, with compression, complicating labor and delivery, antepartum condition or complication
C0157282|ICD9CM|AB|663.13|Cord around neck-antepar
C0157283|ICD9CM|HT|663.2|Other and unspecified cord entanglement, with compression, complicating labor and delivery
C0157284|ICD9CM|PT|663.20|Other and unspecified cord entanglement, with compression, complicating labor and delivery, unspecified as to episode of care or not applicable
C0157284|ICD9CM|AB|663.20|Cord compress NEC-unspec
C0157285|ICD9CM|PT|663.21|Other and unspecified cord entanglement, with compression, complicating labor and delivery, delivered, with or without mention of antepartum condition
C0157285|ICD9CM|AB|663.21|Cord compress NEC-deliv
C0157286|ICD9CM|PT|663.23|Other and unspecified cord entanglement, with compression, complicating labor and delivery, antepartum condition or complication
C0157286|ICD9CM|AB|663.23|Cord compres NEC-antepar
C0157287|ICD9CM|HT|663.3|Other and unspecified cord entanglement, without mention of compression, complicating labor and delivery
C0157288|ICD9CM|PT|663.30|Other and unspecified cord entanglement, without mention of compression, complicating labor and delivery, unspecified as to episode of care or not applicable
C0157288|ICD9CM|AB|663.30|Cord entangle NEC-unspec
C0157289|ICD9CM|PT|663.31|Other and unspecified cord entanglement, without mention of compression, complicating labor and delivery, delivered, with or without mention of antepartum condition
C0157289|ICD9CM|AB|663.31|Cord entangle NEC-deliv
C0157290|ICD9CM|PT|663.33|Other and unspecified cord entanglement, without mention of compression, complicating labor and delivery, antepartum condition or complication
C0157290|ICD9CM|AB|663.33|Cord entangl NEC-antepar
C0157291|ICD9CM|HT|663.4|Short cord complicating labor and delivery
C0157292|ICD9CM|AB|663.40|Short cord-unspecified
C0157292|ICD9CM|PT|663.40|Short cord complicating labor and delivery, unspecified as to episode of care or not applicable
C0157293|ICD9CM|AB|663.41|Short cord-delivered
C0157293|ICD9CM|PT|663.41|Short cord complicating labor and delivery, delivered, with or without mention of antepartum condition
C0157294|ICD9CM|PT|663.43|Short cord complicating labor and delivery, antepartum condition or complication
C0157294|ICD9CM|AB|663.43|Short cord-antepartum
C0157297|ICD9CM|PT|663.51|Vasa previa complicating labor and delivery, delivered, with or without mention of antepartum condition
C0157297|ICD9CM|AB|663.51|Vasa previa-delivered
C0157299|ICD9CM|HT|663.6|Vascular lesions of cord complicating labor and delivery
C0157300|ICD9CM|PT|663.60|Vascular lesions of cord complicating labor and delivery, unspecified as to episode of care or not applicable
C0157300|ICD9CM|AB|663.60|Vasc lesion cord-unspec
C0157301|ICD9CM|PT|663.61|Vascular lesions of cord complicating labor and delivery, delivered, with or without mention of antepartum condition
C0157301|ICD9CM|AB|663.61|Vasc lesion cord-deliver
C0157302|ICD9CM|PT|663.63|Vascular lesions of cord complicating labor and delivery, antepartum condition or complication
C0157302|ICD9CM|AB|663.63|Vasc lesion cord-antepar
C0157303|ICD9CM|HT|663.8|Other umbilical cord complications during labor and delivery
C0157304|ICD9CM|PT|663.80|Other umbilical cord complications complicating labor and delivery, unspecified as to episode of care or not applicable
C0157304|ICD9CM|AB|663.80|Cord complicat NEC-unsp
C0157305|ICD9CM|PT|663.81|Other umbilical cord complications complicating labor and delivery, delivered, with or without mention of antepartum condition
C0157305|ICD9CM|AB|663.81|Cord complicat NEC-deliv
C0157306|ICD9CM|PT|663.83|Other umbilical cord complications complicating labor and delivery, antepartum condition or complication
C0157306|ICD9CM|AB|663.83|Cord compl NEC-antepart
C0157307|ICD9CM|HT|663|Umbilical cord complications during labor and delivery
C0157307|ICD9CM|HT|663.9|Unspecified umbilical cord complication during labor and delivery
C0157308|ICD9CM|PT|663.90|Unspecified umbilical cord complication complicating labor and delivery, unspecified as to episode of care or not applicable
C0157308|ICD9CM|AB|663.90|Cord complicat NOS-unsp
C0157309|ICD9CM|PT|663.91|Unspecified umbilical cord complication complicating labor and delivery, delivered, with or without mention of antepartum condition
C0157309|ICD9CM|AB|663.91|Cord complicat NOS-deliv
C0157310|ICD9CM|PT|663.93|Unspecified umbilical cord complication complicating labor and delivery, antepartum condition or complication
C0157310|ICD9CM|AB|663.93|Cord compl NOS-antepart
C0157311|ICD9CM|HT|664|Trauma to perineum and vulva during delivery
C0157313|ICD9CM|PT|664.00|First-degree perineal laceration, unspecified as to episode of care or not applicable
C0157313|ICD9CM|AB|664.00|Del w 1 deg lacerat-unsp
C0157315|ICD9CM|PT|664.04|First-degree perineal laceration, postpartum condition or complication
C0157315|ICD9CM|AB|664.04|Del w 1 deg lac-postpart
C0157317|ICD9CM|PT|664.10|Second-degree perineal laceration, unspecified as to episode of care or not applicable
C0157317|ICD9CM|AB|664.10|Del w 2 deg lacerat-unsp
C0157321|ICD9CM|PT|664.20|Third-degree perineal laceration, unspecified as to episode of care or not applicable
C0157321|ICD9CM|AB|664.20|Del w 3 deg lacerat-unsp
C0157323|ICD9CM|PT|664.24|Third-degree perineal laceration, postpartum condition or complication
C0157323|ICD9CM|AB|664.24|Del w 3 deg lac-postpart
C0157325|ICD9CM|PT|664.30|Fourth-degree perineal laceration, unspecified as to episode of care or not applicable
C0157325|ICD9CM|AB|664.30|Del w 4 deg lacerat-unsp
C0157327|ICD9CM|PT|664.34|Fourth-degree perineal laceration, postpartum condition or complication
C0157327|ICD9CM|AB|664.34|Del w 4 deg lac-postpart
C0157329|ICD9CM|PT|664.40|Unspecified perineal laceration, unspecified as to episode of care or not applicable
C0157329|ICD9CM|AB|664.40|Ob perineal lac NOS-unsp
C0157331|ICD9CM|PT|664.44|Unspecified perineal laceration, postpartum condition or complication
C0157331|ICD9CM|AB|664.44|Perineal lac NOS-postpar
C0157332|ICD9CM|HT|664.5|Vulvar and perineal hematoma during delivery
C0157333|ICD9CM|PT|664.50|Vulvar and perineal hematoma, unspecified as to episode of care or not applicable
C0157333|ICD9CM|AB|664.50|Ob perineal hematom-unsp
C0157334|ICD9CM|PT|664.51|Vulvar and perineal hematoma, delivered, with or without mention of antepartum condition
C0157334|ICD9CM|AB|664.51|Ob perineal hematoma-del
C0157335|ICD9CM|PT|664.54|Vulvar and perineal hematoma, postpartum condition or complication
C0157335|ICD9CM|AB|664.54|Perin hematoma-postpart
C0157336|ICD9CM|HT|664.8|Other specified trauma to perineum and vulva during delivery
C0157337|ICD9CM|PT|664.80|Other specified trauma to perineum and vulva, unspecified as to episode of care or not applicable
C0157337|ICD9CM|AB|664.80|Ob perin traum NEC-unsp
C0157338|ICD9CM|PT|664.81|Other specified trauma to perineum and vulva, delivered, with or without mention of antepartum condition
C0157338|ICD9CM|AB|664.81|Ob perineal trau NEC-del
C0157339|ICD9CM|PT|664.84|Other specified trauma to perineum and vulva, postpartum condition or complication
C0157339|ICD9CM|AB|664.84|Perin traum NEC-postpart
C0157340|ICD9CM|HT|664.9|Unspecified trauma to perineum and vulva during delivery
C0157341|ICD9CM|PT|664.90|Unspecified trauma to perineum and vulva, unspecified as to episode of care or not applicable
C0157341|ICD9CM|AB|664.90|Ob perin traum NOS-unsp
C0157342|ICD9CM|PT|664.91|Unspecified trauma to perineum and vulva, delivered, with or without mention of antepartum condition
C0157342|ICD9CM|AB|664.91|Ob perineal trau NOS-del
C0157343|ICD9CM|PT|664.94|Unspecified trauma to perineum and vulva, postpartum condition or complication
C0157343|ICD9CM|AB|664.94|Perin traum NOS-postpart
C0157344|ICD9CM|HT|665|Other obstetrical trauma
C0157345|ICD9CM|HT|665.0|Rupture of uterus before onset of labor
C0157346|ICD9CM|PT|665.00|Rupture of uterus before onset of labor, unspecified as to episode of care or not applicable
C0157346|ICD9CM|AB|665.00|Prelabor rupt uter-unsp
C0157347|ICD9CM|PT|665.01|Rupture of uterus before onset of labor, delivered, with or without mention of antepartum condition
C0157347|ICD9CM|AB|665.01|Prelabor rupt uterus-del
C0157350|ICD9CM|PT|665.10|Rupture of uterus during labor, unspecified as to episode of care or not applicable
C0157350|ICD9CM|AB|665.10|Rupture uterus NOS-unsp
C0157351|ICD9CM|PT|665.11|Rupture of uterus during labor, delivered, with or without mention of antepartum condition
C0157351|ICD9CM|AB|665.11|Rupture uterus NOS-deliv
C0157355|ICD9CM|PT|665.20|Inversion of uterus, unspecified as to episode of care or not applicable
C0157355|ICD9CM|AB|665.20|Inversion of uterus-unsp
C0157356|ICD9CM|PT|665.22|Inversion of uterus, delivered, with mention of postpartum complication
C0157356|ICD9CM|AB|665.22|Invers uterus-del w p/p
C0157357|ICD9CM|PT|665.24|Inversion of uterus, postpartum condition or complication
C0157357|ICD9CM|AB|665.24|Invers uterus-postpart
C0157358|ICD9CM|HT|665.3|Obstetrical laceration of cervix
C0157358|ICD9CM|PT|665.31|Laceration of cervix, delivered, with or without mention of antepartum condition
C0157358|ICD9CM|AB|665.31|Lacerat of cervix-deliv
C0157359|ICD9CM|PT|665.30|Laceration of cervix, unspecified as to episode of care or not applicable
C0157359|ICD9CM|AB|665.30|Lacerat of cervix-unspec
C0157361|ICD9CM|PT|665.34|Laceration of cervix, postpartum condition or complication
C0157361|ICD9CM|AB|665.34|Lacer of cervix-postpart
C0157362|ICD9CM|HT|665.4|High vaginal laceration during and after labor
C0157363|ICD9CM|PT|665.40|High vaginal laceration, unspecified as to episode of care or not applicable
C0157363|ICD9CM|AB|665.40|High vaginal lacer-unsp
C0157364|ICD9CM|PT|665.41|High vaginal laceration, delivered, with or without mention of antepartum condition
C0157364|ICD9CM|AB|665.41|High vaginal lacer-deliv
C0157365|ICD9CM|PT|665.44|High vaginal laceration, postpartum condition or complication
C0157365|ICD9CM|AB|665.44|High vaginal lac-postpar
C0157366|ICD9CM|HT|665.5|Other obstetrical injury to pelvic organs
C0157367|ICD9CM|PT|665.50|Other injury to pelvic organs, unspecified as to episode of care or not applicable
C0157367|ICD9CM|AB|665.50|Ob inj pelv org NEC-unsp
C0157368|ICD9CM|PT|665.51|Other injury to pelvic organs, delivered, with or without mention of antepartum condition
C0157368|ICD9CM|AB|665.51|Ob inj pelv org NEC-del
C0157369|ICD9CM|PT|665.54|Other injury to pelvic organs, postpartum condition or complication
C0157369|ICD9CM|AB|665.54|Inj pelv org NEC-postpar
C0157371|ICD9CM|PT|665.60|Damage to pelvic joints and ligaments, unspecified as to episode of care or not applicable
C0157371|ICD9CM|AB|665.60|Damage to pelvic jt-unsp
C0157373|ICD9CM|PT|665.64|Damage to pelvic joints and ligaments, postpartum condition or complication
C0157373|ICD9CM|AB|665.64|Damage pelvic jt-postpar
C0157375|ICD9CM|PT|665.70|Pelvic hematoma, unspecified as to episode of care or not applicable
C0157375|ICD9CM|AB|665.70|Ob pelvic hematoma-unsp
C0157377|ICD9CM|PT|665.72|Pelvic hematoma, delivered with mention of postpartum complication
C0157377|ICD9CM|AB|665.72|Pelvic hematom-del w pp
C0157378|ICD9CM|PT|665.74|Pelvic hematoma, postpartum condition or complication
C0157378|ICD9CM|AB|665.74|Pelvic hematoma-postpart
C0157379|ICD9CM|HT|665.8|Other specified obstetrical trauma
C0157380|ICD9CM|PT|665.80|Other specified obstetrical trauma, unspecified as to episode of care or not applicable
C0157380|ICD9CM|AB|665.80|Ob trauma NEC-unspec
C0157381|ICD9CM|PT|665.81|Other specified obstetrical trauma, delivered, with or without mention of antepartum condition
C0157381|ICD9CM|AB|665.81|Ob trauma NEC-delivered
C0157382|ICD9CM|PT|665.82|Other specified obstetrical trauma, delivered, with mention of postpartum complication
C0157382|ICD9CM|AB|665.82|Ob trauma NEC-del w p/p
C0157383|ICD9CM|PT|665.83|Other specified obstetrical trauma, antepartum condition or complication
C0157383|ICD9CM|AB|665.83|Ob trauma NEC-antepartum
C0157384|ICD9CM|PT|665.84|Other specified obstetrical trauma, postpartum condition or complication
C0157384|ICD9CM|AB|665.84|Ob trauma NEC-postpartum
C0157386|ICD9CM|PT|665.90|Unspecified obstetrical trauma, unspecified as to episode of care or not applicable
C0157386|ICD9CM|AB|665.90|Ob trauma NOS-unspec
C0157387|ICD9CM|PT|665.91|Unspecified obstetrical trauma, delivered, with or without mention of antepartum condition
C0157387|ICD9CM|AB|665.91|Ob trauma NOS-delivered
C0157388|ICD9CM|PT|665.92|Unspecified obstetrical trauma, delivered, with mention of postpartum complication
C0157388|ICD9CM|AB|665.92|Ob trauma NOS-del w p/p
C0157389|ICD9CM|PT|665.93|Unspecified obstetrical trauma, antepartum condition or complication
C0157389|ICD9CM|AB|665.93|Ob trauma NOS-antepartum
C0157390|ICD9CM|PT|665.94|Unspecified obstetrical trauma, postpartum condition or complication
C0157390|ICD9CM|AB|665.94|Ob trauma NOS-postpartum
C0157392|ICD9CM|PT|666.00|Third-stage postpartum hemorrhage, unspecified as to episode of care or not applicable
C0157392|ICD9CM|AB|666.00|Third-stage hem-unspec
C0157393|ICD9CM|PT|666.02|Third-stage postpartum hemorrhage, delivered, with mention of postpartum complication
C0157393|ICD9CM|AB|666.02|Thrd-stage hem-del w p/p
C0157394|ICD9CM|PT|666.10|Other immediate postpartum hemorrhage, unspecified as to episode of care or not applicable
C0157394|ICD9CM|AB|666.10|Postpartum hem NEC-unsp
C0157395|ICD9CM|PT|666.12|Other immediate postpartum hemorrhage, delivered, with mention of postpartum complication
C0157395|ICD9CM|AB|666.12|Postpa hem NEC-del w p/p
C0157398|ICD9CM|PT|666.22|Delayed and secondary postpartum hemorrhage, delivered, with mention of postpartum complication
C0157398|ICD9CM|AB|666.22|Delay p/p hem-del w p/p
C0157401|ICD9CM|PT|666.30|Postpartum coagulation defects, unspecified as to episode of care or not applicable
C0157401|ICD9CM|AB|666.30|Postpart coagul def-unsp
C0157402|ICD9CM|PT|666.32|Postpartum coagulation defects, delivered, with mention of postpartum complication
C0157402|ICD9CM|AB|666.32|P/p coag def-del w p/p
C0157403|ICD9CM|HT|666.3|Postpartum coagulation defects
C0157403|ICD9CM|AB|666.34|Postpart coag def-postpa
C0157403|ICD9CM|PT|666.34|Postpartum coagulation defects, postpartum condition or complication
C0157404|ICD9CM|HT|667|Retained placenta or membranes, without hemorrhage
C0157405|ICD9CM|PT|667.00|Retained placenta without hemorrhage, unspecified as to episode of care or not applicable
C0157405|ICD9CM|AB|667.00|Retain placenta NOS-unsp
C0157406|ICD9CM|PT|667.02|Retained placenta without hemorrhage, delivered, with mention of postpartum complication
C0157406|ICD9CM|AB|667.02|Retnd plac NOS-del w p/p
C0157407|ICD9CM|PT|667.04|Retained placenta without hemorrhage, postpartum condition or complication
C0157407|ICD9CM|AB|667.04|Retain plac NOS-postpart
C0157408|ICD9CM|HT|667.1|Retained portions of placenta or membranes, without hemorrhage
C0157409|ICD9CM|PT|667.10|Retained portions of placenta or membranes, without hemorrhage, unspecified as to episode of care or not applicable
C0157409|ICD9CM|AB|667.10|Retain prod concept-unsp
C0157410|ICD9CM|PT|667.12|Retained portions of placenta or membranes, without hemorrhage, delivered, with mention of postpartum complication
C0157410|ICD9CM|AB|667.12|Ret prod conc-del w p/p
C0157411|ICD9CM|PT|667.14|Retained portions of placenta or membranes, without hemorrhage, postpartum condition or complication
C0157411|ICD9CM|AB|667.14|Ret prod concept-postpar
C0157412|ICD9CM|HT|668|Complications of the administration of anesthetic or other sedation in labor and delivery
C0157413|ICD9CM|HT|668.0|Pulmonary complications of anesthesia or other sedation in labor and delivery
C0157414|ICD9CM|PT|668.00|Pulmonary complications of anesthesia or other sedation in labor and delivery, unspecified as to episode of care or not applicable
C0157414|ICD9CM|AB|668.00|Pulm compl in del-unspec
C0157415|ICD9CM|PT|668.01|Pulmonary complications of anesthesia or other sedation in labor and delivery, delivered, with or without mention of antepartum condition
C0157415|ICD9CM|AB|668.01|Pulm compl in del-deliv
C0157416|ICD9CM|PT|668.02|Pulmonary complications of anesthesia or other sedation in labor and delivery, delivered, with mention of postpartum complication
C0157416|ICD9CM|AB|668.02|Pulm complic-del w p/p
C0157417|ICD9CM|PT|668.03|Pulmonary complications of anesthesia or other sedation in labor and delivery, antepartum condition or complication
C0157417|ICD9CM|AB|668.03|Pulm complicat-antepart
C0157418|ICD9CM|PT|668.04|Pulmonary complications of anesthesia or other sedation in labor and delivery, postpartum condition or complication
C0157418|ICD9CM|AB|668.04|Pulm complicat-postpart
C0157420|ICD9CM|PT|668.10|Cardiac complications of anesthesia or other sedation in labor and delivery, unspecified as to episode of care or not applicable
C0157420|ICD9CM|AB|668.10|Heart compl in del-unsp
C0157421|ICD9CM|PT|668.11|Cardiac complications of anesthesia or other sedation in labor and delivery, delivered, with or without mention of antepartum condition
C0157421|ICD9CM|AB|668.11|Heart compl in del-deliv
C0157422|ICD9CM|PT|668.12|Cardiac complications of anesthesia or other sedation in labor and delivery, delivered, with mention of postpartum complication
C0157422|ICD9CM|AB|668.12|Heart compl-del w p/p
C0157423|ICD9CM|PT|668.13|Cardiac complications of anesthesia or other sedation in labor and delivery, antepartum condition or complication
C0157423|ICD9CM|AB|668.13|Heart complic-antepart
C0157424|ICD9CM|PT|668.14|Cardiac complications of anesthesia or other sedation in labor and delivery, postpartum condition or complication
C0157424|ICD9CM|AB|668.14|Heart complic-postpart
C0157425|ICD9CM|HT|668.2|Central nervous system complications of anesthesia or other sedation in labor and delivery
C0157426|ICD9CM|PT|668.20|Central nervous system complications of anesthesia or other sedation in labor and delivery, unspecified as to episode of care or not applicable
C0157426|ICD9CM|AB|668.20|Cns compl labor/del-unsp
C0157427|ICD9CM|PT|668.21|Central nervous system complications of anesthesia or other sedation in labor and delivery, delivered, with or without mention of antepartum condition
C0157427|ICD9CM|AB|668.21|Cns compl lab/del-deliv
C0157428|ICD9CM|PT|668.22|Central nervous system complications of anesthesia or other sedation in labor and delivery, delivered, with mention of postpartum complication
C0157428|ICD9CM|AB|668.22|Cns complic-del w p/p
C0157429|ICD9CM|PT|668.23|Central nervous system complications of anesthesia or other sedation in labor and delivery, antepartum condition or complication
C0157429|ICD9CM|AB|668.23|Cns compl in del-antepar
C0157430|ICD9CM|PT|668.24|Central nervous system complications of anesthesia or other sedation in labor and delivery, postpartum condition or complication
C0157430|ICD9CM|AB|668.24|Cns compl in del-postpar
C0157431|ICD9CM|HT|668.8|Other complications of anesthesia or other sedation in labor and delivery
C0157432|ICD9CM|PT|668.80|Other complications of anesthesia or other sedation in labor and delivery, unspecified as to episode of care or not applicable
C0157432|ICD9CM|AB|668.80|Anesth comp del NEC-unsp
C0157434|ICD9CM|PT|668.82|Other complications of anesthesia or other sedation in labor and delivery, delivered, with mention of postpartum complication
C0157434|ICD9CM|AB|668.82|Anesth compl NEC-del p/p
C0157435|ICD9CM|PT|668.83|Other complications of anesthesia or other sedation in labor and delivery, antepartum condition or complication
C0157435|ICD9CM|AB|668.83|Anesth compl antepartum
C0157436|ICD9CM|PT|668.84|Other complications of anesthesia or other sedation in labor and delivery, postpartum condition or complication
C0157436|ICD9CM|PT|668.81|Other complications of anesthesia or other sedation in labor and delivery, delivered, with or without mention of antepartum condition
C0157436|ICD9CM|AB|668.81|Anesth compl NEC-deliver
C0157436|ICD9CM|AB|668.84|Anesth compl-postpartum
C0157437|ICD9CM|HT|668.9|Unspecified complication of anesthesia or other sedation in labor and delivery
C0157438|ICD9CM|PT|668.90|Unspecified complication of anesthesia and other sedation in labor and delivery, unspecified as to episode of care or not applicable
C0157438|ICD9CM|AB|668.90|Anesth comp del NOS-unsp
C0157439|ICD9CM|PT|668.91|Unspecified complication of anesthesia and other sedation in labor and delivery, delivered, with or without mention of antepartum condition
C0157439|ICD9CM|AB|668.91|Anesth compl NOS-deliver
C0157440|ICD9CM|PT|668.92|Unspecified complication of anesthesia and other sedation in labor and delivery, delivered, with mention of postpartum complication
C0157440|ICD9CM|AB|668.92|Anesth compl NOS-del p/p
C0157441|ICD9CM|PT|668.93|Unspecified complication of anesthesia and other sedation in labor and delivery, antepartum condition or complication
C0157441|ICD9CM|AB|668.93|Anesth compl-antepartum
C0157442|ICD9CM|PT|668.94|Unspecified complication of anesthesia and other sedation in labor and delivery, postpartum condition or complication
C0157442|ICD9CM|AB|668.94|Anesth compl-postpartum
C0157443|ICD9CM|HT|669.8|Other complications of labor and delivery
C0157445|ICD9CM|PT|669.00|Maternal distress complicating labor and delivery, unspecified as to episode of care or not applicable
C0157445|ICD9CM|AB|669.00|Maternal distress-unspec
C0157446|ICD9CM|PT|669.01|Maternal distress complicating labor and delivery, delivered, with or without mention of antepartum condition
C0157446|ICD9CM|AB|669.01|Maternal distress-deliv
C0157447|ICD9CM|PT|669.02|Maternal distress complicating labor and delivery, delivered, with mention of postpartum complication
C0157447|ICD9CM|AB|669.02|Matern distres-del w p/p
C0157448|ICD9CM|PT|669.03|Maternal distress complicating labor and delivery, antepartum condition or complication
C0157448|ICD9CM|AB|669.03|Matern distress-antepar
C0157449|ICD9CM|PT|669.04|Maternal distress complicating labor and delivery, postpartum condition or complication
C0157449|ICD9CM|AB|669.04|Matern distress-postpart
C0157450|ICD9CM|HT|669.1|Shock during or following labor and delivery
C0157451|ICD9CM|PT|669.10|Shock during or following labor and delivery, unspecified as to episode of care or not applicable
C0157451|ICD9CM|AB|669.10|Obstetric shock-unspec
C0157452|ICD9CM|PT|669.11|Shock during or following labor and delivery, delivered, with or without mention of antepartum condition
C0157452|ICD9CM|AB|669.11|Obstetric shock-deliver
C0157453|ICD9CM|PT|669.12|Shock during or following labor and delivery, delivered, with mention of postpartum complication
C0157453|ICD9CM|AB|669.12|Obstet shock-deliv w p/p
C0157454|ICD9CM|PT|669.13|Shock during or following labor and delivery, antepartum condition or complication
C0157454|ICD9CM|AB|669.13|Obstetric shock-antepar
C0157455|ICD9CM|PT|669.14|Shock during or following labor and delivery, postpartum condition or complication
C0157455|ICD9CM|AB|669.14|Obstetric shock-postpart
C0157456|ICD9CM|PT|669.20|Maternal hypotension syndrome, unspecified as to episode of care or not applicable
C0157456|ICD9CM|AB|669.20|Matern hypotens syn-unsp
C0157457|ICD9CM|PT|669.21|Maternal hypotension syndrome, delivered, with or without mention of antepartum condition
C0157457|ICD9CM|AB|669.21|Matern hypoten syn-deliv
C0157458|ICD9CM|PT|669.22|Maternal hypotension syndrome, delivered, with mention of postpartum complication
C0157458|ICD9CM|AB|669.22|Matern hypoten-del w p/p
C0157459|ICD9CM|AB|669.23|Matern hypotens-antepar
C0157459|ICD9CM|PT|669.23|Maternal hypotension syndrome, antepartum condition or complication
C0157460|ICD9CM|AB|669.24|Matern hypotens-postpart
C0157460|ICD9CM|PT|669.24|Maternal hypotension syndrome, postpartum condition or complication
C0157462|ICD9CM|PT|669.30|Acute kidney failure following labor and delivery, unspecified as to episode of care or not applicable
C0157462|ICD9CM|AB|669.30|Ac kidny fail w del-unsp
C0157463|ICD9CM|PT|669.32|Acute kidney failure following labor and delivery, delivered, with mention of postpartum complication
C0157463|ICD9CM|AB|669.32|Ac kidney fail-del w p/p
C0157464|ICD9CM|PT|669.34|Acute kidney failure following labor and delivery, postpartum condition or complication
C0157464|ICD9CM|AB|669.34|Ac kidney fail-postpart
C0157465|ICD9CM|HT|669.4|Other complications of obstetrical surgery and procedures
C0157466|ICD9CM|PT|669.40|Other complications of obstetrical surgery and procedures, unspecified as to episode of care or not applicable
C0157466|ICD9CM|AB|669.40|Oth ob surg compl-unspec
C0157467|ICD9CM|PT|669.41|Other complications of obstetrical surgery and procedures, delivered, with or without mention of antepartum condition
C0157467|ICD9CM|AB|669.41|Oth ob compl-delivered
C0157468|ICD9CM|PT|669.42|Other complications of obstetrical surgery and procedures, delivered, with mention of postpartum complication
C0157468|ICD9CM|AB|669.42|Oth ob compl-deliv w p/p
C0157469|ICD9CM|PT|669.44|Other complications of obstetrical surgery and procedures, postpartum condition or complication
C0157469|ICD9CM|AB|669.44|Oth ob surg compl-postpa
C0157470|ICD9CM|HT|669.5|Forceps or vacuum extractor delivery without mention of indication
C0157471|ICD9CM|PT|669.50|Forceps or vacuum extractor delivery without mention of indication, unspecified as to episode of care or not applicable
C0157471|ICD9CM|AB|669.50|Forcep deliv NOS-unspec
C0157472|ICD9CM|PT|669.51|Forceps or vacuum extractor delivery without mention of indication, delivered, with or without mention of antepartum condition
C0157472|ICD9CM|AB|669.51|Forcep deliv NOS-deliver
C0157474|ICD9CM|PT|669.60|Breech extraction, without mention of indication, unspecified as to episode of care or not applicable
C0157474|ICD9CM|AB|669.60|Breech extr NOS-unspec
C0157475|ICD9CM|PT|669.61|Breech extraction, without mention of indication, delivered, with or without mention of antepartum condition
C0157475|ICD9CM|AB|669.61|Breech extr NOS-deliver
C0157477|ICD9CM|PT|669.70|Cesarean delivery, without mention of indication, unspecified as to episode of care or not applicable
C0157477|ICD9CM|AB|669.70|Cesarean deliv NOS-unsp
C0157478|ICD9CM|PT|669.71|Cesarean delivery, without mention of indication, delivered, with or without mention of antepartum condition
C0157478|ICD9CM|AB|669.71|Cesarean delivery NOS
C0157479|ICD9CM|PT|669.80|Other complications of labor and delivery, unspecified as to episode of care or not applicable
C0157479|ICD9CM|AB|669.80|Compl lab/deliv NEC-unsp
C0157480|ICD9CM|PT|669.81|Other complications of labor and delivery, delivered, with or without mention of antepartum condition
C0157480|ICD9CM|AB|669.81|Comp lab/deliv NEC-deliv
C0157481|ICD9CM|PT|669.82|Other complications of labor and delivery, delivered, with mention of postpartum complication
C0157481|ICD9CM|AB|669.82|Compl del NEC-del w p/p
C0157482|ICD9CM|PT|669.83|Other complications of labor and delivery, antepartum condition or complication
C0157482|ICD9CM|AB|669.83|Compl deliv NEC-antepar
C0157483|ICD9CM|PT|669.84|Other complications of labor and delivery, postpartum condition or complication
C0157483|ICD9CM|AB|669.84|Compl deliv NEC-postpart
C0157484|ICD9CM|PT|669.90|Unspecified complication of labor and delivery, unspecified as to episode of care or not applicable
C0157484|ICD9CM|AB|669.90|Compl lab/deliv NOS-unsp
C0157485|ICD9CM|PT|669.91|Unspecified complication of labor and delivery, delivered, with or without mention of antepartum condition
C0157485|ICD9CM|AB|669.91|Comp lab/deliv NOS-deliv
C0157486|ICD9CM|PT|669.92|Unspecified complication of labor and delivery, delivered, with mention of postpartum complication
C0157486|ICD9CM|AB|669.92|Compl del NOS-del w p/p
C0157487|ICD9CM|PT|669.93|Unspecified complication of labor and delivery, antepartum condition or complication
C0157487|ICD9CM|AB|669.93|Compl deliv NOS-antepar
C0157488|ICD9CM|PT|669.94|Unspecified complication of labor and delivery, postpartum condition or complication
C0157488|ICD9CM|AB|669.94|Compl deliv NOS-postpart
C0157489|ICD9CM|HT|670|Major puerperal infection
C0157489|ICD9CM|HT|670.0|Major puerperal infection, unspecified
C0157491|ICD9CM|PT|670.02|Major puerperal infection, delivered, with mention of postpartum complication
C0157491|ICD9CM|AB|670.02|Maj puer inf NOS-del p/p
C0157495|ICD9CM|PT|671.00|Varicose veins of legs complicating pregnancy and the puerperium, unspecified as to episode of care or not applicable
C0157495|ICD9CM|AB|671.00|Varic vein leg preg-unsp
C0157496|ICD9CM|PT|671.01|Varicose veins of legs complicating pregnancy and the puerperium, delivered, with or without mention of antepartum condition
C0157496|ICD9CM|AB|671.01|Varicose vein leg-deliv
C0157497|ICD9CM|PT|671.02|Varicose veins of legs complicating pregnancy and the puerperium, delivered, with mention of postpartum complication
C0157497|ICD9CM|AB|671.02|Varic vein leg-del w p/p
C0157498|ICD9CM|PT|671.03|Varicose veins of legs complicating pregnancy and the puerperium, antepartum condition or complication
C0157498|ICD9CM|AB|671.03|Varic vein leg-antepart
C0157499|ICD9CM|PT|671.04|Varicose veins of legs complicating pregnancy and the puerperium, postpartum condition or complication
C0157499|ICD9CM|AB|671.04|Varic vein leg-postpart
C0157501|ICD9CM|PT|671.10|Varicose veins of vulva and perineum complicating pregnancy and the puerperium, unspecified as to episode of care or not applicable
C0157501|ICD9CM|AB|671.10|Varic vulva preg-unspec
C0157502|ICD9CM|PT|671.11|Varicose veins of vulva and perineum complicating pregnancy and the puerperium, delivered, with or without mention of antepartum condition
C0157502|ICD9CM|AB|671.11|Varicose vulva-delivered
C0157503|ICD9CM|PT|671.12|Varicose veins of vulva and perineum complicating pregnancy and the puerperium, delivered, with mention of postpartum complication
C0157503|ICD9CM|AB|671.12|Varicose vulva-del w p/p
C0157504|ICD9CM|PT|671.13|Varicose veins of vulva and perineum complicating pregnancy and the puerperium, antepartum condition or complication
C0157504|ICD9CM|AB|671.13|Varicose vulva-antepart
C0157505|ICD9CM|PT|671.14|Varicose veins of vulva and perineum complicating pregnancy and the puerperium, postpartum condition or complication
C0157505|ICD9CM|AB|671.14|Varicose vulva-postpart
C0157508|ICD9CM|PT|671.21|Superficial thrombophlebitis complicating pregnancy and the puerperium, delivered, with or without mention of antepartum condition
C0157508|ICD9CM|AB|671.21|Thrombophlebitis-deliver
C0157509|ICD9CM|PT|671.22|Superficial thrombophlebitis complicating pregnancy and the puerperium, delivered, with mention of postpartum complication
C0157509|ICD9CM|AB|671.22|Thrombophleb-deliv w p/p
C0157514|ICD9CM|PT|671.31|Deep phlebothrombosis, antepartum, delivered, with or without mention of antepartum condition
C0157514|ICD9CM|AB|671.31|Deep throm antepar-deliv
C0157516|ICD9CM|PT|671.40|Deep phlebothrombosis, postpartum, unspecified as to episode of care or not applicable
C0157516|ICD9CM|AB|671.40|Deep thromb postpar-unsp
C0157517|ICD9CM|PT|671.42|Deep phlebothrombosis, postpartum, delivered, with mention of postpartum complication
C0157517|ICD9CM|AB|671.42|Thromb postpar-del w p/p
C0157519|ICD9CM|PT|671.50|Other phlebitis and thrombosis complicating pregnancy and the puerperium, unspecified as to episode of care or not applicable
C0157519|ICD9CM|AB|671.50|Thrombosis NEC preg-unsp
C0157520|ICD9CM|PT|671.51|Other phlebitis and thrombosis complicating pregnancy and the puerperium, delivered, with or without mention of antepartum condition
C0157520|ICD9CM|AB|671.51|Thrombosis NEC-delivered
C0157521|ICD9CM|PT|671.52|Other phlebitis and thrombosis complicating pregnancy and the puerperium, delivered, with mention of postpartum complication
C0157521|ICD9CM|AB|671.52|Thromb NEC-deliv w p/p
C0157522|ICD9CM|PT|671.53|Other phlebitis and thrombosis complicating pregnancy and the puerperium, antepartum condition or complication
C0157522|ICD9CM|AB|671.53|Thrombosis NEC-antepart
C0157523|ICD9CM|PT|671.54|Other phlebitis and thrombosis complicating pregnancy and the puerperium, postpartum condition or complication
C0157523|ICD9CM|AB|671.54|Thrombosis NEC-postpart
C0157524|ICD9CM|HT|671.8|Other venous complications in pregnancy and the puerperium
C0157525|ICD9CM|PT|671.80|Other venous complications of pregnancy and the puerperium, unspecified as to episode of care or not applicable
C0157525|ICD9CM|AB|671.80|Ven compl preg NEC-unsp
C0157526|ICD9CM|PT|671.81|Other venous complications of pregnancy and the puerperium, delivered, with or without mention of antepartum condition
C0157526|ICD9CM|AB|671.81|Venous compl NEC-deliver
C0157527|ICD9CM|PT|671.82|Other venous complications of pregnancy and the puerperium, delivered, with mention of postpartum complication
C0157527|ICD9CM|AB|671.82|Ven comp NEC-deliv w p/p
C0157532|ICD9CM|PT|671.91|Unspecified venous complication of pregnancy and the puerperium, delivered, with or without mention of antepartum condition
C0157532|ICD9CM|AB|671.91|Venous compl NOS-deliver
C0157533|ICD9CM|PT|671.92|Unspecified venous complication of pregnancy and the puerperium, delivered, with mention of postpartum complication
C0157533|ICD9CM|AB|671.92|Ven comp NOS-deliv w p/p
C0157535|ICD9CM|PT|671.94|Unspecified venous complication of pregnancy and the puerperium, postpartum condition or complication
C0157535|ICD9CM|AB|671.94|Venous compl NOS-postpar
C0157536|ICD9CM|HT|672.0|Pyrexia of unknown origin during the puerperium
C0157536|ICD9CM|HT|672|Pyrexia of unknown origin during the puerperium
C0157540|ICD9CM|HT|673|Obstetrical pulmonary embolism
C0157541|ICD9CM|HT|673.0|Obstetrical air embolism
C0157542|ICD9CM|PT|673.00|Obstetrical air embolism, unspecified as to episode of care or not applicable
C0157542|ICD9CM|AB|673.00|Ob air embolism-unspec
C0157543|ICD9CM|PT|673.01|Obstetrical air embolism, delivered, with or without mention of antepartum condition
C0157543|ICD9CM|AB|673.01|Ob air embolism-deliver
C0157544|ICD9CM|PT|673.02|Obstetrical air embolism, delivered, with mention of postpartum complication
C0157544|ICD9CM|AB|673.02|Ob air embol-deliv w p/p
C0157545|ICD9CM|PT|673.03|Obstetrical air embolism, antepartum condition or complication
C0157545|ICD9CM|AB|673.03|Ob air embolism-antepart
C0157546|ICD9CM|PT|673.04|Obstetrical air embolism, postpartum condition or complication
C0157546|ICD9CM|AB|673.04|Ob air embolism-postpart
C0157548|ICD9CM|PT|673.11|Amniotic fluid embolism, delivered, with or without mention of antepartum condition
C0157548|ICD9CM|AB|673.11|Amniotic embolism-deliv
C0157549|ICD9CM|PT|673.12|Amniotic fluid embolism, delivered, with mention of postpartum complication
C0157549|ICD9CM|AB|673.12|Amniot embol-deliv w p/p
C0157550|ICD9CM|PT|673.13|Amniotic fluid embolism, antepartum condition or complication
C0157550|ICD9CM|AB|673.13|Amniotic embol-antepart
C0157551|ICD9CM|PT|673.14|Amniotic fluid embolism, postpartum condition or complication
C0157551|ICD9CM|AB|673.14|Amniotic embol-postpart
C0157552|ICD9CM|HT|673.2|Obstetrical blood-clot embolism
C0157552|ICD9CM|PT|673.20|Obstetrical blood-clot embolism, unspecified as to episode of care or not applicable
C0157552|ICD9CM|AB|673.20|Ob pulm embol NOS-unspec
C0157554|ICD9CM|PT|673.21|Obstetrical blood-clot embolism, delivered, with or without mention of antepartum condition
C0157554|ICD9CM|AB|673.21|Pulm embol NOS-delivered
C0157555|ICD9CM|PT|673.22|Obstetrical blood-clot embolism, delivered, with mention of postpartum complication
C0157555|ICD9CM|AB|673.22|Pulm embol NOS-del w p/p
C0157556|ICD9CM|PT|673.23|Obstetrical blood-clot embolism, antepartum condition or complication
C0157556|ICD9CM|AB|673.23|Pulm embol NOS-antepart
C0157557|ICD9CM|PT|673.24|Obstetrical blood-clot embolism, postpartum condition or complication
C0157557|ICD9CM|AB|673.24|Pulm embol NOS-postpart
C0157560|ICD9CM|PT|673.31|Obstetrical pyemic and septic embolism, delivered, with or without mention of antepartum condition
C0157560|ICD9CM|AB|673.31|Ob pyemic embol-deliver
C0157561|ICD9CM|PT|673.32|Obstetrical pyemic and septic embolism, delivered, with mention of postpartum complication
C0157561|ICD9CM|AB|673.32|Ob pyem embol-del w p/p
C0157562|ICD9CM|PT|673.33|Obstetrical pyemic and septic embolism, antepartum condition or complication
C0157562|ICD9CM|AB|673.33|Ob pyemic embol-antepart
C0157563|ICD9CM|PT|673.34|Obstetrical pyemic and septic embolism, postpartum condition or complication
C0157563|ICD9CM|AB|673.34|Ob pyemic embol-postpart
C0157564|ICD9CM|HT|673.8|Other obstetrical pulmonary embolism
C0157565|ICD9CM|PT|673.80|Other obstetrical pulmonary embolism, unspecified as to episode of care or not applicable
C0157565|ICD9CM|AB|673.80|Ob pulmon embol NEC-unsp
C0157566|ICD9CM|PT|673.81|Other obstetrical pulmonary embolism, delivered, with or without mention of antepartum condition
C0157566|ICD9CM|AB|673.81|Pulmon embol NEC-deliver
C0157567|ICD9CM|PT|673.82|Other obstetrical pulmonary embolism, delivered, with mention of postpartum complication
C0157567|ICD9CM|AB|673.82|Pulm embol NEC-del w p/p
C0157568|ICD9CM|PT|673.83|Other obstetrical pulmonary embolism, antepartum condition or complication
C0157568|ICD9CM|AB|673.83|Pulmon embol NEC-antepar
C0157569|ICD9CM|PT|673.84|Other obstetrical pulmonary embolism, postpartum condition or complication
C0157569|ICD9CM|AB|673.84|Pulmon embol NEC-postpar
C0157571|ICD9CM|HT|674.0|Cerebrovascular disorders in the puerperium
C0157572|ICD9CM|PT|674.00|Cerebrovascular disorders in the puerperium, unspecified as to episode of care or not applicable
C0157572|ICD9CM|AB|674.00|Puerp cerebvasc dis-unsp
C0157573|ICD9CM|PT|674.01|Cerebrovascular disorders in the puerperium, delivered, with or without mention of antepartum condition
C0157573|ICD9CM|AB|674.01|Puerp cerebvas dis-deliv
C0157574|ICD9CM|PT|674.02|Cerebrovascular disorders in the puerperium, delivered, with mention of postpartum complication
C0157574|ICD9CM|AB|674.02|Cerebvas dis-deliv w p/p
C0157575|ICD9CM|PT|674.03|Cerebrovascular disorders in the puerperium, antepartum condition or complication
C0157575|ICD9CM|AB|674.03|Cerebrovasc dis-antepart
C0157578|ICD9CM|PT|674.10|Disruption of cesarean wound, unspecified as to episode of care or not applicable
C0157578|ICD9CM|AB|674.10|Disrupt c-sect wnd-unsp
C0157579|ICD9CM|PT|674.12|Disruption of cesarean wound, delivered, with mention of postpartum complication
C0157579|ICD9CM|AB|674.12|Disrupt c-sect-del w p/p
C0157582|ICD9CM|PT|674.20|Disruption of perineal wound, unspecified as to episode of care or not applicable
C0157582|ICD9CM|AB|674.20|Disrupt perineum-unspec
C0157583|ICD9CM|PT|674.22|Disruption of perineal wound, delivered, with mention of postpartum complication
C0157583|ICD9CM|AB|674.22|Disrupt perin-del w p/p
C0157585|ICD9CM|HT|674.3|Other complications of obstetrical surgical wounds
C0157586|ICD9CM|PT|674.30|Other complications of obstetrical surgical wounds, unspecified as to episode of care or not applicable
C0157586|ICD9CM|AB|674.30|Ob surg compl NEC-unspec
C0157587|ICD9CM|PT|674.32|Other complications of obstetrical surgical wounds, delivered, with mention of postpartum complication
C0157587|ICD9CM|AB|674.32|Ob surg compl-del w p/p
C0157588|ICD9CM|PT|674.34|Other complications of obstetrical surgical wounds, postpartum condition or complication
C0157588|ICD9CM|AB|674.34|Ob surg comp NEC-postpar
C0157589|ICD9CM|PT|674.40|Placental polyp, unspecified as to episode of care or not applicable
C0157589|ICD9CM|AB|674.40|Placental polyp-unspec
C0157590|ICD9CM|PT|674.42|Placental polyp, delivered, with mention of postpartum complication
C0157590|ICD9CM|AB|674.42|Placent polyp-del w p/p
C0157591|ICD9CM|AB|674.44|Placental polyp-postpart
C0157591|ICD9CM|PT|674.44|Placental polyp, postpartum condition or complication
C0157592|ICD9CM|HT|674.8|Other complications of the puerperium
C0157594|ICD9CM|PT|674.82|Other complications of puerperium, delivered, with mention of postpartum complication
C0157594|ICD9CM|AB|674.82|Puerp comp NEC-del w p/p
C0157597|ICD9CM|PT|674.92|Unspecified complications of puerperium, delivered, with mention of postpartum complication
C0157597|ICD9CM|AB|674.92|Puerp comp NOS-del w p/p
C0157600|ICD9CM|PT|675.00|Infections of nipple associated with childbirth, unspecified as to episode of care or not applicable
C0157600|ICD9CM|AB|675.00|Infect nipple preg-unsp
C0157601|ICD9CM|PT|675.01|Infections of nipple associated with childbirth, delivered, with or without mention of antepartum condition
C0157601|ICD9CM|AB|675.01|Infect nipple-delivered
C0157602|ICD9CM|PT|675.02|Infections of nipple associated with childbirth, delivered, with mention of postpartum complication
C0157602|ICD9CM|AB|675.02|Infect nipple-del w p/p
C0157603|ICD9CM|PT|675.03|Infections of nipple associated with childbirth, antepartum condition or complication
C0157603|ICD9CM|AB|675.03|Infect nipple-antepartum
C0157604|ICD9CM|PT|675.04|Infections of nipple associated with childbirth, postpartum condition or complication
C0157604|ICD9CM|AB|675.04|Infect nipple-postpartum
C0157606|ICD9CM|PT|675.10|Abscess of breast associated with childbirth, unspecified as to episode of care or not applicable
C0157606|ICD9CM|AB|675.10|Breast abscess preg-unsp
C0157607|ICD9CM|PT|675.11|Abscess of breast associated with childbirth, delivered, with or without mention of antepartum condition
C0157607|ICD9CM|AB|675.11|Breast abscess-delivered
C0157608|ICD9CM|PT|675.12|Abscess of breast associated with childbirth, delivered, with mention of postpartum complication
C0157608|ICD9CM|AB|675.12|Breast abscess-del w p/p
C0157611|ICD9CM|HT|675.2|Nonpurulent mastitis associated with childbirth
C0157612|ICD9CM|PT|675.20|Nonpurulent mastitis associated with childbirth, unspecified as to episode of care or not applicable
C0157612|ICD9CM|AB|675.20|Mastitis in preg-unspec
C0157613|ICD9CM|PT|675.21|Nonpurulent mastitis associated with childbirth, delivered, with or without mention of antepartum condition
C0157613|ICD9CM|AB|675.21|Mastitis-delivered
C0157614|ICD9CM|PT|675.22|Nonpurulent mastitis associated with childbirth, delivered, with mention of postpartum complication
C0157614|ICD9CM|AB|675.22|Mastitis-deliv w p/p
C0157617|ICD9CM|HT|675.8|Other specified infections of the breast and nipple associated with childbirth
C0157618|ICD9CM|PT|675.80|Other specified infections of the breast and nipple associated with childbirth, unspecified as to episode of care or not applicable
C0157618|ICD9CM|AB|675.80|Breast inf preg NEC-unsp
C0157619|ICD9CM|PT|675.81|Other specified infections of the breast and nipple associated with childbirth, delivered, with or without mention of antepartum condition
C0157619|ICD9CM|AB|675.81|Breast infect NEC-deliv
C0157620|ICD9CM|PT|675.82|Other specified infections of the breast and nipple associated with childbirth, delivered, with mention of postpartum complication
C0157620|ICD9CM|AB|675.82|Breast inf NEC-del w p/p
C0157621|ICD9CM|PT|675.83|Other specified infections of the breast and nipple associated with childbirth, antepartum condition or complication
C0157621|ICD9CM|AB|675.83|Breast inf NEC-antepart
C0157622|ICD9CM|PT|675.84|Other specified infections of the breast and nipple associated with childbirth, postpartum condition or complication
C0157622|ICD9CM|AB|675.84|Breast inf NEC-postpart
C0157623|ICD9CM|HT|675.9|Unspecified infection of the breast and nipple associated with childbirth
C0157623|ICD9CM|HT|675|Infections of the breast and nipple associated with childbirth
C0157624|ICD9CM|PT|675.90|Unspecified infection of the breast and nipple associated with childbirth, unspecified as to episode of care or not applicable
C0157624|ICD9CM|AB|675.90|Breast inf preg NOS-unsp
C0157625|ICD9CM|PT|675.91|Unspecified infection of the breast and nipple associated with childbirth, delivered, with or without mention of antepartum condition
C0157625|ICD9CM|AB|675.91|Breast infect NOS-deliv
C0157626|ICD9CM|PT|675.92|Unspecified infection of the breast and nipple associated with childbirth, delivered, with mention of postpartum complication
C0157626|ICD9CM|AB|675.92|Breast inf NOS-del w p/p
C0157627|ICD9CM|PT|675.93|Unspecified infection of the breast and nipple associated with childbirth, antepartum condition or complication
C0157627|ICD9CM|AB|675.93|Breast inf NOS-antepart
C0157628|ICD9CM|PT|675.94|Unspecified infection of the breast and nipple associated with childbirth, postpartum condition or complication
C0157628|ICD9CM|AB|675.94|Breast inf NOS-postpart
C0157629|ICD9CM|HT|676|Other disorders of the breast associated with childbirth and disorders of lactation
C0157630|ICD9CM|HT|676.0|Retracted nipple associated with childbirth
C0157631|ICD9CM|PT|676.00|Retracted nipple associated with childbirth, unspecified as to episode of care or not applicable
C0157631|ICD9CM|AB|676.00|Retract nipple preg-unsp
C0157632|ICD9CM|PT|676.01|Retracted nipple associated with childbirth, delivered, with or without mention of antepartum condition
C0157632|ICD9CM|AB|676.01|Retracted nipple-deliver
C0157633|ICD9CM|PT|676.02|Retracted nipple associated with childbirth, delivered, with mention of postpartum complication
C0157633|ICD9CM|AB|676.02|Retract nipple-del w p/p
C0157634|ICD9CM|PT|676.03|Retracted nipple associated with childbirth, antepartum condition or complication
C0157634|ICD9CM|AB|676.03|Retract nipple-antepart
C0157635|ICD9CM|PT|676.04|Retracted nipple associated with childbirth, postpartum condition or complication
C0157635|ICD9CM|AB|676.04|Retract nipple-postpart
C0157636|ICD9CM|HT|676.1|Cracked nipple associated with childbirth
C0157637|ICD9CM|PT|676.10|Cracked nipple associated with childbirth, unspecified as to episode of care or not applicable
C0157637|ICD9CM|AB|676.10|Cracked nipple preg-unsp
C0157638|ICD9CM|PT|676.11|Cracked nipple associated with childbirth, delivered, with or without mention of antepartum condition
C0157638|ICD9CM|AB|676.11|Cracked nipple-delivered
C0157639|ICD9CM|PT|676.12|Cracked nipple associated with childbirth, delivered, with mention of postpartum complication
C0157639|ICD9CM|AB|676.12|Cracked nipple-del w p/p
C0157640|ICD9CM|PT|676.13|Cracked nipple associated with childbirth, antepartum condition or complication
C0157640|ICD9CM|AB|676.13|Cracked nipple-antepart
C0157641|ICD9CM|PT|676.14|Cracked nipple associated with childbirth, postpartum condition or complication
C0157641|ICD9CM|AB|676.14|Cracked nipple-postpart
C0157642|ICD9CM|HT|676.2|Engorgement of breasts associated with childbirth
C0157643|ICD9CM|PT|676.20|Engorgement of breasts associated with childbirth, unspecified as to episode of care or not applicable
C0157643|ICD9CM|AB|676.20|Breast engorge-unspec
C0157644|ICD9CM|PT|676.21|Engorgement of breasts associated with childbirth, delivered, with or without mention of antepartum condition
C0157644|ICD9CM|AB|676.21|Breast engorge-delivered
C0157645|ICD9CM|PT|676.22|Engorgement of breasts associated with childbirth, delivered, with mention of postpartum complication
C0157645|ICD9CM|AB|676.22|Breast engorge-del w p/p
C0157646|ICD9CM|PT|676.23|Engorgement of breasts associated with childbirth, antepartum condition or complication
C0157646|ICD9CM|AB|676.23|Breast engorge-antepart
C0157647|ICD9CM|PT|676.24|Engorgement of breasts associated with childbirth, postpartum condition or complication
C0157647|ICD9CM|AB|676.24|Breast engorge-postpart
C0157648|ICD9CM|HT|676.3|Other and unspecified disorder of breast associated with childbirth
C0157649|ICD9CM|PT|676.30|Other and unspecified disorder of breast associated with childbirth, unspecified as to episode of care or not applicable
C0157649|ICD9CM|AB|676.30|Breast dis preg NEC-unsp
C0157650|ICD9CM|PT|676.31|Other and unspecified disorder of breast associated with childbirth, delivered, with or without mention of antepartum condition
C0157650|ICD9CM|AB|676.31|Breast dis NEC-delivered
C0157651|ICD9CM|PT|676.32|Other and unspecified disorder of breast associated with childbirth, delivered, with mention of postpartum complication
C0157651|ICD9CM|AB|676.32|Breast dis NEC-del w p/p
C0157652|ICD9CM|PT|676.33|Other and unspecified disorder of breast associated with childbirth, antepartum condition or complication
C0157652|ICD9CM|AB|676.33|Breast dis NEC-antepart
C0157653|ICD9CM|PT|676.34|Other and unspecified disorder of breast associated with childbirth, postpartum condition or complication
C0157653|ICD9CM|AB|676.34|Breast dis NEC-postpart
C0157655|ICD9CM|PT|676.41|Failure of lactation, delivered, with or without mention of antepartum condition
C0157655|ICD9CM|AB|676.41|Lactation fail-delivered
C0157656|ICD9CM|PT|676.44|Failure of lactation, postpartum condition or complication
C0157656|ICD9CM|PT|676.42|Failure of lactation, delivered, with mention of postpartum complication
C0157656|ICD9CM|AB|676.44|Lactation fail-postpart
C0157656|ICD9CM|AB|676.42|Lactation fail-del w p/p
C0157657|ICD9CM|PT|676.43|Failure of lactation, antepartum condition or complication
C0157657|ICD9CM|AB|676.43|Lactation fail-antepart
C0157660|ICD9CM|PT|676.51|Suppressed lactation, delivered, with or without mention of antepartum condition
C0157660|ICD9CM|AB|676.51|Suppr lactation-deliver
C0157661|ICD9CM|PT|676.54|Suppressed lactation, postpartum condition or complication
C0157661|ICD9CM|PT|676.52|Suppressed lactation, delivered, with mention of postpartum complication
C0157661|ICD9CM|AB|676.52|Suppr lactat-del w p/p
C0157661|ICD9CM|AB|676.54|Suppr lactation-postpart
C0157662|ICD9CM|PT|676.53|Suppressed lactation, antepartum condition or complication
C0157662|ICD9CM|AB|676.53|Suppr lactation-antepar
C0157665|ICD9CM|AB|676.61|Galactorrhea-delivered
C0157665|ICD9CM|PT|676.61|Galactorrhea associated with childbirth, delivered, with or without mention of antepartum condition
C0157666|ICD9CM|PT|676.62|Galactorrhea associated with childbirth, delivered, with mention of postpartum complication
C0157666|ICD9CM|AB|676.62|Galactorrhea-del w p/p
C0157667|ICD9CM|PT|676.63|Galactorrhea associated with childbirth, antepartum condition or complication
C0157667|ICD9CM|AB|676.63|Galactorrhea-antepartum
C0157668|ICD9CM|PT|676.64|Galactorrhea associated with childbirth, postpartum condition or complication
C0157668|ICD9CM|AB|676.64|Galactorrhea-postpartum
C0157669|ICD9CM|HT|676.8|Other disorders of lactation
C0157669|ICD9CM|PT|676.80|Other disorders of lactation, unspecified as to episode of care or not applicable
C0157669|ICD9CM|AB|676.80|Lactation dis NEC-unspec
C0157671|ICD9CM|PT|676.81|Other disorders of lactation, delivered, with or without mention of antepartum condition
C0157671|ICD9CM|AB|676.81|Lactation dis NEC-deliv
C0157672|ICD9CM|PT|676.84|Other disorders of lactation, postpartum condition or complication
C0157672|ICD9CM|PT|676.82|Other disorders of lactation, delivered, with mention of postpartum complication
C0157672|ICD9CM|AB|676.84|Lactat dis NEC-postpart
C0157672|ICD9CM|AB|676.82|Lactat dis NEC-del w p/p
C0157673|ICD9CM|PT|676.83|Other disorders of lactation, antepartum condition or complication
C0157673|ICD9CM|AB|676.83|Lactat dis NEC-antepart
C0157676|ICD9CM|PT|676.91|Unspecified disorder of lactation, delivered, with or without mention of antepartum condition
C0157676|ICD9CM|AB|676.91|Lactation dis NOS-deliv
C0157677|ICD9CM|PT|676.92|Unspecified disorder of lactation, delivered, with mention of postpartum complication
C0157677|ICD9CM|AB|676.92|Lactat dis NOS-del w p/p
C0157678|ICD9CM|PT|676.93|Unspecified disorder of lactation, antepartum condition or complication
C0157678|ICD9CM|AB|676.93|Lactat dis NOS-antepart
C0157679|ICD9CM|PT|676.94|Unspecified disorder of lactation, postpartum condition or complication
C0157679|ICD9CM|AB|676.94|Lactat dis NOS-postpart
C0157680|ICD9CM|HT|680|Carbuncle and furuncle
C0157681|ICD9CM|PT|680.0|Carbuncle and furuncle of face
C0157681|ICD9CM|AB|680.0|Carbuncle of face
C0157682|ICD9CM|PT|680.1|Carbuncle and furuncle of neck
C0157682|ICD9CM|AB|680.1|Carbuncle of neck
C0157683|ICD9CM|PT|680.2|Carbuncle and furuncle of trunk
C0157683|ICD9CM|AB|680.2|Carbuncle of trunk
C0157684|ICD9CM|PT|680.3|Carbuncle and furuncle of upper arm and forearm
C0157684|ICD9CM|AB|680.3|Carbuncle of arm
C0157685|ICD9CM|PT|680.4|Carbuncle and furuncle of hand
C0157685|ICD9CM|AB|680.4|Carbuncle of hand
C0157686|ICD9CM|PT|680.5|Carbuncle and furuncle of buttock
C0157686|ICD9CM|AB|680.5|Carbuncle of buttock
C0157687|ICD9CM|PT|680.6|Carbuncle and furuncle of leg, except foot
C0157687|ICD9CM|AB|680.6|Carbuncle of leg
C0157688|ICD9CM|PT|680.7|Carbuncle and furuncle of foot
C0157688|ICD9CM|AB|680.7|Carbuncle of foot
C0157689|ICD9CM|PT|680.8|Carbuncle and furuncle of other specified sites
C0157689|ICD9CM|AB|680.8|Carbuncle, site NEC
C0157690|ICD9CM|HT|681|Cellulitis and abscess of finger and toe
C0157691|ICD9CM|HT|681.0|Cellulitis and abscess of finger
C0157691|ICD9CM|AB|681.00|Cellulitis, finger NOS
C0157691|ICD9CM|PT|681.00|Cellulitis and abscess of finger, unspecified
C0157692|ICD9CM|PT|681.02|Onychia and paronychia of finger
C0157692|ICD9CM|AB|681.02|Onychia of finger
C0157693|ICD9CM|HT|681.1|Cellulitis and abscess of toe
C0157693|ICD9CM|AB|681.10|Cellulitis, toe NOS
C0157693|ICD9CM|PT|681.10|Cellulitis and abscess of toe, unspecified
C0157694|ICD9CM|PT|681.11|Onychia and paronychia of toe
C0157694|ICD9CM|AB|681.11|Onychia of toe
C0157695|ICD9CM|HT|682|Other cellulitis and abscess
C0157696|ICD9CM|PT|682.0|Cellulitis and abscess of face
C0157696|ICD9CM|AB|682.0|Cellulitis of face
C0157697|ICD9CM|PT|682.1|Cellulitis and abscess of neck
C0157697|ICD9CM|AB|682.1|Cellulitis of neck
C0157698|ICD9CM|PT|682.2|Cellulitis and abscess of trunk
C0157698|ICD9CM|AB|682.2|Cellulitis of trunk
C0157699|ICD9CM|PT|682.3|Cellulitis and abscess of upper arm and forearm
C0157699|ICD9CM|AB|682.3|Cellulitis of arm
C0157701|ICD9CM|PT|682.5|Cellulitis and abscess of buttock
C0157701|ICD9CM|AB|682.5|Cellulitis of buttock
C0157702|ICD9CM|PT|682.6|Cellulitis and abscess of leg, except foot
C0157702|ICD9CM|AB|682.6|Cellulitis of leg
C0157704|ICD9CM|PT|682.8|Cellulitis and abscess of other specified sites
C0157704|ICD9CM|AB|682.8|Cellulitis, site NEC
C0157705|ICD9CM|AB|683|Acute lymphadenitis
C0157705|ICD9CM|PT|683|Acute lymphadenitis
C0157707|ICD9CM|HT|686|Other local infections of skin and subcutaneous tissue
C0157708|ICD9CM|PT|692.0|Contact dermatitis and other eczema due to detergents
C0157708|ICD9CM|AB|692.0|Detergent dermatitis
C0157709|ICD9CM|PT|692.1|Contact dermatitis and other eczema due to oils and greases
C0157709|ICD9CM|AB|692.1|Oil & grease dermatitis
C0157710|ICD9CM|PT|692.2|Contact dermatitis and other eczema due to solvents
C0157710|ICD9CM|AB|692.2|Solvent dermatitis
C0157711|ICD9CM|PT|692.3|Contact dermatitis and other eczema due to drugs and medicines in contact with skin
C0157711|ICD9CM|AB|692.3|Topical med dermatitis
C0157712|ICD9CM|PT|692.4|Contact dermatitis and other eczema due to other chemical products
C0157712|ICD9CM|AB|692.4|Chemical dermatitis NEC
C0157713|ICD9CM|PT|692.5|Contact dermatitis and other eczema due to food in contact with skin
C0157713|ICD9CM|AB|692.5|Topical food dermatitis
C0157714|ICD9CM|PT|692.6|Contact dermatitis and other eczema due to plants [except food]
C0157714|ICD9CM|AB|692.6|Dermatitis due to plant
C0157715|ICD9CM|HT|692.7|Contact dermatitis and other eczema due to solar radiation
C0157718|ICD9CM|HT|693|Dermatitis due to substances taken internally
C0157718|ICD9CM|PT|693.9|Dermatitis due to unspecified substance taken internally
C0157718|ICD9CM|AB|693.9|Dermat d/t int agent NOS
C0157719|ICD9CM|PT|693.8|Dermatitis due to other specified substances taken internally
C0157719|ICD9CM|AB|693.8|Dermat d/t int agent NEC
C0157721|ICD9CM|PT|694.61|Benign mucous membrane pemphigoid with ocular involvement
C0157721|ICD9CM|AB|694.61|Ocular pemphigus
C0157723|ICD9CM|HT|696|Psoriasis and similar disorders
C0157724|ICD9CM|HT|698|Pruritus and related conditions
C0157725|ICD9CM|PT|698.8|Other specified pruritic conditions
C0157725|ICD9CM|AB|698.8|Pruritic conditions NEC
C0157726|ICD9CM|AB|700|Corns and callosities
C0157726|ICD9CM|PT|700|Corns and callosities
C0157727|ICD9CM|HT|701|Other hypertrophic and atrophic conditions of skin
C0157729|ICD9CM|PT|701.5|Other abnormal granulation tissue
C0157729|ICD9CM|AB|701.5|Abnormal granulation NEC
C0157730|ICD9CM|PT|702.8|Other specified dermatoses
C0157730|ICD9CM|AB|702.8|Other specf dermatoses
C0157731|ICD9CM|PT|703.8|Other specified diseases of nail
C0157731|ICD9CM|AB|703.8|Diseases of nail NEC
C0157733|ICD9CM|PT|704.2|Abnormalities of the hair
C0157733|ICD9CM|AB|704.2|Abnormalities of hair
C0157734|ICD9CM|AB|704.3|Variations in hair color
C0157734|ICD9CM|PT|704.3|Variations in hair color
C0157735|ICD9CM|HT|705.8|Other specified disorders of sweat glands
C0157735|ICD9CM|PT|705.89|Other specified disorders of sweat glands
C0157735|ICD9CM|AB|705.89|Sweat gland disorder NEC
C0157736|ICD9CM|PT|706.8|Other specified diseases of sebaceous glands
C0157736|ICD9CM|AB|706.8|Sebaceous gland dis NEC
C0157738|ICD9CM|HT|707|Chronic ulcer of skin
C0157740|ICD9CM|PT|707.8|Chronic ulcer of other specified sites
C0157740|ICD9CM|AB|707.8|Chronic skin ulcer NEC
C0157741|ICD9CM|AB|708.1|Idiopathic urticaria
C0157741|ICD9CM|PT|708.1|Idiopathic urticaria
C0157742|ICD9CM|PT|708.2|Urticaria due to cold and heat
C0157742|ICD9CM|AB|708.2|Urticaria from cold/heat
C0157743|ICD9CM|AB|708.4|Vibratory urticaria
C0157743|ICD9CM|PT|708.4|Vibratory urticaria
C0157746|ICD9CM|PT|709.4|Foreign body granuloma of skin and subcutaneous tissue
C0157746|ICD9CM|AB|709.4|Foreign body granul-skin
C0157748|ICD9CM|PT|710.8|Other specified diffuse diseases of connective tissue
C0157748|ICD9CM|AB|710.8|Diff connect tis dis NEC
C0157749|ICD9CM|HT|711|Arthropathy associated with infections
C0157756|ICD9CM|PT|711.07|Pyogenic arthritis, ankle and foot
C0157756|ICD9CM|AB|711.07|Pyogen arthritis-ankle
C0157760|ICD9CM|PT|711.10|Arthropathy associated with Reiter's disease and nonspecific urethritis, site unspecified
C0157760|ICD9CM|HT|711.1|Arthropathy associated with Reiter's disease and nonspecific urethritis
C0157760|ICD9CM|AB|711.10|Reiter arthritis-unspec
C0157761|ICD9CM|PT|711.11|Arthropathy associated with Reiter's disease and nonspecific urethritis, shoulder region
C0157761|ICD9CM|AB|711.11|Reiter arthritis-shlder
C0157762|ICD9CM|PT|711.12|Arthropathy associated with Reiter's disease and nonspecific urethritis, upper arm
C0157762|ICD9CM|AB|711.12|Reiter arthritis-up/arm
C0157763|ICD9CM|PT|711.13|Arthropathy associated with Reiter's disease and nonspecific urethritis, forearm
C0157763|ICD9CM|AB|711.13|Reiter arthritis-forearm
C0157764|ICD9CM|PT|711.14|Arthropathy associated with Reiter's disease and nonspecific urethritis, hand
C0157764|ICD9CM|AB|711.14|Reiter arthritis-hand
C0157765|ICD9CM|PT|711.15|Arthropathy associated with Reiter's disease and nonspecific urethritis, pelvic region and thigh
C0157765|ICD9CM|AB|711.15|Reiter arthritis-pelvis
C0157766|ICD9CM|PT|711.16|Arthropathy associated with Reiter's disease and nonspecific urethritis, lower leg
C0157766|ICD9CM|AB|711.16|Reiter arthritis-l/leg
C0157767|ICD9CM|PT|711.17|Arthropathy associated with Reiter's disease and nonspecific urethritis, ankle and foot
C0157767|ICD9CM|AB|711.17|Reiter arthritis-ankle
C0157768|ICD9CM|PT|711.18|Arthropathy associated with Reiter's disease and nonspecific urethritis, other specified sites
C0157768|ICD9CM|AB|711.18|Reiter arthritis NEC
C0157769|ICD9CM|PT|711.19|Arthropathy associated with Reiter's disease and nonspecific urethritis, multiple sites
C0157769|ICD9CM|AB|711.19|Reiter arthritis-mult
C0157770|ICD9CM|HT|711.2|Arthropathy in Behcet's syndrome
C0157770|ICD9CM|PT|711.20|Arthropathy in Behcet's syndrome, site unspecified
C0157770|ICD9CM|AB|711.20|Behcet arthritis-unspec
C0157787|ICD9CM|PT|711.38|Postdysenteric arthropathy, other specified sites
C0157787|ICD9CM|AB|711.38|Dysenter arthrit NEC
C0157790|ICD9CM|PT|711.40|Arthropathy associated with other bacterial diseases, site unspecified
C0157790|ICD9CM|HT|711.4|Arthropathy associated with other bacterial diseases
C0157790|ICD9CM|AB|711.40|Bact arthritis-unspec
C0157801|ICD9CM|PT|711.50|Arthropathy associated with other viral diseases, site unspecified
C0157801|ICD9CM|HT|711.5|Arthropathy associated with other viral diseases
C0157801|ICD9CM|AB|711.50|Viral arthritis-unspec
C0157805|ICD9CM|PT|711.54|Arthropathy associated with other viral diseases, hand
C0157805|ICD9CM|AB|711.54|Viral arthritis-hand
C0157821|ICD9CM|PT|711.69|Arthropathy associated with mycoses, involving multiple sites
C0157821|ICD9CM|AB|711.69|Mycotic arthritis-mult
C0157822|ICD9CM|HT|711.7|Arthropathy associated with helminthiasis
C0157824|ICD9CM|PT|711.71|Arthropathy associated with helminthiasis, shoulder region
C0157824|ICD9CM|AB|711.71|Helminth arthrit-shlder
C0157833|ICD9CM|PT|711.80|Arthropathy associated with other infectious and parasitic diseases, site unspecified
C0157833|ICD9CM|HT|711.8|Arthropathy associated with other infectious and parasitic diseases
C0157833|ICD9CM|AB|711.80|Inf arthritis NEC-unspec
C0157834|ICD9CM|PT|711.81|Arthropathy associated with other infectious and parasitic diseases, shoulder region
C0157834|ICD9CM|AB|711.81|Inf arthritis NEC-shlder
C0157835|ICD9CM|PT|711.82|Arthropathy associated with other infectious and parasitic diseases, upper arm
C0157835|ICD9CM|AB|711.82|Inf arthritis NEC-up/arm
C0157836|ICD9CM|PT|711.83|Arthropathy associated with other infectious and parasitic diseases, forearm
C0157836|ICD9CM|AB|711.83|Inf arthrit NEC-forearm
C0157837|ICD9CM|PT|711.84|Arthropathy associated with other infectious and parasitic diseases, hand
C0157837|ICD9CM|AB|711.84|Inf arthritis NEC-hand
C0157838|ICD9CM|PT|711.85|Arthropathy associated with other infectious and parasitic diseases, pelvic region and thigh
C0157838|ICD9CM|AB|711.85|Inf arthritis NEC-pelvis
C0157839|ICD9CM|PT|711.86|Arthropathy associated with other infectious and parasitic diseases, lower leg
C0157839|ICD9CM|AB|711.86|Inf arthritis NEC-l/leg
C0157840|ICD9CM|PT|711.87|Arthropathy associated with other infectious and parasitic diseases, ankle and foot
C0157840|ICD9CM|AB|711.87|Inf arthritis NEC-ankle
C0157841|ICD9CM|PT|711.88|Arthropathy associated with other infectious and parasitic diseases, other specified sites
C0157841|ICD9CM|AB|711.88|Inf arthrit NEC-oth site
C0157842|ICD9CM|PT|711.89|Arthropathy associated with other infectious and parasitic diseases, multiple sites
C0157842|ICD9CM|AB|711.89|Inf arthritis NEC-mult
C0157843|ICD9CM|PT|711.91|Unspecified infective arthritis, shoulder region
C0157843|ICD9CM|AB|711.91|Inf arthritis NOS-shlder
C0157844|ICD9CM|PT|711.92|Unspecified infective arthritis, upper arm
C0157844|ICD9CM|AB|711.92|Inf arthritis NOS-up/arm
C0157845|ICD9CM|PT|711.93|Unspecified infective arthritis, forearm
C0157845|ICD9CM|AB|711.93|Inf arthrit NOS-forearm
C0157846|ICD9CM|PT|711.94|Unspecified infective arthritis, hand
C0157846|ICD9CM|AB|711.94|Inf arthrit NOS-hand
C0157847|ICD9CM|PT|711.95|Unspecified infective arthritis, pelvic region and thigh
C0157847|ICD9CM|AB|711.95|Inf arthrit NOS-pelvis
C0157848|ICD9CM|PT|711.96|Unspecified infective arthritis, lower leg
C0157848|ICD9CM|AB|711.96|Inf arthrit NOS-l/leg
C0157849|ICD9CM|PT|711.97|Unspecified infective arthritis, ankle and foot
C0157849|ICD9CM|AB|711.97|Inf arthrit NOS-ankle
C0157850|ICD9CM|PT|711.98|Unspecified infective arthritis, other specified sites
C0157850|ICD9CM|AB|711.98|Inf arthrit NOS-oth site
C0157851|ICD9CM|PT|711.99|Unspecified infective arthritis, multiple sites
C0157851|ICD9CM|AB|711.99|Inf arthritis NOS-mult
C0157852|ICD9CM|HT|712.1|Chondrocalcinosis due to dicalcium phosphate crystals
C0157874|ICD9CM|PT|712.30|Chondrocalcinosis, unspecified, site unspecified
C0157874|ICD9CM|AB|712.30|Chondrocalcin NOS-unspec
C0157884|ICD9CM|HT|712.8|Other specified crystal arthropathies
C0157884|ICD9CM|PT|712.80|Other specified crystal arthropathies, site unspecified
C0157884|ICD9CM|AB|712.80|Cryst arthrop NEC-unspec
C0157892|ICD9CM|PT|712.88|Other specified crystal arthropathies, other specified sites
C0157892|ICD9CM|AB|712.88|Cry arthrop NEC-oth site
C0157904|ICD9CM|HT|713|Arthropathy associated with other disorders classified elsewhere
C0157911|ICD9CM|PT|713.7|Other general diseases with articular involvement
C0157911|ICD9CM|AB|713.7|Arthrop w system dis NEC
C0157913|ICD9CM|HT|714|Rheumatoid arthritis and other inflammatory polyarthropathies
C0157914|ICD9CM|PT|714.2|Other rheumatoid arthritis with visceral or systemic involvement
C0157914|ICD9CM|AB|714.2|Syst rheum arthritis NEC
C0157916|ICD9CM|PT|714.31|Polyarticular juvenile rheumatoid arthritis, acute
C0157916|ICD9CM|AB|714.31|Polyart juv rheum arthr
C0157917|ICD9CM|PT|714.32|Pauciarticular juvenile rheumatoid arthritis
C0157917|ICD9CM|AB|714.32|Pauciart juv rheum arthr
C0157918|ICD9CM|PT|714.33|Monoarticular juvenile rheumatoid arthritis
C0157918|ICD9CM|AB|714.33|Monoart juv rheum arthr
C0157919|ICD9CM|HT|714.8|Other specified inflammatory polyarthropathies
C0157919|ICD9CM|PT|714.89|Other specified inflammatory polyarthropathies
C0157919|ICD9CM|AB|714.89|Inflamm polyarthrop NEC
C0157923|ICD9CM|PT|715.00|Osteoarthrosis, generalized, site unspecified
C0157923|ICD9CM|AB|715.00|General osteoarthrosis
C0157924|ICD9CM|PT|715.04|Osteoarthrosis, generalized, hand
C0157924|ICD9CM|AB|715.04|Gen osteoarthros-hand
C0157926|ICD9CM|HT|715.1|Osteoarthrosis, localized, primary
C0157926|ICD9CM|PT|715.10|Osteoarthrosis, localized, primary, site unspecified
C0157926|ICD9CM|AB|715.10|Loc prim osteoart-unspec
C0157937|ICD9CM|PT|715.20|Osteoarthrosis, localized, secondary, site unspecified
C0157937|ICD9CM|AB|715.20|Loc 2nd osteoarth-unspec
C0157938|ICD9CM|PT|715.21|Osteoarthrosis, localized, secondary, shoulder region
C0157938|ICD9CM|AB|715.21|Loc 2nd osteoarth-shlder
C0157939|ICD9CM|PT|715.22|Osteoarthrosis, localized, secondary, upper arm
C0157939|ICD9CM|AB|715.22|Loc 2nd osteoarth-up/arm
C0157940|ICD9CM|PT|715.23|Osteoarthrosis, localized, secondary, forearm
C0157940|ICD9CM|AB|715.23|Loc 2nd osteoart-forearm
C0157941|ICD9CM|PT|715.24|Osteoarthrosis, localized, secondary, hand
C0157941|ICD9CM|AB|715.24|Loc 2nd osteoarthro-hand
C0157942|ICD9CM|PT|715.25|Osteoarthrosis, localized, secondary, pelvic region and thigh
C0157942|ICD9CM|AB|715.25|Loc 2nd osteoarth-pelvis
C0157943|ICD9CM|PT|715.26|Osteoarthrosis, localized, secondary, lower leg
C0157943|ICD9CM|AB|715.26|Loc 2nd osteoarthr-l/leg
C0157944|ICD9CM|PT|715.27|Osteoarthrosis, localized, secondary, ankle and foot
C0157944|ICD9CM|AB|715.27|Loc 2nd osteoarthr-ankle
C0157945|ICD9CM|PT|715.28|Osteoarthrosis, localized, secondary, other specified sites
C0157945|ICD9CM|AB|715.28|Loc 2nd osteoarthros NEC
C0157946|ICD9CM|HT|715.3|Osteoarthrosis, localized, not specified whether primary or secondary
C0157947|ICD9CM|PT|715.30|Osteoarthrosis, localized, not specified whether primary or secondary, site unspecified
C0157947|ICD9CM|AB|715.30|Loc osteoarth NOS-unspec
C0157948|ICD9CM|PT|715.31|Osteoarthrosis, localized, not specified whether primary or secondary, shoulder region
C0157948|ICD9CM|AB|715.31|Loc osteoarth NOS-shlder
C0157949|ICD9CM|PT|715.32|Osteoarthrosis, localized, not specified whether primary or secondary, upper arm
C0157949|ICD9CM|AB|715.32|Loc osteoarth NOS-up/arm
C0157950|ICD9CM|PT|715.33|Osteoarthrosis, localized, not specified whether primary or secondary, forearm
C0157950|ICD9CM|AB|715.33|Loc osteoart NOS-forearm
C0157951|ICD9CM|PT|715.34|Osteoarthrosis, localized, not specified whether primary or secondary, hand
C0157951|ICD9CM|AB|715.34|Loc osteoarth NOS-hand
C0157952|ICD9CM|PT|715.35|Osteoarthrosis, localized, not specified whether primary or secondary, pelvic region and thigh
C0157952|ICD9CM|AB|715.35|Loc osteoarth NOS-pelvis
C0157953|ICD9CM|PT|715.36|Osteoarthrosis, localized, not specified whether primary or secondary, lower leg
C0157953|ICD9CM|AB|715.36|Loc osteoarth NOS-l/leg
C0157954|ICD9CM|PT|715.37|Osteoarthrosis, localized, not specified whether primary or secondary, ankle and foot
C0157954|ICD9CM|AB|715.37|Loc osteoarth NOS-ankle
C0157955|ICD9CM|PT|715.38|Osteoarthrosis, localized, not specified whether primary or secondary, other specified sites
C0157955|ICD9CM|AB|715.38|Loc osteoar NOS-site NEC
C0157957|ICD9CM|PT|715.80|Osteoarthrosis involving, or with mention of more than one site, but not specified as generalized, site unspecified
C0157957|ICD9CM|AB|715.80|Osteoarthrosis-mult site
C0157958|ICD9CM|PT|715.89|Osteoarthrosis involving, or with mention of more than one site, but not specified as generalized, multiple sites
C0157958|ICD9CM|AB|715.89|Osteoarthrosis-mult site
C0157959|ICD9CM|PT|715.90|Osteoarthrosis, unspecified whether generalized or localized, site unspecified
C0157959|ICD9CM|AB|715.90|Osteoarthros NOS-unspec
C0157960|ICD9CM|PT|715.91|Osteoarthrosis, unspecified whether generalized or localized, shoulder region
C0157960|ICD9CM|AB|715.91|Osteoarthros NOS-shlder
C0157961|ICD9CM|PT|715.92|Osteoarthrosis, unspecified whether generalized or localized, upper arm
C0157961|ICD9CM|AB|715.92|Osteoarthros NOS-up/arm
C0157962|ICD9CM|PT|715.93|Osteoarthrosis, unspecified whether generalized or localized, forearm
C0157962|ICD9CM|AB|715.93|Osteoarthros NOS-forearm
C0157963|ICD9CM|PT|715.94|Osteoarthrosis, unspecified whether generalized or localized, hand
C0157963|ICD9CM|AB|715.94|Osteoarthros NOS-hand
C0157964|ICD9CM|PT|715.95|Osteoarthrosis, unspecified whether generalized or localized, pelvic region and thigh
C0157964|ICD9CM|AB|715.95|Osteoarthros NOS-pelvis
C0157965|ICD9CM|PT|715.96|Osteoarthrosis, unspecified whether generalized or localized, lower leg
C0157965|ICD9CM|AB|715.96|Osteoarthros NOS-l/leg
C0157966|ICD9CM|PT|715.97|Osteoarthrosis, unspecified whether generalized or localized, ankle and foot
C0157966|ICD9CM|AB|715.97|Osteoarthros NOS-ankle
C0157967|ICD9CM|PT|715.98|Osteoarthrosis, unspecified whether generalized or localized, other specified sites
C0157967|ICD9CM|AB|715.98|Osteoarthro NOS-oth site
C0157969|ICD9CM|PT|716.01|Kaschin-Beck disease, shoulder region
C0157969|ICD9CM|AB|716.01|Kaschin-beck dis-shlder
C0157970|ICD9CM|PT|716.02|Kaschin-Beck disease, upper arm
C0157970|ICD9CM|AB|716.02|Kaschin-beck dis-up/arm
C0157971|ICD9CM|AB|716.03|Kaschin-beck dis-forearm
C0157971|ICD9CM|PT|716.03|Kaschin-Beck disease, forearm
C0157972|ICD9CM|AB|716.04|Kaschin-beck dis-hand
C0157972|ICD9CM|PT|716.04|Kaschin-Beck disease, hand
C0157974|ICD9CM|PT|716.06|Kaschin-Beck disease, lower leg
C0157974|ICD9CM|AB|716.06|Kaschin-beck dis-l/leg
C0157977|ICD9CM|PT|716.09|Kaschin-Beck disease, multiple sites
C0157977|ICD9CM|AB|716.09|Kaschin-beck dis-mult
C0157987|ICD9CM|HT|716.2|Allergic arthritis
C0157987|ICD9CM|PT|716.20|Allergic arthritis, site unspecified
C0157987|ICD9CM|AB|716.20|Allerg arthritis-unspec
C0157997|ICD9CM|HT|716.3|Climacteric arthritis
C0157997|ICD9CM|PT|716.30|Climacteric arthritis, site unspecified
C0157997|ICD9CM|AB|716.30|Climact arthritis-unspec
C0158004|ICD9CM|PT|716.37|Climacteric arthritis, ankle and foot
C0158004|ICD9CM|AB|716.37|Climact arthritis-ankle
C0158007|ICD9CM|PT|716.41|Transient arthropathy, shoulder region
C0158007|ICD9CM|AB|716.41|Trans arthropathy-shlder
C0158017|ICD9CM|PT|716.51|Unspecified polyarthropathy or polyarthritis, shoulder region
C0158017|ICD9CM|AB|716.51|Polyarthritis NOS-shlder
C0158018|ICD9CM|PT|716.52|Unspecified polyarthropathy or polyarthritis, upper arm
C0158018|ICD9CM|AB|716.52|Polyarthritis NOS-up/arm
C0158019|ICD9CM|PT|716.53|Unspecified polyarthropathy or polyarthritis, forearm
C0158019|ICD9CM|AB|716.53|Polyarthrit NOS-forearm
C0158020|ICD9CM|PT|716.54|Unspecified polyarthropathy or polyarthritis, hand
C0158020|ICD9CM|AB|716.54|Polyarthritis NOS-hand
C0158021|ICD9CM|PT|716.55|Unspecified polyarthropathy or polyarthritis, pelvic region and thigh
C0158021|ICD9CM|AB|716.55|Polyarthritis NOS-pelvis
C0158022|ICD9CM|PT|716.56|Unspecified polyarthropathy or polyarthritis, lower leg
C0158022|ICD9CM|AB|716.56|Polyarthritis NOS-l/leg
C0158023|ICD9CM|PT|716.57|Unspecified polyarthropathy or polyarthritis, ankle and foot
C0158023|ICD9CM|AB|716.57|Polyarthritis NOS-ankle
C0158024|ICD9CM|PT|716.58|Unspecified polyarthropathy or polyarthritis, other specified sites
C0158024|ICD9CM|AB|716.58|Polyarthrit NOS-oth site
C0158026|ICD9CM|HT|716.6|Unspecified monoarthritis
C0158026|ICD9CM|PT|716.60|Unspecified monoarthritis, site unspecified
C0158026|ICD9CM|AB|716.60|Monoarthritis NOS-unspec
C0158044|ICD9CM|PT|716.91|Arthropathy, unspecified, shoulder region
C0158044|ICD9CM|AB|716.91|Arthropathy NOS-shlder
C0158045|ICD9CM|PT|716.92|Arthropathy, unspecified, upper arm
C0158045|ICD9CM|AB|716.92|Arthropathy NOS-up/arm
C0158048|ICD9CM|PT|716.95|Arthropathy, unspecified, pelvic region and thigh
C0158048|ICD9CM|AB|716.95|Arthropathy NOS-pelvis
C0158049|ICD9CM|PT|716.96|Arthropathy, unspecified, lower leg
C0158049|ICD9CM|AB|716.96|Arthropathy NOS-l/leg
C0158050|ICD9CM|PT|716.97|Arthropathy, unspecified, ankle and foot
C0158050|ICD9CM|AB|716.97|Arthropathy NOS-ankle
C0158051|ICD9CM|PT|716.98|Arthropathy, unspecified, other specified sites
C0158051|ICD9CM|AB|716.98|Arthropathy NOS-oth site
C0158052|ICD9CM|PT|716.99|Arthropathy, unspecified, multiple sites
C0158052|ICD9CM|AB|716.99|Arthropathy NOS-mult
C0158053|ICD9CM|HT|717|Internal derangement of knee
C0158053|ICD9CM|PT|717.9|Unspecified internal derangement of knee
C0158053|ICD9CM|AB|717.9|Int derangement knee NOS
C0158054|ICD9CM|PT|717.0|Old bucket handle tear of medial meniscus
C0158054|ICD9CM|AB|717.0|Old bucket tear med men
C0158055|ICD9CM|PT|717.1|Derangement of anterior horn of medial meniscus
C0158055|ICD9CM|AB|717.1|Derang ant med meniscus
C0158056|ICD9CM|PT|717.2|Derangement of posterior horn of medial meniscus
C0158056|ICD9CM|AB|717.2|Derang post med meniscus
C0158057|ICD9CM|PT|717.3|Other and unspecified derangement of medial meniscus
C0158057|ICD9CM|AB|717.3|Derang med meniscus NEC
C0158058|ICD9CM|HT|717.4|Derangement of lateral meniscus
C0158058|ICD9CM|PT|717.40|Derangement of lateral meniscus, unspecified
C0158058|ICD9CM|AB|717.40|Derang lat meniscus NOS
C0158060|ICD9CM|PT|717.42|Derangement of anterior horn of lateral meniscus
C0158060|ICD9CM|AB|717.42|Derange ant lat meniscus
C0158061|ICD9CM|PT|717.43|Derangement of posterior horn of lateral meniscus
C0158061|ICD9CM|AB|717.43|Derang post lat meniscus
C0158062|ICD9CM|PT|717.49|Other derangement of lateral meniscus
C0158062|ICD9CM|AB|717.49|Derang lat meniscus NEC
C0158065|ICD9CM|HT|717.8|Other internal derangement of knee
C0158065|ICD9CM|PT|717.89|Other internal derangement of knee
C0158065|ICD9CM|AB|717.89|Int derangement knee NEC
C0158066|ICD9CM|PT|717.81|Old disruption of lateral collateral ligament
C0158066|ICD9CM|AB|717.81|Old disrupt lat collat
C0158067|ICD9CM|PT|717.82|Old disruption of medial collateral ligament
C0158067|ICD9CM|AB|717.82|Old disrupt med collat
C0158068|ICD9CM|PT|717.83|Old disruption of anterior cruciate ligament
C0158068|ICD9CM|AB|717.83|Old disrupt ant cruciate
C0158069|ICD9CM|PT|717.84|Old disruption of posterior cruciate ligament
C0158069|ICD9CM|AB|717.84|Old disrupt post cruciat
C0158070|ICD9CM|PT|717.85|Old disruption of other ligaments of knee
C0158070|ICD9CM|AB|717.85|Old disrupt knee lig NEC
C0158072|ICD9CM|HT|718|Other derangement of joint
C0158073|ICD9CM|HT|718.0|Articular cartilage disorder
C0158073|ICD9CM|PT|718.00|Articular cartilage disorder, site unspecified
C0158073|ICD9CM|AB|718.00|Artic cartil dis-unspec
C0158077|ICD9CM|PT|718.04|Articular cartilage disorder, hand
C0158077|ICD9CM|AB|718.04|Artic cartil dis-hand
C0158082|ICD9CM|PT|718.11|Loose body in joint, shoulder region
C0158082|ICD9CM|AB|718.11|Loose body-shlder
C0158083|ICD9CM|PT|718.12|Loose body in joint, upper arm
C0158083|ICD9CM|AB|718.12|Loose body-up/arm
C0158084|ICD9CM|PT|718.13|Loose body in joint, forearm
C0158084|ICD9CM|AB|718.13|Loose body-forearm
C0158085|ICD9CM|PT|718.14|Loose body in joint, hand
C0158085|ICD9CM|AB|718.14|Loose body-hand
C0158086|ICD9CM|PT|718.15|Loose body in joint, pelvic region and thigh
C0158086|ICD9CM|AB|718.15|Loose body-pelvis
C0158087|ICD9CM|PT|718.17|Loose body in joint, ankle and foot
C0158087|ICD9CM|AB|718.17|Loose body-ankle
C0158088|ICD9CM|PT|718.19|Loose body in joint, multiple sites
C0158088|ICD9CM|AB|718.19|Loose body-mult joints
C0158090|ICD9CM|HT|718.2|Pathological dislocation
C0158090|ICD9CM|PT|718.20|Pathological dislocation of joint, site unspecified
C0158090|ICD9CM|AB|718.20|Pathol dislocat-unspec
C0158091|ICD9CM|PT|718.21|Pathological dislocation of joint, shoulder region
C0158091|ICD9CM|AB|718.21|Pathol dislocat-shlder
C0158094|ICD9CM|PT|718.24|Pathological dislocation of joint, hand
C0158094|ICD9CM|AB|718.24|Pathol dislocat-hand
C0158095|ICD9CM|PT|718.25|Pathological dislocation of joint, pelvic region and thigh
C0158095|ICD9CM|AB|718.25|Pathol dislocat-pelvis
C0158098|ICD9CM|PT|718.28|Pathological dislocation of joint, other specified sites
C0158098|ICD9CM|AB|718.28|Pathol dislocat-jt NEC
C0158100|ICD9CM|HT|718.3|Recurrent dislocation of joint
C0158100|ICD9CM|PT|718.30|Recurrent dislocation of joint, site unspecified
C0158100|ICD9CM|AB|718.30|Recur dislocat-unspec
C0158105|ICD9CM|PT|718.35|Recurrent dislocation of joint, pelvic region and thigh
C0158105|ICD9CM|AB|718.35|Recur dislocat-pelvis
C0158108|ICD9CM|PT|718.38|Recurrent dislocation of joint, other specified sites
C0158108|ICD9CM|AB|718.38|Recur dislocat-jt NEC
C0158110|ICD9CM|PT|718.41|Contracture of joint, shoulder region
C0158110|ICD9CM|AB|718.41|Jt contracture-shlder
C0158111|ICD9CM|PT|718.42|Contracture of joint, upper arm
C0158111|ICD9CM|AB|718.42|Jt contracture-up/arm
C0158112|ICD9CM|PT|718.43|Contracture of joint, forearm
C0158112|ICD9CM|AB|718.43|Jt contracture-forearm
C0158113|ICD9CM|PT|718.44|Contracture of joint, hand
C0158113|ICD9CM|AB|718.44|Jt contracture-hand
C0158115|ICD9CM|PT|718.46|Contracture of joint, lower leg
C0158115|ICD9CM|AB|718.46|Jt contracture-l/leg
C0158117|ICD9CM|PT|718.48|Contracture of joint, other specified sites
C0158117|ICD9CM|AB|718.48|Jt contracture-jt NEC
C0158118|ICD9CM|PT|718.49|Contracture of joint, multiple sites
C0158118|ICD9CM|AB|718.49|Jt contracture-mult jts
C0158119|ICD9CM|PT|718.51|Ankylosis of joint, shoulder region
C0158119|ICD9CM|AB|718.51|Ankylosis-shoulder
C0158120|ICD9CM|PT|718.52|Ankylosis of joint, upper arm
C0158120|ICD9CM|AB|718.52|Ankylosis-upper/arm
C0158121|ICD9CM|PT|718.53|Ankylosis of joint, forearm
C0158121|ICD9CM|AB|718.53|Ankylosis-forearm
C0158122|ICD9CM|PT|718.54|Ankylosis of joint, hand
C0158122|ICD9CM|AB|718.54|Ankylosis-hand
C0158123|ICD9CM|PT|718.55|Ankylosis of joint, pelvic region and thigh
C0158123|ICD9CM|AB|718.55|Ankylosis-pelvis
C0158124|ICD9CM|PT|718.56|Ankylosis of joint, lower leg
C0158124|ICD9CM|AB|718.56|Ankylosis-lower/leg
C0158126|ICD9CM|PT|718.58|Ankylosis of joint, other specified sites
C0158126|ICD9CM|AB|718.58|Ankylosis-joint NEC
C0158127|ICD9CM|PT|718.59|Ankylosis of joint, multiple sites
C0158127|ICD9CM|AB|718.59|Ankylosis-mult joints
C0158128|ICD9CM|HT|718.6|Unspecified intrapelvic protrusion of acetabulum
C0158129|ICD9CM|PT|718.65|Unspecified intrapelvic protrusion of acetabulum, pelvic region and thigh
C0158129|ICD9CM|AB|718.65|Protrusio acetabuli NOS
C0158140|ICD9CM|HT|718.9|Unspecified derangement of joint
C0158140|ICD9CM|PT|718.90|Unspecified derangement of joint, site unspecified
C0158140|ICD9CM|AB|718.90|Jt derangmnt NOS-unsp jt
C0158150|ICD9CM|PT|719.01|Effusion of joint, shoulder region
C0158150|ICD9CM|AB|719.01|Joint effusion-shlder
C0158151|ICD9CM|PT|719.02|Effusion of joint, upper arm
C0158151|ICD9CM|AB|719.02|Joint effusion-up/arm
C0158152|ICD9CM|AB|719.03|Joint effusion-forearm
C0158152|ICD9CM|PT|719.03|Effusion of joint, forearm
C0158153|ICD9CM|AB|719.04|Joint effusion-hand
C0158153|ICD9CM|PT|719.04|Effusion of joint, hand
C0158155|ICD9CM|PT|719.06|Effusion of joint, lower leg
C0158155|ICD9CM|AB|719.06|Joint effusion-l/leg
C0158156|ICD9CM|PT|719.07|Effusion of joint, ankle and foot
C0158156|ICD9CM|AB|719.07|Joint effusion-ankle
C0158157|ICD9CM|PT|719.08|Effusion of joint, other specified sites
C0158157|ICD9CM|AB|719.08|Joint effusion-jt NEC
C0158158|ICD9CM|PT|719.09|Effusion of joint, multiple sites
C0158158|ICD9CM|AB|719.09|Joint effusion-mult jts
C0158159|ICD9CM|PT|719.11|Hemarthrosis, shoulder region
C0158159|ICD9CM|AB|719.11|Hemarthrosis-shlder
C0158162|ICD9CM|PT|719.14|Hemarthrosis, hand
C0158162|ICD9CM|AB|719.14|Hemarthrosis-hand
C0158167|ICD9CM|PT|719.19|Hemarthrosis, multiple sites
C0158167|ICD9CM|AB|719.19|Hemarthrosis-mult jts
C0158168|ICD9CM|HT|719.2|Villonodular synovitis
C0158168|ICD9CM|PT|719.20|Villonodular synovitis, site unspecified
C0158168|ICD9CM|AB|719.20|Villonod synovit-unspec
C0158169|ICD9CM|PT|719.21|Villonodular synovitis, shoulder region
C0158169|ICD9CM|AB|719.21|Villonod synovit-shlder
C0158175|ICD9CM|PT|719.27|Villonodular synovitis, ankle and foot
C0158175|ICD9CM|AB|719.27|Villonod synovit-ankle
C0158178|ICD9CM|PT|719.31|Palindromic rheumatism, shoulder region
C0158178|ICD9CM|AB|719.31|Palindrom rheum-shlder
C0158181|ICD9CM|PT|719.34|Palindromic rheumatism, hand
C0158181|ICD9CM|AB|719.34|Palindrom rheum-hand
C0158186|ICD9CM|PT|719.39|Palindromic rheumatism, multiple sites
C0158186|ICD9CM|AB|719.39|Palindrom rheum-mult jts
C0158194|ICD9CM|PT|719.48|Pain in joint, other specified sites
C0158194|ICD9CM|AB|719.48|Joint pain-jt NEC
C0158195|ICD9CM|PT|719.50|Stiffness of joint, not elsewhere classified, site unspecified
C0158195|ICD9CM|AB|719.50|Jt stiffness NEC-unspec
C0158196|ICD9CM|PT|719.51|Stiffness of joint, not elsewhere classified, shoulder region
C0158196|ICD9CM|AB|719.51|Jt stiffness NEC-shlder
C0158197|ICD9CM|PT|719.52|Stiffness of joint, not elsewhere classified, upper arm
C0158197|ICD9CM|AB|719.52|Jt stiffness NEC-up/arm
C0158198|ICD9CM|PT|719.53|Stiffness of joint, not elsewhere classified, forearm
C0158198|ICD9CM|AB|719.53|Jt stiffnes NEC-forearm
C0158199|ICD9CM|PT|719.54|Stiffness of joint, not elsewhere classified, hand
C0158199|ICD9CM|AB|719.54|Jt stiffness NEC-hand
C0158200|ICD9CM|PT|719.55|Stiffness of joint, not elsewhere classified, pelvic region and thigh
C0158200|ICD9CM|AB|719.55|Jt stiffness NEC-pelvis
C0158201|ICD9CM|PT|719.56|Stiffness of joint, not elsewhere classified, lower leg
C0158201|ICD9CM|AB|719.56|Jt stiffness NEC-l/leg
C0158202|ICD9CM|PT|719.57|Stiffness of joint, not elsewhere classified, ankle and foot
C0158202|ICD9CM|AB|719.57|Jt stiffness NEC-ankle
C0158203|MTH|PN|NOCODE|Stiffness of joint, NEC, involving other specified sites in ICD9CM
C0158203|ICD9CM|PT|719.58|Stiffness of joint, not elsewhere classified, other specified sites
C0158203|ICD9CM|AB|719.58|Jt stiffness NEC-oth jt
C0158204|ICD9CM|PT|719.59|Stiffness of joint, not elsewhere classified, multiple sites
C0158204|ICD9CM|AB|719.59|Jt stiffness NEC-mult jt
C0158205|ICD9CM|HT|719.6|Other symptoms referable to joint
C0158206|ICD9CM|PT|719.61|Other symptoms referable to joint, shoulder region
C0158206|ICD9CM|AB|719.61|Joint symptom NEC-shlder
C0158207|ICD9CM|PT|719.62|Other symptoms referable to joint, upper arm
C0158207|ICD9CM|AB|719.62|Joint symptom NEC-up/arm
C0158208|ICD9CM|PT|719.63|Other symptoms referable to joint, forearm
C0158208|ICD9CM|AB|719.63|Joint sympt NEC-forearm
C0158209|ICD9CM|PT|719.64|Other symptoms referable to joint, hand
C0158209|ICD9CM|AB|719.64|Joint symptom NEC-hand
C0158210|ICD9CM|PT|719.65|Other symptoms referable to joint, pelvic region and thigh
C0158210|ICD9CM|AB|719.65|Joint symptom NEC-pelvis
C0158211|ICD9CM|PT|719.66|Other symptoms referable to joint, lower leg
C0158211|ICD9CM|AB|719.66|Joint symptom NEC-l/leg
C0158212|ICD9CM|PT|719.67|Other symptoms referable to joint, ankle and foot
C0158212|ICD9CM|AB|719.67|Joint symptom NEC-ankle
C0158213|ICD9CM|PT|719.68|Other symptoms referable to joint, other specified sites
C0158213|ICD9CM|AB|719.68|Joint symptom NEC-oth jt
C0158214|ICD9CM|PT|719.69|Other symptoms referable to joint, multiple sites
C0158214|ICD9CM|AB|719.69|Joint sympt NEC-mult jts
C0158222|ICD9CM|PT|719.81|Other specified disorders of joint, shoulder region
C0158222|ICD9CM|AB|719.81|Joint dis NEC-shlder
C0158223|ICD9CM|PT|719.82|Other specified disorders of joint, upper arm
C0158223|ICD9CM|AB|719.82|Joint dis NEC-up/arm
C0158224|ICD9CM|PT|719.83|Other specified disorders of joint, forearm
C0158224|ICD9CM|AB|719.83|Joint dis NEC-forearm
C0158225|ICD9CM|PT|719.84|Other specified disorders of joint, hand
C0158225|ICD9CM|AB|719.84|Joint dis NEC-hand
C0158226|ICD9CM|PT|719.85|Other specified disorders of joint, pelvic region and thigh
C0158226|ICD9CM|AB|719.85|Joint dis NEC-pelvis
C0158227|ICD9CM|PT|719.86|Other specified disorders of joint, lower leg
C0158227|ICD9CM|AB|719.86|Joint dis NEC-l/leg
C0158228|ICD9CM|PT|719.87|Other specified disorders of joint, ankle and foot
C0158228|ICD9CM|AB|719.87|Joint dis NEC-ankle
C0158229|ICD9CM|PT|719.88|Other specified disorders of joint, other specified sites
C0158229|ICD9CM|AB|719.88|Joint dis NEC-oth jt
C0158230|ICD9CM|PT|719.89|Other specified disorders of joint, multiple sites
C0158230|ICD9CM|AB|719.89|Joint dis NEC-mult jts
C0158231|ICD9CM|PT|719.91|Unspecified disorder of joint, shoulder region
C0158231|ICD9CM|AB|719.91|Joint dis NOS-shlder
C0158232|ICD9CM|PT|719.92|Unspecified disorder of joint, upper arm
C0158232|ICD9CM|AB|719.92|Joint dis NOS-up/arm
C0158233|ICD9CM|PT|719.93|Unspecified disorder of joint, forearm
C0158233|ICD9CM|AB|719.93|Joint dis NOS-forearm
C0158234|ICD9CM|PT|719.94|Unspecified disorder of joint, hand
C0158234|ICD9CM|AB|716.94|Arthropathy NOS-hand
C0158234|ICD9CM|PT|716.94|Arthropathy, unspecified, hand
C0158234|ICD9CM|AB|719.94|Joint dis NOS-hand
C0158235|ICD9CM|PT|719.95|Unspecified disorder of joint, pelvic region and thigh
C0158235|ICD9CM|AB|719.95|Joint dis NOS-pelvis
C0158236|ICD9CM|PT|719.96|Unspecified disorder of joint, lower leg
C0158236|ICD9CM|AB|719.96|Joint dis NOS-l/leg
C0158239|ICD9CM|PT|719.99|Unspecified disorder of joint, multiple sites
C0158239|ICD9CM|AB|719.99|Joint dis NOS-mult jts
C0158240|ICD9CM|HT|721|Spondylosis and allied disorders
C0158241|ICD9CM|PT|721.0|Cervical spondylosis without myelopathy
C0158241|ICD9CM|AB|721.0|Cervical spondylosis
C0158242|ICD9CM|PT|721.1|Cervical spondylosis with myelopathy
C0158242|ICD9CM|AB|721.1|Cerv spondyl w myelopath
C0158243|ICD9CM|PT|721.2|Thoracic spondylosis without myelopathy
C0158243|ICD9CM|AB|721.2|Thoracic spondylosis
C0158244|ICD9CM|PT|721.3|Lumbosacral spondylosis without myelopathy
C0158244|ICD9CM|AB|721.3|Lumbosacral spondylosis
C0158245|ICD9CM|HT|721.4|Thoracic or lumbar spondylosis with myelopathy
C0158246|ICD9CM|PT|721.41|Spondylosis with myelopathy, thoracic region
C0158246|ICD9CM|AB|721.41|Spond compr thor sp cord
C0158247|ICD9CM|PT|721.42|Spondylosis with myelopathy, lumbar region
C0158247|ICD9CM|AB|721.42|Spond compr lumb sp cord
C0158248|ICD9CM|AB|721.5|Kissing spine
C0158248|ICD9CM|PT|721.5|Kissing spine
C0158249|ICD9CM|PT|721.8|Other allied disorders of spine
C0158249|ICD9CM|AB|721.8|Spinal disorders NEC
C0158252|ICD9CM|HT|722|Intervertebral disc disorders
C0158253|ICD9CM|PT|722.0|Displacement of cervical intervertebral disc without myelopathy
C0158253|ICD9CM|AB|722.0|Cervical disc displacmnt
C0158254|ICD9CM|HT|722.1|Displacement of thoracic or lumbar intervertebral disc without myelopathy
C0158255|ICD9CM|PT|722.10|Displacement of lumbar intervertebral disc without myelopathy
C0158255|ICD9CM|AB|722.10|Lumbar disc displacement
C0158256|ICD9CM|PT|722.11|Displacement of thoracic intervertebral disc without myelopathy
C0158256|ICD9CM|AB|722.11|Thoracic disc displacmnt
C0158259|ICD9CM|PT|722.31|Schmorl's nodes, thoracic region
C0158259|ICD9CM|AB|722.31|Schmorls node-thoracic
C0158260|ICD9CM|PT|722.32|Schmorl's nodes, lumbar region
C0158260|ICD9CM|AB|722.32|Schmorls node-lumbar
C0158261|ICD9CM|PT|722.39|Schmorl's nodes, other region
C0158261|ICD9CM|AB|722.39|Schmorls node-region NEC
C0158262|ICD9CM|PT|722.4|Degeneration of cervical intervertebral disc
C0158262|ICD9CM|AB|722.4|Cervical disc degen
C0158263|ICD9CM|HT|722.5|Degeneration of thoracic or lumbar intervertebral disc
C0158264|ICD9CM|PT|722.51|Degeneration of thoracic or thoracolumbar intervertebral disc
C0158264|ICD9CM|AB|722.51|Thoracic disc degen
C0158265|ICD9CM|PT|722.52|Degeneration of lumbar or lumbosacral intervertebral disc
C0158265|ICD9CM|AB|722.52|Lumb/lumbosac disc degen
C0158266|ICD9CM|PT|722.6|Degeneration of intervertebral disc, site unspecified
C0158266|ICD9CM|AB|722.6|Disc degeneration NOS
C0158267|ICD9CM|HT|722.7|Intervertebral disc disorder with myelopathy
C0158268|ICD9CM|PT|722.71|Intervertebral disc disorder with myelopathy, cervical region
C0158268|ICD9CM|AB|722.71|Cerv disc dis w myelopat
C0158269|ICD9CM|PT|722.72|Intervertebral disc disorder with myelopathy, thoracic region
C0158269|ICD9CM|AB|722.72|Thor disc dis w myelopat
C0158270|ICD9CM|PT|722.73|Intervertebral disc disorder with myelopathy, lumbar region
C0158270|ICD9CM|AB|722.73|Lumb disc dis w myelopat
C0158272|ICD9CM|PT|722.81|Postlaminectomy syndrome, cervical region
C0158272|ICD9CM|AB|722.81|Postlaminect synd-cerv
C0158273|ICD9CM|PT|722.82|Postlaminectomy syndrome, thoracic region
C0158273|ICD9CM|AB|722.82|Postlaminect synd-thorac
C0158274|ICD9CM|PT|722.83|Postlaminectomy syndrome, lumbar region
C0158274|ICD9CM|AB|722.83|Postlaminect synd-lumbar
C0158275|ICD9CM|HT|722.9|Other and unspecified disc disorder
C0158276|ICD9CM|PT|722.91|Other and unspecified disc disorder, cervical region
C0158276|ICD9CM|AB|722.91|Disc dis NEC/NOS-cerv
C0158277|ICD9CM|PT|722.92|Other and unspecified disc disorder, thoracic region
C0158277|ICD9CM|AB|722.92|Disc dis NEC/NOS-thorac
C0158278|ICD9CM|PT|722.93|Other and unspecified disc disorder, lumbar region
C0158278|ICD9CM|AB|722.93|Disc dis NEC/NOS-lumbar
C0158279|ICD9CM|HT|723|Other disorders of cervical region
C0158280|ICD9CM|PT|723.0|Spinal stenosis in cervical region
C0158280|ICD9CM|AB|723.0|Cervical spinal stenosis
C0158281|ICD9CM|AB|723.3|Cervicobrachial syndrome
C0158281|ICD9CM|PT|723.3|Cervicobrachial syndrome (diffuse)
C0158284|MTH|PN|NOCODE|Cervical syndrome NEC in ICD9CM_2014
C0158284|ICD9CM|PT|723.8|Other syndromes affecting cervical region
C0158284|ICD9CM|AB|723.8|Cervical syndrome NEC
C0158285|ICD9CM|PT|723.9|Unspecified musculoskeletal disorders and symptoms referable to neck
C0158285|ICD9CM|AB|723.9|Neck disorder/sympt NOS
C0158287|ICD9CM|PT|724.01|Spinal stenosis, thoracic region
C0158287|ICD9CM|AB|724.01|Spinal stenosis-thoracic
C0158289|ICD9CM|PT|724.09|Spinal stenosis, other region
C0158289|ICD9CM|AB|724.09|Spinal stenosis-oth site
C0158291|ICD9CM|PT|724.4|Thoracic or lumbosacral neuritis or radiculitis, unspecified
C0158291|ICD9CM|AB|724.4|Lumbosacral neuritis NOS
C0158292|ICD9CM|AB|724.6|Disorders of sacrum
C0158292|ICD9CM|PT|724.6|Disorders of sacrum
C0158293|ICD9CM|HT|724.7|Disorders of coccyx
C0158293|ICD9CM|AB|724.70|Disorder of coccyx NOS
C0158293|ICD9CM|PT|724.70|Unspecified disorder of coccyx
C0158295|ICD9CM|AB|724.71|Hypermobility of coccyx
C0158295|ICD9CM|PT|724.71|Hypermobility of coccyx
C0158296|ICD9CM|PT|724.79|Other disorders of coccyx
C0158296|ICD9CM|AB|724.79|Disorder of coccyx NEC
C0158297|ICD9CM|PT|724.8|Other symptoms referable to back
C0158297|ICD9CM|AB|724.8|Other back symptoms
C0158298|ICD9CM|HT|724|Other and unspecified disorders of back
C0158298|ICD9CM|PT|724.9|Other unspecified back disorders
C0158298|ICD9CM|AB|724.9|Back disorder NOS
C0158301|ICD9CM|HT|726.1|Rotator cuff syndrome of shoulder and allied disorders
C0158302|ICD9CM|PT|726.10|Disorders of bursae and tendons in shoulder region, unspecified
C0158302|ICD9CM|AB|726.10|Rotator cuff synd NOS
C0158303|ICD9CM|PT|726.11|Calcifying tendinitis of shoulder
C0158303|ICD9CM|AB|726.11|Calcif tendinitis shlder
C0158304|ICD9CM|AB|726.12|Bicipital tenosynovitis
C0158304|ICD9CM|PT|726.12|Bicipital tenosynovitis
C0158305|ICD9CM|PT|726.19|Other specified disorders of bursae and tendons in shoulder region
C0158305|ICD9CM|AB|726.19|Rotator cuff dis NEC
C0158307|ICD9CM|HT|726.3|Enthesopathy of elbow region
C0158307|ICD9CM|AB|726.30|Elbow enthesopathy NOS
C0158307|ICD9CM|PT|726.30|Enthesopathy of elbow, unspecified
C0158309|ICD9CM|AB|726.31|Medial epicondylitis
C0158309|ICD9CM|PT|726.31|Medial epicondylitis
C0158310|ICD9CM|PT|726.39|Other enthesopathy of elbow region
C0158310|ICD9CM|AB|726.39|Elbow enthesopathy NEC
C0158311|ICD9CM|PT|726.4|Enthesopathy of wrist and carpus
C0158311|ICD9CM|AB|726.4|Enthesopathy of wrist
C0158312|ICD9CM|PT|726.5|Enthesopathy of hip region
C0158312|ICD9CM|AB|726.5|Enthesopathy of hip
C0158313|ICD9CM|HT|726.6|Enthesopathy of knee
C0158313|ICD9CM|AB|726.60|Enthesopathy of knee NOS
C0158313|ICD9CM|PT|726.60|Enthesopathy of knee, unspecified
C0158314|ICD9CM|PT|726.61|Pes anserinus tendinitis or bursitis
C0158314|ICD9CM|AB|726.61|Pes anserinus tendinitis
C0158315|ICD9CM|PT|726.62|Tibial collateral ligament bursitis
C0158315|ICD9CM|AB|726.62|Tibial coll lig bursitis
C0158316|ICD9CM|PT|726.63|Fibular collateral ligament bursitis
C0158316|ICD9CM|AB|726.63|Fibula coll lig bursitis
C0158317|ICD9CM|AB|726.64|Patellar tendinitis
C0158317|ICD9CM|PT|726.64|Patellar tendinitis
C0158318|ICD9CM|PT|726.69|Other enthesopathy of knee
C0158318|ICD9CM|AB|726.69|Enthesopathy of knee NEC
C0158319|ICD9CM|HT|726.7|Enthesopathy of ankle and tarsus
C0158319|ICD9CM|PT|726.70|Enthesopathy of ankle and tarsus, unspecified
C0158319|ICD9CM|AB|726.70|Ankle enthesopathy NOS
C0158321|ICD9CM|AB|726.72|Tibialis tendinitis
C0158321|ICD9CM|PT|726.72|Tibialis tendinitis
C0158322|ICD9CM|AB|726.73|Calcaneal spur
C0158322|ICD9CM|PT|726.73|Calcaneal spur
C0158323|ICD9CM|PT|726.79|Other enthesopathy of ankle and tarsus
C0158323|ICD9CM|AB|726.79|Ankle enthesopathy NEC
C0158324|ICD9CM|PT|726.8|Other peripheral enthesopathies
C0158324|ICD9CM|AB|726.8|Periph enthesopathy NEC
C0158326|ICD9CM|HT|727|Other disorders of synovium, tendon, and bursa
C0158326|ICD9CM|HT|727.8|Other disorders of synovium, tendon, and bursa
C0158326|ICD9CM|PT|727.89|Other disorders of synovium, tendon, and bursa
C0158326|ICD9CM|AB|727.89|Synov/tend/bursa dis NEC
C0158327|ICD9CM|PT|727.01|Synovitis and tenosynovitis in diseases classified elsewhere
C0158327|ICD9CM|AB|727.01|Synovitis in oth dis
C0158331|ICD9CM|PT|727.06|Tenosynovitis of foot and ankle
C0158331|ICD9CM|AB|727.06|Tenosynovitis foot/ankle
C0158332|ICD9CM|PT|727.2|Specific bursitides often of occupational origin
C0158332|ICD9CM|AB|727.2|Occupational bursitis
C0158334|ICD9CM|AB|727.41|Ganglion of joint
C0158334|ICD9CM|PT|727.41|Ganglion of joint
C0158335|ICD9CM|PT|727.42|Ganglion of tendon sheath
C0158335|ICD9CM|AB|727.42|Ganglion of tendon
C0158336|ICD9CM|PT|727.49|Other ganglion and cyst of synovium, tendon, and bursa
C0158336|ICD9CM|AB|727.49|Bursal cyst NEC
C0158337|ICD9CM|HT|727.5|Rupture of synovium
C0158337|ICD9CM|AB|727.50|Rupture of synovium NOS
C0158337|ICD9CM|PT|727.50|Rupture of synovium, unspecified
C0158338|ICD9CM|PT|727.59|Other rupture of synovium
C0158338|ICD9CM|AB|727.59|Rupture of synovium NEC
C0158339|ICD9CM|HT|727.6|Rupture of tendon, nontraumatic
C0158339|ICD9CM|PT|727.60|Nontraumatic rupture of unspecified tendon
C0158339|ICD9CM|AB|727.60|Nontraum tendon rupt NOS
C0158342|ICD9CM|PT|727.62|Nontraumatic rupture of tendons of biceps (long head)
C0158342|ICD9CM|AB|727.62|Biceps tendon rupture
C0158344|ICD9CM|PT|727.64|Nontraumatic rupture of flexor tendons of hand and wrist
C0158344|ICD9CM|AB|727.64|Rupt flexor tendon hand
C0158345|ICD9CM|PT|727.65|Nontraumatic rupture of quadriceps tendon
C0158345|ICD9CM|AB|727.65|Rupture quadricep tendon
C0158346|ICD9CM|AB|727.66|Rupture patellar tendon
C0158346|ICD9CM|PT|727.66|Nontraumatic rupture of patellar tendon
C0158347|ICD9CM|AB|727.67|Rupture achilles tendon
C0158347|ICD9CM|PT|727.67|Nontraumatic rupture of achilles tendon
C0158348|ICD9CM|PT|727.68|Nontraumatic rupture of other tendons of foot and ankle
C0158348|ICD9CM|AB|727.68|Rupture tendon foot NEC
C0158349|ICD9CM|PT|727.69|Nontraumatic rupture of other tendon
C0158349|ICD9CM|AB|727.69|Nontraum tendon rupt NEC
C0158350|ICD9CM|AB|727.81|Contracture of tendon
C0158350|ICD9CM|PT|727.81|Contracture of tendon (sheath)
C0158351|ICD9CM|PT|727.9|Unspecified disorder of synovium, tendon, and bursa
C0158351|ICD9CM|AB|727.9|Synov/tend/bursa dis NOS
C0158352|ICD9CM|HT|728|Disorders of muscle, ligament, and fascia
C0158352|ICD9CM|PT|728.9|Unspecified disorder of muscle, ligament, and fascia
C0158352|ICD9CM|AB|728.9|Muscle/ligament dis NOS
C0158353|ICD9CM|AB|728.0|Infective myositis
C0158353|ICD9CM|PT|728.0|Infective myositis
C0158355|ICD9CM|PT|728.10|Calcification and ossification, unspecified
C0158355|ICD9CM|AB|728.10|Muscular calcificat NOS
C0158357|ICD9CM|PT|728.13|Postoperative heterotopic calcification
C0158357|ICD9CM|AB|728.13|Postop heterotopic calc
C0158358|ICD9CM|PT|728.19|Other muscular calcification and ossification
C0158358|ICD9CM|AB|728.19|Muscular calcificat NEC
C0158359|ICD9CM|AB|728.4|Laxity of ligament
C0158359|ICD9CM|PT|728.4|Laxity of ligament
C0158360|ICD9CM|AB|728.71|Plantar fibromatosis
C0158360|ICD9CM|PT|728.71|Plantar fascial fibromatosis
C0158361|ICD9CM|HT|728.8|Other disorders of muscle, ligament, and fascia
C0158361|ICD9CM|PT|728.89|Other disorders of muscle, ligament, and fascia
C0158361|ICD9CM|AB|728.89|Muscle/ligament dis NEC
C0158362|ICD9CM|AB|728.81|Interstitial myositis
C0158362|ICD9CM|PT|728.81|Interstitial myositis
C0158363|ICD9CM|PT|728.83|Rupture of muscle, nontraumatic
C0158363|ICD9CM|AB|728.83|Nontraum muscle rupture
C0158364|ICD9CM|AB|728.84|Diastasis of muscle
C0158364|ICD9CM|PT|728.84|Diastasis of muscle
C0158366|ICD9CM|PT|729.31|Hypertrophy of fat pad, knee
C0158366|ICD9CM|AB|729.31|Hypertrophy of fat pad
C0158367|ICD9CM|PT|729.39|Panniculitis, other site
C0158367|ICD9CM|AB|729.39|Panniculitis, site NEC
C0158368|ICD9CM|PT|729.6|Residual foreign body in soft tissue
C0158368|ICD9CM|AB|729.6|Old FB in soft tissue
C0158369|ICD9CM|AB|729.81|Swelling of limb
C0158369|ICD9CM|PT|729.81|Swelling of limb
C0158370|ICD9CM|HT|729|Other disorders of soft tissues
C0158370|ICD9CM|PT|729.99|Other disorders of soft tissue
C0158370|ICD9CM|HT|729.9|Other and unspecified disorders of soft tissue
C0158370|ICD9CM|AB|729.99|Soft tissue disorder NEC
C0158371|ICD9CM|HT|730.0|Acute osteomyelitis
C0158371|ICD9CM|PT|730.00|Acute osteomyelitis, site unspecified
C0158371|ICD9CM|AB|730.00|Ac osteomyelitis-unspec
C0158372|ICD9CM|PT|730.01|Acute osteomyelitis, shoulder region
C0158372|ICD9CM|AB|730.01|Ac osteomyelitis-shlder
C0158373|ICD9CM|PT|730.02|Acute osteomyelitis, upper arm
C0158373|ICD9CM|AB|730.02|Ac osteomyelitis-up/arm
C0158374|ICD9CM|PT|730.03|Acute osteomyelitis, forearm
C0158374|ICD9CM|AB|730.03|Ac osteomyelitis-forearm
C0158375|ICD9CM|PT|730.04|Acute osteomyelitis, hand
C0158375|ICD9CM|AB|730.04|Ac osteomyelitis-hand
C0158377|ICD9CM|PT|730.06|Acute osteomyelitis, lower leg
C0158377|ICD9CM|AB|730.06|Ac osteomyelitis-l/leg
C0158380|ICD9CM|PT|730.09|Acute osteomyelitis, multiple sites
C0158380|ICD9CM|AB|730.09|Ac osteomyelitis-mult
C0158381|ICD9CM|PT|730.11|Chronic osteomyelitis, shoulder region
C0158381|ICD9CM|AB|730.11|Chr osteomyelit-shlder
C0158382|ICD9CM|PT|730.12|Chronic osteomyelitis, upper arm
C0158382|ICD9CM|AB|730.12|Chr osteomyelit-up/arm
C0158383|ICD9CM|PT|730.13|Chronic osteomyelitis, forearm
C0158383|ICD9CM|AB|730.13|Chr osteomyelit-forearm
C0158384|ICD9CM|PT|730.14|Chronic osteomyelitis, hand
C0158384|ICD9CM|AB|730.14|Chr osteomyelit-hand
C0158386|ICD9CM|PT|730.16|Chronic osteomyelitis, lower leg
C0158386|ICD9CM|AB|730.16|Chr osteomyelit-l/leg
C0158395|ICD9CM|PT|730.26|Unspecified osteomyelitis, lower leg
C0158395|ICD9CM|AB|730.26|Osteomyelitis NOS-l/leg
C0158396|ICD9CM|PT|730.27|Unspecified osteomyelitis, ankle and foot
C0158396|ICD9CM|AB|730.27|Osteomyelitis NOS-ankle
C0158401|ICD9CM|PT|730.32|Periostitis, without mention of osteomyelitis, upper arm
C0158401|ICD9CM|AB|730.32|Periostitis-up/arm
C0158402|ICD9CM|AB|730.33|Periostitis-forearm
C0158402|ICD9CM|PT|730.33|Periostitis, without mention of osteomyelitis, forearm
C0158403|ICD9CM|AB|730.34|Periostitis-hand
C0158403|ICD9CM|PT|730.34|Periostitis, without mention of osteomyelitis, hand
C0158405|ICD9CM|PT|730.36|Periostitis, without mention of osteomyelitis, lower leg
C0158405|ICD9CM|AB|730.36|Periostitis-l/leg
C0158406|ICD9CM|PT|730.37|Periostitis, without mention of osteomyelitis, ankle and foot
C0158406|ICD9CM|AB|730.37|Periostitis-ankle
C0158407|ICD9CM|PT|730.39|Periostitis, without mention of osteomyelitis, multiple sites
C0158407|ICD9CM|AB|730.39|Periostitis-mult
C0158408|ICD9CM|HT|730.7|Osteopathy resulting from poliomyelitis
C0158408|ICD9CM|PT|730.70|Osteopathy resulting from poliomyelitis, site unspecified
C0158408|ICD9CM|AB|730.70|Polio osteopathy-unspec
C0158420|ICD9CM|PT|730.81|Other infections involving bone in diseases classified elsewhere, shoulder region
C0158420|ICD9CM|AB|730.81|Bone infect NEC-shlder
C0158421|ICD9CM|PT|730.82|Other infections involving bone in diseases classified elsewhere, upper arm
C0158421|ICD9CM|AB|730.82|Bone infect NEC-up/arm
C0158422|ICD9CM|PT|730.83|Other infections involving bone in diseases classified elsewhere, forearm
C0158422|ICD9CM|AB|730.83|Bone infect NEC-forearm
C0158423|ICD9CM|PT|730.84|Other infections involving bone in diseases classified elsewhere, hand
C0158423|ICD9CM|AB|730.84|Bone infect NEC-hand
C0158424|ICD9CM|PT|730.85|Other infections involving bone in diseases classified elsewhere, pelvic region and thigh
C0158424|ICD9CM|AB|730.85|Bone infect NEC-pelvis
C0158425|ICD9CM|PT|730.86|Other infections involving bone in diseases classified elsewhere, lower leg
C0158425|ICD9CM|AB|730.86|Bone infect NEC-l/leg
C0158426|ICD9CM|PT|730.87|Other infections involving bone in diseases classified elsewhere, ankle and foot
C0158426|ICD9CM|AB|730.87|Bone infect NEC-ankle
C0158427|ICD9CM|PT|730.88|Other infections involving bone in diseases classified elsewhere, other specified sites
C0158427|ICD9CM|AB|730.88|Bone infect NEC-oth site
C0158428|ICD9CM|PT|730.89|Other infections involving bone in diseases classified elsewhere, multiple sites
C0158428|ICD9CM|AB|730.89|Bone infect NEC-mult
C0158434|ICD9CM|PT|730.25|Unspecified osteomyelitis, pelvic region and thigh
C0158434|ICD9CM|PT|730.95|Unspecified infection of bone, pelvic region and thigh
C0158434|ICD9CM|AB|730.25|Osteomyelitis NOS-pelvis
C0158434|ICD9CM|AB|730.95|Bone infect NOS-pelvis
C0158437|ICD9CM|PT|730.98|Unspecified infection of bone, other specified sites
C0158437|ICD9CM|AB|730.98|Bone infect NOS-oth site
C0158438|ICD9CM|PT|730.99|Unspecified infection of bone, multiple sites
C0158438|ICD9CM|AB|730.99|Bone infect NOS-mult
C0158439|ICD9CM|PT|731.1|Osteitis deformans in diseases classified elsewhere
C0158439|ICD9CM|AB|731.1|Osteitis def in oth dis
C0158440|ICD9CM|PT|731.8|Other bone involvement in diseases classified elsewhere
C0158440|ICD9CM|AB|731.8|Bone involv in oth dis
C0158441|ICD9CM|PT|732.2|Nontraumatic slipped upper femoral epiphysis
C0158441|ICD9CM|AB|732.2|Femoral epiphysiolysis
C0158442|ICD9CM|PT|732.3|Juvenile osteochondrosis of upper extremity
C0158442|ICD9CM|AB|732.3|Juv osteochondrosis arm
C0158444|ICD9CM|PT|732.5|Juvenile osteochondrosis of foot
C0158444|ICD9CM|AB|732.5|Juv osteochondrosis foot
C0158445|ICD9CM|PT|732.6|Other juvenile osteochondrosis
C0158445|ICD9CM|AB|732.6|Juv osteochondrosis NEC
C0158447|ICD9CM|AB|733.02|Idiopathic osteoporosis
C0158447|ICD9CM|PT|733.02|Idiopathic osteoporosis
C0158449|ICD9CM|PT|733.41|Aseptic necrosis of head of humerus
C0158449|ICD9CM|AB|733.41|Aseptic necrosis humerus
C0158450|ICD9CM|PT|733.43|Aseptic necrosis of medial femoral condyle
C0158450|ICD9CM|AB|733.43|Asept necro femur condyl
C0158451|ICD9CM|PT|733.44|Aseptic necrosis of talus
C0158451|ICD9CM|AB|733.44|Aseptic necrosis talus
C0158452|ICD9CM|PT|733.49|Aseptic necrosis of bone, other
C0158452|ICD9CM|AB|733.49|Asept necrosis bone NEC
C0158453|ICD9CM|HT|733.8|Malunion and nonunion of fracture
C0158454|ICD9CM|AB|733.81|Malunion of fracture
C0158454|ICD9CM|PT|733.81|Malunion of fracture
C0158456|ICD9CM|PT|733.91|Arrest of bone development or growth
C0158456|ICD9CM|AB|733.91|Arrest of bone growth
C0158457|ICD9CM|HT|735|Acquired deformities of toe
C0158457|ICD9CM|PT|735.9|Unspecified acquired deformity of toe
C0158457|ICD9CM|AB|735.9|Acq deformity of toe NOS
C0158458|ICD9CM|PT|735.0|Hallux valgus (acquired)
C0158458|ICD9CM|AB|735.0|Hallux valgus
C0158461|ICD9CM|AB|736.74|Claw foot, acquired
C0158461|ICD9CM|PT|736.74|Claw foot, acquired
C0158461|ICD9CM|PT|735.5|Claw toe (acquired)
C0158461|ICD9CM|AB|735.5|Claw toe
C0158463|ICD9CM|HT|736|Other acquired deformities of limbs
C0158464|ICD9CM|HT|736.0|Acquired deformities of forearm, excluding fingers
C0158465|ICD9CM|PT|736.01|Cubitus valgus (acquired)
C0158465|ICD9CM|AB|736.01|Cubitus valgus
C0158466|ICD9CM|PT|736.02|Cubitus varus (acquired)
C0158466|ICD9CM|AB|736.02|Cubitus varus
C0158467|ICD9CM|PT|736.03|Valgus deformity of wrist (acquired)
C0158467|ICD9CM|AB|736.03|Valgus deformity wrist
C0158468|ICD9CM|PT|736.04|Varus deformity of wrist (acquired)
C0158468|ICD9CM|AB|736.04|Varus deformity wrist
C0158470|ICD9CM|PT|736.06|Claw hand (acquired)
C0158470|ICD9CM|AB|736.06|Claw hand
C0158471|ICD9CM|AB|736.07|Club hand, acquired
C0158471|ICD9CM|PT|736.07|Club hand, acquired
C0158472|ICD9CM|PT|736.09|Other acquired deformities of forearm, excluding fingers
C0158472|ICD9CM|AB|736.09|Forearm deformity NEC
C0158473|ICD9CM|AB|736.1|Mallet finger
C0158473|ICD9CM|PT|736.1|Mallet finger
C0158476|ICD9CM|AB|736.21|Boutonniere deformity
C0158476|ICD9CM|PT|736.21|Boutonniere deformity
C0158477|ICD9CM|AB|736.22|Swan-neck deformity
C0158477|ICD9CM|PT|736.22|Swan-neck deformity
C0158478|ICD9CM|PT|736.30|Unspecified acquired deformity of hip
C0158478|ICD9CM|HT|736.3|Acquired deformities of hip
C0158478|ICD9CM|AB|736.30|Acq hip deformity NOS
C0158480|ICD9CM|PT|736.31|Coxa valga (acquired)
C0158480|ICD9CM|AB|736.31|Coxa valga
C0158481|ICD9CM|PT|736.32|Coxa vara (acquired)
C0158481|ICD9CM|AB|736.32|Coxa vara
C0158482|ICD9CM|PT|736.39|Other acquired deformities of hip
C0158482|ICD9CM|AB|736.39|Acq hip deformity NEC
C0158483|ICD9CM|HT|736.4|Genu valgum or varum (acquired)
C0158484|ICD9CM|PT|736.41|Genu valgum (acquired)
C0158484|ICD9CM|AB|736.41|Genu valgum
C0158485|ICD9CM|PT|736.42|Genu varum (acquired)
C0158485|ICD9CM|AB|736.42|Genu varum
C0158486|ICD9CM|PT|736.5|Genu recurvatum (acquired)
C0158486|ICD9CM|AB|736.5|Genu recurvatum
C0158487|ICD9CM|PT|736.6|Other acquired deformities of knee
C0158487|ICD9CM|AB|736.6|Acq knee deformity NEC
C0158488|ICD9CM|HT|736.7|Other acquired deformities of ankle and foot
C0158488|ICD9CM|PT|736.79|Other acquired deformities of ankle and foot
C0158488|ICD9CM|AB|736.79|Acq ankle-foot def NEC
C0158489|ICD9CM|PT|736.71|Acquired equinovarus deformity
C0158489|ICD9CM|AB|736.71|Acq equinovarus
C0158490|ICD9CM|PT|736.72|Equinus deformity of foot, acquired
C0158490|ICD9CM|AB|736.72|Acq equinus deformity
C0158493|ICD9CM|PT|736.75|Cavovarus deformity of foot, acquired
C0158493|ICD9CM|AB|736.75|Acq cavovarus deformity
C0158494|ICD9CM|PT|736.76|Other acquired calcaneus deformity
C0158494|ICD9CM|AB|736.76|Calcaneus deformity NEC
C0158495|ICD9CM|HT|736.8|Acquired deformities of other parts of limbs
C0158497|ICD9CM|PT|737.0|Adolescent postural kyphosis
C0158497|ICD9CM|AB|737.0|Adoles postural kyphosis
C0158498|ICD9CM|AB|737.11|Radiation kyphosis
C0158498|ICD9CM|PT|737.11|Kyphosis due to radiation
C0158499|ICD9CM|AB|737.12|Postlaminectomy kyphosis
C0158499|ICD9CM|PT|737.12|Kyphosis, postlaminectomy
C0158500|ICD9CM|PT|737.21|Lordosis, postlaminectomy
C0158500|ICD9CM|AB|737.21|Postlaminectomy lordosis
C0158501|ICD9CM|PT|737.22|Other postsurgical lordosis
C0158501|ICD9CM|AB|737.22|Oth postsurgery lordosis
C0158502|ICD9CM|PT|737.31|Resolving infantile idiopathic scoliosis
C0158502|ICD9CM|AB|737.31|Resolv idiopath scolios
C0158503|ICD9CM|PT|737.32|Progressive infantile idiopathic scoliosis
C0158503|ICD9CM|AB|737.32|Progr idiopath scoliosis
C0158504|ICD9CM|PT|737.33|Scoliosis due to radiation
C0158504|ICD9CM|AB|737.33|Radiation scoliosis
C0158505|ICD9CM|AB|737.34|Thoracogenic scoliosis
C0158505|ICD9CM|PT|737.34|Thoracogenic scoliosis
C0158506|ICD9CM|HT|737.4|Curvature of spine associated with other conditions
C0158506|ICD9CM|AB|737.9|Curvature of spine NOS
C0158506|ICD9CM|PT|737.40|Curvature of spine, unspecified, associated with other conditions
C0158506|ICD9CM|PT|737.9|Unspecified curvature of spine
C0158506|ICD9CM|AB|737.40|Spin curv NOS in oth dis
C0158507|ICD9CM|PT|737.41|Kyphosis associated with other conditions
C0158507|ICD9CM|AB|737.41|Kyphosis in oth dis
C0158508|ICD9CM|PT|737.42|Lordosis associated with other conditions
C0158508|ICD9CM|AB|737.42|Lordosis in oth dis
C0158509|ICD9CM|PT|737.43|Scoliosis associated with other conditions
C0158509|ICD9CM|AB|737.43|Scoliosis in oth dis
C0158510|ICD9CM|HT|738|Other acquired musculoskeletal deformity
C0158511|ICD9CM|HT|738.1|Other acquired deformity of head
C0158512|ICD9CM|PT|738.2|Acquired deformity of neck
C0158512|ICD9CM|AB|738.2|Acq neck deformity
C0158514|ICD9CM|PT|738.5|Other acquired deformity of back or spine
C0158514|ICD9CM|AB|738.5|Other acq back deformity
C0158515|ICD9CM|PT|738.6|Acquired deformity of pelvis
C0158515|ICD9CM|AB|738.6|Acq pelvic deformity
C0158516|ICD9CM|AB|738.7|Cauliflower ear
C0158516|ICD9CM|PT|738.7|Cauliflower ear
C0158517|ICD9CM|PT|738.8|Acquired deformity of other specified site
C0158517|ICD9CM|AB|738.8|Acq deformity NEC
C0158530|ICD9CM|HT|740|Anencephalus and similar anomalies
C0158534|ICD9CM|AB|741.90|Spina bifida
C0158534|ICD9CM|HT|741.9|Spina bifida without mention of hydrocephalus
C0158534|ICD9CM|PT|741.90|Spina bifida without mention of hydrocephalus, unspecified region
C0158535|ICD9CM|PT|741.91|Spina bifida without mention of hydrocephalus, cervical region
C0158535|ICD9CM|AB|741.91|Spina bifida-cerv
C0158536|ICD9CM|PT|741.92|Spina bifida without mention of hydrocephalus, dorsal (thoracic) region
C0158536|ICD9CM|AB|741.92|Spina bifida-dorsal
C0158537|ICD9CM|PT|741.93|Spina bifida without mention of hydrocephalus, lumbar region
C0158537|ICD9CM|AB|741.93|Spina bifida-lumbar
C0158538|ICD9CM|HT|742|Other congenital anomalies of nervous system
C0158543|ICD9CM|PT|743.03|Cystic eyeball, congenital
C0158543|ICD9CM|AB|743.03|Congen cystic eyeball
C0158545|ICD9CM|PT|743.12|Microphthalmos associated with other anomalies of eye and adnexa
C0158545|ICD9CM|AB|743.12|Microphth w oth eye anom
C0158547|ICD9CM|PT|743.22|Buphthalmos associated with other ocular anomalies
C0158547|ICD9CM|AB|743.22|Buphthal w oth eye anom
C0158548|ICD9CM|HT|743.3|Congenital cataract and lens anomalies
C0158549|ICD9CM|PT|743.31|Congenital capsular and subcapsular cataract
C0158549|ICD9CM|AB|743.31|Capsular cataract
C0158551|ICD9CM|PT|743.33|Congenital nuclear cataract
C0158551|ICD9CM|AB|743.33|Nuclear cataract
C0158552|ICD9CM|PT|743.34|Total and subtotal cataract, congenital
C0158552|ICD9CM|AB|743.34|Cong tot/subtot cataract
C0158553|ICD9CM|PT|743.36|Congenital anomalies of lens shape
C0158553|ICD9CM|AB|743.36|Anomalies of lens shape
C0158554|ICD9CM|PT|743.39|Other congenital cataract and lens anomalies
C0158554|ICD9CM|AB|743.39|Cong catar/lens anom NEC
C0158555|ICD9CM|HT|743.4|Coloboma and other anomalies of anterior segment
C0158557|ICD9CM|PT|743.42|Corneal opacities, interfering with vision, congenital
C0158557|ICD9CM|AB|743.42|Cong cornea opac aff vis
C0158558|ICD9CM|PT|743.43|Other corneal opacities, congenital
C0158558|ICD9CM|AB|743.43|Cong corneal opacit NEC
C0158560|ICD9CM|PT|743.46|Other specified congenital anomalies of iris and ciliary body
C0158560|ICD9CM|AB|743.46|Anom iris & cil body NEC
C0158562|ICD9CM|PT|743.48|Multiple and combined congenital anomalies of anterior segment
C0158562|ICD9CM|AB|743.48|Mult anom anter seg-eye
C0158564|ICD9CM|AB|743.51|Vitreous anomalies
C0158564|ICD9CM|PT|743.51|Vitreous anomalies
C0158566|ICD9CM|PT|743.53|Chorioretinal degeneration, congenital
C0158566|ICD9CM|AB|743.53|Cong chorioretinal degen
C0158567|ICD9CM|PT|743.54|Congenital folds and cysts of posterior segment
C0158567|ICD9CM|AB|743.54|Cong fold/cyst post eye
C0158568|ICD9CM|PT|743.55|Congenital macular changes
C0158568|ICD9CM|AB|743.55|Cong macular change-eye
C0158571|ICD9CM|PT|743.59|Other congenital anomalies of posterior segment
C0158571|ICD9CM|AB|743.59|Post segmnt anom NEC-eye
C0158572|ICD9CM|HT|743.6|Congenital anomalies of eyelids, lacrimal system, and orbit
C0158575|ICD9CM|PT|743.63|Other specified congenital anomalies of eyelid
C0158575|ICD9CM|AB|743.63|Spec anom of eyelid NEC
C0158576|ICD9CM|PT|743.64|Specified congenital anomalies of lacrimal gland
C0158576|ICD9CM|AB|743.64|Spec lacrimal gland anom
C0158577|ICD9CM|PT|743.65|Specified congenital anomalies of lacrimal passages
C0158577|ICD9CM|AB|743.65|Spec lacrimal pass anom
C0158579|ICD9CM|PT|743.69|Other congenital anomalies of eyelids, lacrimal system, and orbit
C0158579|ICD9CM|AB|743.69|Anom eyelid/lacr/orb NEC
C0158581|ICD9CM|HT|744|Congenital anomalies of ear, face, and neck
C0158587|ICD9CM|PT|744.04|Anomalies of ear ossicles
C0158587|ICD9CM|AB|744.04|Anomalies ear ossicles
C0158589|ICD9CM|PT|744.09|Other anomalies of ear causing impairment of hearing
C0158589|ICD9CM|AB|744.09|Ear anom NEC/impair hear
C0158591|ICD9CM|PT|744.21|Absence of ear lobe, congenital
C0158591|ICD9CM|AB|744.21|Cong absence of ear lobe
C0158592|ICD9CM|PT|744.24|Specified anomalies of Eustachian tube
C0158592|ICD9CM|AB|744.24|Eustachian tube anom NEC
C0158595|ICD9CM|HT|744.4|Branchial cleft cyst or fistula; preauricular sinus
C0158598|ICD9CM|PT|744.46|Preauricular sinus or fistula
C0158598|ICD9CM|AB|744.46|Preauricular sinus/fistu
C0158599|ICD9CM|AB|744.47|Preauricular cyst
C0158599|ICD9CM|PT|744.47|Preauricular cyst
C0158606|ICD9CM|HT|745|Bulbus cordis anomalies and anomalies of cardiac septal closure
C0158608|ICD9CM|PT|745.19|Other transposition of great vessels
C0158608|ICD9CM|AB|745.19|Transpos great vess NEC
C0158609|ICD9CM|PT|745.8|Other bulbus cordis anomalies and anomalies of cardiac septal closure
C0158609|ICD9CM|AB|745.8|Septal closure anom NEC
C0158610|ICD9CM|PT|745.9|Unspecified defect of septal closure
C0158610|ICD9CM|AB|745.9|Septal closure anom NOS
C0158611|ICD9CM|HT|746|Other congenital anomalies of heart
C0158616|ICD9CM|PT|746.1|Tricuspid atresia and stenosis, congenital
C0158616|ICD9CM|AB|746.1|Cong tricusp atres/sten
C0158617|ICD9CM|PT|746.4|Congenital insufficiency of aortic valve
C0158617|ICD9CM|AB|746.4|Cong aorta valv insuffic
C0158618|ICD9CM|PT|746.5|Congenital mitral stenosis
C0158618|ICD9CM|AB|746.5|Congen mitral stenosis
C0158619|ICD9CM|PT|746.6|Congenital mitral insufficiency
C0158619|ICD9CM|AB|746.6|Cong mitral insufficienc
C0158621|ICD9CM|PT|746.81|Subaortic stenosis
C0158621|ICD9CM|AB|746.81|Cong subaortic stenosis
C0158623|ICD9CM|AB|746.85|Coronary artery anomaly
C0158623|ICD9CM|PT|746.85|Coronary artery anomaly
C0158625|ICD9CM|HT|747|Other congenital anomalies of circulatory system
C0158629|ICD9CM|AB|747.21|Anomalies of aortic arch
C0158629|ICD9CM|PT|747.21|Anomalies of aortic arch
C0158632|ICD9CM|AB|747.40|Great vein anomaly NOS
C0158632|ICD9CM|HT|747.4|Anomalies of great veins, congenital
C0158632|ICD9CM|PT|747.40|Anomaly of great veins, unspecified
C0158634|ICD9CM|PT|747.42|Partial anomalous pulmonary venous connection
C0158634|ICD9CM|AB|747.42|Part anom pulm ven conn
C0158635|ICD9CM|PT|747.5|Absence or hypoplasia of umbilical artery
C0158635|ICD9CM|AB|747.5|Umbilical artery absence
C0158638|ICD9CM|PT|747.81|Anomalies of cerebrovascular system
C0158638|ICD9CM|AB|747.81|Cerebrovascular anomaly
C0158641|ICD9CM|AB|748.4|Congenital cystic lung
C0158641|ICD9CM|PT|748.4|Congenital cystic lung
C0158644|ICD9CM|AB|748.60|Lung anomaly NOS
C0158644|ICD9CM|PT|748.60|Anomaly of lung, unspecified
C0158646|ICD9CM|HT|749.2|Cleft palate with cleft lip
C0158646|ICD9CM|HT|749|Cleft palate and cleft lip
C0158646|ICD9CM|AB|749.20|Cleft palate & lip NOS
C0158646|ICD9CM|PT|749.20|Cleft palate with cleft lip, unspecified
C0158647|ICD9CM|PT|749.01|Cleft palate, unilateral, complete
C0158647|ICD9CM|AB|749.01|Unilat cleft palate-comp
C0158648|ICD9CM|PT|749.02|Cleft palate, unilateral, incomplete
C0158648|ICD9CM|AB|749.02|Unilat cleft palate-inc
C0158649|ICD9CM|PT|749.03|Cleft palate, bilateral, complete
C0158649|ICD9CM|AB|749.03|Bilat cleft palate-compl
C0158650|ICD9CM|PT|749.04|Cleft palate, bilateral, incomplete
C0158650|ICD9CM|AB|749.04|Bilat cleft palate-inc
C0158651|ICD9CM|PT|749.11|Cleft lip, unilateral, complete
C0158651|ICD9CM|AB|749.11|Unilat cleft lip-compl
C0158652|ICD9CM|PT|749.12|Cleft lip, unilateral, incomplete
C0158652|ICD9CM|AB|749.12|Unilat cleft lip-imcompl
C0158653|ICD9CM|PT|749.13|Cleft lip, bilateral, complete
C0158653|ICD9CM|AB|749.13|Bilat cleft lip-complete
C0158654|ICD9CM|PT|749.14|Cleft lip, bilateral, incomplete
C0158654|ICD9CM|AB|749.14|Bilat cleft lip-incompl
C0158655|ICD9CM|PT|749.21|Cleft palate with cleft lip, unilateral, complete
C0158655|ICD9CM|AB|749.21|Unil cleft palat/lip-com
C0158656|ICD9CM|PT|749.22|Cleft palate with cleft lip, unilateral, incomplete
C0158656|ICD9CM|AB|749.22|Unil cleft palat/lip-inc
C0158657|ICD9CM|PT|749.23|Cleft palate with cleft lip, bilateral, complete
C0158657|ICD9CM|AB|749.23|Bilat clft palat/lip-com
C0158658|ICD9CM|PT|749.24|Cleft palate with cleft lip, bilateral, incomplete
C0158658|ICD9CM|AB|749.24|Bilat clft palat/lip-inc
C0158659|ICD9CM|PT|749.25|Other combinations of cleft palate with cleft lip
C0158659|ICD9CM|AB|749.25|Cleft palate & lip NEC
C0158662|ICD9CM|PT|750.10|Congenital anomaly of tongue, unspecified
C0158662|ICD9CM|AB|750.10|Tongue anomaly NOS
C0158663|ICD9CM|AB|750.11|Aglossia
C0158663|ICD9CM|PT|750.11|Aglossia
C0158664|ICD9CM|PT|750.12|Congenital adhesions of tongue
C0158664|ICD9CM|AB|750.12|Cong adhesions of tongue
C0158667|ICD9CM|AB|750.21|Salivary gland absence
C0158667|ICD9CM|PT|750.21|Absence of salivary gland
C0158669|ICD9CM|PT|750.24|Congenital fistula of salivary gland
C0158669|ICD9CM|AB|750.24|Cong salivary fistula
C0158670|ICD9CM|PT|750.25|Congenital fistula of lip
C0158670|ICD9CM|AB|750.25|Congenital lip fistula
C0158671|ICD9CM|PT|750.26|Other specified anomalies of mouth
C0158671|ICD9CM|AB|750.26|Mouth anomaly NEC
C0158673|ICD9CM|PT|750.29|Other specified anomalies of pharynx
C0158673|ICD9CM|AB|750.29|Pharyngeal anomaly NEC
C0158674|ICD9CM|AB|750.6|Congenital hiatus hernia
C0158674|ICD9CM|PT|750.6|Congenital hiatus hernia
C0158678|ICD9CM|HT|751|Other congenital anomalies of digestive system
C0158679|ICD9CM|PT|751.4|Anomalies of intestinal fixation
C0158679|ICD9CM|AB|751.4|Intestinal fixation anom
C0158681|ICD9CM|HT|751.6|Anomalies of gallbladder, bile ducts, and liver
C0158684|ICD9CM|PT|751.7|Anomalies of pancreas
C0158684|ICD9CM|AB|751.7|Pancreas anomalies
C0158687|ICD9CM|HT|752|Congenital anomalies of genital organs
C0158687|ICD9CM|PT|752.9|Unspecified anomaly of genital organs
C0158687|ICD9CM|AB|752.9|Genital organ anom NOS
C0158688|ICD9CM|AB|752.0|Anomalies of ovaries
C0158688|ICD9CM|PT|752.0|Anomalies of ovaries
C0158689|ICD9CM|HT|752.1|Anomalies of fallopian tubes and broad ligaments, congenital
C0158689|ICD9CM|PT|752.10|Unspecified anomaly of fallopian tubes and broad ligaments
C0158689|ICD9CM|AB|752.10|Tubal/broad lig anom NOS
C0158694|ICD9CM|HT|752.4|Anomalies of cervix, vagina, and external female genitalia, congenital
C0158694|ICD9CM|PT|752.40|Unspecified anomaly of cervix, vagina, and external female genitalia
C0158694|ICD9CM|AB|752.40|Cervix/fem gen anom NOS
C0158695|ICD9CM|PT|752.41|Embryonic cyst of cervix, vagina, and external female genitalia
C0158695|ICD9CM|AB|752.41|Embryon cyst fem gen NEC
C0158698|ICD9CM|HT|753|Congenital anomalies of urinary system
C0158698|ICD9CM|PT|753.9|Unspecified anomaly of urinary system
C0158698|ICD9CM|AB|753.9|Urinary anomaly NOS
C0158699|ICD9CM|PT|753.0|Renal agenesis and dysgenesis
C0158699|ICD9CM|AB|753.0|Renal agenesis
C0158707|ICD9CM|PT|753.8|Other specified anomalies of bladder and urethra
C0158707|ICD9CM|AB|753.8|Cystourethral anom NEC
C0158709|ICD9CM|HT|754|Certain congenital musculoskeletal deformities
C0158712|ICD9CM|PT|754.2|Congenital musculoskeletal deformities of spine
C0158712|ICD9CM|AB|754.2|Cong postural deformity
C0158713|ICD9CM|PT|754.31|Congenital dislocation of hip, bilateral
C0158713|ICD9CM|AB|754.31|Congen hip disloc, bilat
C0158715|ICD9CM|PT|754.33|Congenital subluxation of hip, bilateral
C0158715|ICD9CM|AB|754.33|Cong hip sublux, bilat
C0158716|ICD9CM|PT|754.35|Congenital dislocation of one hip with subluxation of other hip
C0158716|ICD9CM|AB|754.35|Cong hip disloc w sublux
C0158718|ICD9CM|PT|754.41|Congenital dislocation of knee (with genu recurvatum)
C0158718|ICD9CM|AB|754.41|Cong knee dislocation
C0158719|ICD9CM|PT|754.42|Congenital bowing of femur
C0158719|ICD9CM|AB|754.42|Congen bowing of femur
C0158720|ICD9CM|PT|754.43|Congenital bowing of tibia and fibula
C0158720|ICD9CM|AB|754.43|Cong bowing tibia/fibula
C0158722|ICD9CM|HT|754.5|Varus deformities of feet, congenital
C0158722|ICD9CM|AB|754.50|Talipes varus
C0158722|ICD9CM|PT|754.50|Talipes varus
C0158725|ICD9CM|PT|754.59|Other varus deformities of feet
C0158725|ICD9CM|AB|754.59|Cong varus foot def NEC
C0158726|ICD9CM|HT|754.6|Valgus deformities of feet, congenital
C0158728|ICD9CM|PT|754.69|Other valgus deformities of feet
C0158728|ICD9CM|AB|754.69|Cong valgus foot def NEC
C0158729|ICD9CM|HT|754.7|Other congenital deformities of feet
C0158729|ICD9CM|PT|754.79|Other deformities of feet
C0158729|ICD9CM|AB|754.79|Cong foot deform NEC
C0158730|ICD9CM|HT|754.8|Other specified nonteratogenic anomalies
C0158730|ICD9CM|PT|754.89|Other specified nonteratogenic anomalies
C0158730|ICD9CM|AB|754.89|Nonteratogenic anom NEC
C0158731|ICD9CM|AB|754.82|Pectus carinatum
C0158731|ICD9CM|PT|754.82|Pectus carinatum
C0158732|ICD9CM|HT|755|Other congenital anomalies of limbs
C0158733|ICD9CM|PT|755.01|Polydactyly of fingers
C0158733|ICD9CM|AB|755.01|Polydactyly, fingers
C0158734|ICD9CM|PT|755.02|Polydactyly of toes
C0158734|ICD9CM|AB|755.02|Polydactyly, toes
C0158736|ICD9CM|PT|755.12|Syndactyly of fingers with fusion of bone
C0158736|ICD9CM|AB|755.12|Syndactyl fing w fusion
C0158738|ICD9CM|PT|755.14|Syndactyly of toes with fusion of bone
C0158738|ICD9CM|AB|755.14|Syndactyl toe w fusion
C0158743|ICD9CM|PT|755.23|Longitudinal deficiency, combined, involving humerus, radius, and ulna (complete or incomplete)
C0158743|ICD9CM|AB|755.23|Combin longit defic arm
C0158744|ICD9CM|PT|755.24|Longitudinal deficiency, humeral, complete or partial (with or without distal deficiencies, incomplete)
C0158744|ICD9CM|AB|755.24|Longitudin defic humerus
C0158745|ICD9CM|PT|755.25|Longitudinal deficiency, radioulnar, complete or partial (with or without distal deficiencies, incomplete)
C0158745|ICD9CM|AB|755.25|Longitud defic radioulna
C0158746|ICD9CM|PT|755.26|Longitudinal deficiency, radial, complete or partial (with or without distal deficiencies, incomplete)
C0158746|ICD9CM|AB|755.26|Longitud defic radius
C0158747|ICD9CM|PT|755.27|Longitudinal deficiency, ulnar, complete or partial (with or without distal deficiencies, incomplete)
C0158747|ICD9CM|AB|755.27|Longitudinal defic ulna
C0158748|ICD9CM|PT|755.28|Longitudinal deficiency, carpals or metacarpals, complete or partial (with or without incomplete phalangeal deficiency)
C0158748|ICD9CM|AB|755.28|Longitudinal defic hand
C0158752|ICD9CM|PT|755.31|Transverse deficiency of lower limb
C0158752|ICD9CM|AB|755.31|Transverse defic leg
C0158754|ICD9CM|PT|755.33|Longitudinal deficiency, combined, involving femur, tibia, and fibula (complete or incomplete)
C0158754|ICD9CM|AB|755.33|Comb longitudin def leg
C0158755|ICD9CM|PT|755.34|Longitudinal deficiency, femoral, complete or partial (with or without distal deficiencies, incomplete)
C0158755|ICD9CM|AB|755.34|Longitudinal defic femur
C0158756|ICD9CM|PT|755.35|Longitudinal deficiency, tibiofibular, complete or partial (with or without distal deficiencies, incomplete)
C0158756|ICD9CM|AB|755.35|Tibiofibula longit defic
C0158757|ICD9CM|PT|755.36|Longitudinal deficiency, tibia, complete or partial (with or without distal deficiencies, incomplete)
C0158757|ICD9CM|AB|755.36|Longitudinal defic tibia
C0158758|ICD9CM|PT|755.37|Longitudinal deficiency, fibular, complete or partial (with or without distal deficiencies, incomplete)
C0158758|ICD9CM|AB|755.37|Longitudin defic fibula
C0158759|ICD9CM|PT|755.38|Longitudinal deficiency, tarsals or metatarsals, complete or partial (with or without incomplete phalangeal deficiency)
C0158759|ICD9CM|AB|755.38|Longitudinal defic foot
C0158760|ICD9CM|PT|755.51|Congenital deformity of clavicle
C0158760|ICD9CM|AB|755.51|Cong deformity-clavicle
C0158761|ICD9CM|AB|755.53|Radioulnar synostosis
C0158761|ICD9CM|PT|755.53|Radioulnar synostosis
C0158763|ICD9CM|AB|755.57|Macrodactylia (fingers)
C0158763|ICD9CM|PT|755.57|Macrodactylia (fingers)
C0158767|ICD9CM|PT|755.64|Congenital deformity of knee (joint)
C0158767|ICD9CM|AB|755.64|Cong knee deformity
C0158768|ICD9CM|AB|755.65|Macrodactylia of toes
C0158768|ICD9CM|PT|755.65|Macrodactylia of toes
C0158773|ICD9CM|HT|756|Other congenital musculoskeletal anomalies
C0158775|ICD9CM|HT|756.1|Anomalies of spine, congenital
C0158775|ICD9CM|AB|756.10|Anomaly of spine NOS
C0158775|ICD9CM|PT|756.10|Anomaly of spine, unspecified
C0158776|ICD9CM|PT|756.13|Absence of vertebra, congenital
C0158776|ICD9CM|AB|756.13|Cong absence of vertebra
C0158779|ICD9CM|AB|756.2|Cervical rib
C0158779|ICD9CM|PT|756.2|Cervical rib
C0158782|ICD9CM|AB|756.6|Anomalies of diaphragm
C0158782|ICD9CM|PT|756.6|Anomalies of diaphragm
C0158784|ICD9CM|AB|756.82|Accessory muscle
C0158784|ICD9CM|PT|756.82|Accessory muscle
C0158794|ICD9CM|PT|758.4|Balanced autosomal translocation in normal individual
C0158794|ICD9CM|AB|758.4|Balance autosom transloc
C0158795|ICD9CM|HT|759|Other and unspecified congenital anomalies
C0158797|ICD9CM|AB|759.1|Adrenal gland anomaly
C0158797|ICD9CM|PT|759.1|Anomalies of adrenal gland
C0158799|ICD9CM|HT|760|Fetus or newborn affected by maternal conditions which may be unrelated to present pregnancy
C0158801|ICD9CM|PT|760.1|Maternal renal and urinary tract diseases affecting fetus or newborn
C0158801|ICD9CM|AB|760.1|Matern urine dis aff NB
C0158803|ICD9CM|PT|760.3|Other chronic maternal circulatory and respiratory diseases affecting fetus or newborn
C0158803|ICD9CM|AB|760.3|Matern cardioresp aff NB
C0158804|ICD9CM|PT|760.4|Maternal nutritional disorders affecting fetus or newborn
C0158804|ICD9CM|AB|760.4|Matern nutrit dis aff NB
C0158805|ICD9CM|PT|760.5|Maternal injury affecting fetus or newborn
C0158805|ICD9CM|AB|760.5|Maternal injury aff NB
C0158808|ICD9CM|PT|760.70|Unspecified noxious substance affecting fetus or newborn via placenta or breast milk
C0158808|ICD9CM|AB|760.70|Nox sub NOS aff NB/fetus
C0158809|ICD9CM|PT|760.72|Narcotics affecting fetus or newborn via placenta or breast milk
C0158809|ICD9CM|AB|760.72|Matern narc aff NB/fetus
C0158810|ICD9CM|PT|760.73|Hallucinogenic agents affecting fetus or newborn via placenta or breast milk
C0158810|ICD9CM|AB|760.73|Matern halluc af NB/fet
C0158811|ICD9CM|PT|760.74|Anti-infectives affecting fetus or newborn via placenta or breast milk
C0158811|ICD9CM|AB|760.74|Mat anti-inf aff NB/fet
C0158812|ICD9CM|PT|760.75|Cocaine affecting fetus or newborn via placenta or breast milk
C0158812|ICD9CM|AB|760.75|Mat cocaine aff NB/fet
C0158813|ICD9CM|PT|760.79|Other noxious influences affecting fetus or newborn via placenta or breast milk
C0158813|ICD9CM|AB|760.79|Nox sub NEC aff NB/fetus
C0158814|ICD9CM|PT|760.8|Other specified maternal conditions affecting fetus or newborn
C0158814|ICD9CM|AB|760.8|Maternal cond NEC aff NB
C0158816|ICD9CM|HT|761|Fetus or newborn affected by maternal complications of pregnancy
C0158816|ICD9CM|PT|761.9|Unspecified maternal complication of pregnancy affecting fetus or newborn
C0158816|ICD9CM|AB|761.9|Matern compl NOS aff NB
C0158817|ICD9CM|PT|761.0|Incompetent cervix affecting fetus or newborn
C0158817|ICD9CM|AB|761.0|Incompetnt cervix aff NB
C0158819|ICD9CM|PT|761.2|Oligohydramnios affecting fetus or newborn
C0158819|ICD9CM|AB|761.2|Oligohydramnios aff NB
C0158820|ICD9CM|PT|761.3|Polyhydramnios affecting fetus or newborn
C0158820|ICD9CM|AB|761.3|Polyhydramnios aff NB
C0158823|ICD9CM|PT|761.6|Maternal death affecting fetus or newborn
C0158823|ICD9CM|AB|761.6|Maternal death aff NB
C0158825|ICD9CM|PT|761.8|Other specified maternal complications of pregnancy affecting fetus or newborn
C0158825|ICD9CM|AB|761.8|Matern compl NEC aff NB
C0158829|ICD9CM|PT|762.1|Other forms of placental separation and hemorrhage affecting fetus or newborn
C0158829|ICD9CM|AB|762.1|Placenta hem NEC aff NB
C0158831|ICD9CM|PT|762.3|Placental transfusion syndromes affecting fetus or newborn
C0158831|ICD9CM|AB|762.3|Placent transfusion syn
C0158832|ICD9CM|PT|762.4|Prolapsed umbilical cord affecting fetus or newborn
C0158832|ICD9CM|AB|762.4|Prolapsed cord aff NB
C0158835|ICD9CM|PT|762.7|Chorioamnionitis affecting fetus or newborn
C0158835|ICD9CM|AB|762.7|Chorioamnionitis aff NB
C0158836|ICD9CM|PT|762.8|Other specified abnormalities of chorion and amnion affecting fetus or newborn
C0158836|ICD9CM|AB|762.8|Abn amnion NEC aff NB
C0158837|ICD9CM|PT|762.9|Unspecified abnormality of chorion and amnion affecting fetus or newborn
C0158837|ICD9CM|AB|762.9|Abn amnion NOS aff NB
C0158839|ICD9CM|PT|763.0|Breech delivery and extraction affecting fetus or newborn
C0158839|ICD9CM|AB|763.0|Breech del/extrac aff NB
C0158841|ICD9CM|PT|763.2|Forceps delivery affecting fetus or newborn
C0158841|ICD9CM|AB|763.2|Forceps delivery aff NB
C0158842|ICD9CM|PT|763.3|Delivery by vacuum extractor affecting fetus or newborn
C0158842|ICD9CM|AB|763.3|Vacuum extrac del aff NB
C0158843|ICD9CM|PT|763.4|Cesarean delivery affecting fetus or newborn
C0158843|ICD9CM|AB|763.4|Cesarean delivery aff NB
C0158845|ICD9CM|PT|763.6|Precipitate delivery affecting fetus or newborn
C0158845|ICD9CM|AB|763.6|Precipitate del aff NB
C0158846|ICD9CM|PT|763.7|Abnormal uterine contractions affecting fetus or newborn
C0158846|ICD9CM|AB|763.7|Abn uterine contr aff NB
C0158849|ICD9CM|HT|764|Slow fetal growth and fetal malnutrition
C0158851|ICD9CM|PT|764.00|"Light-for-dates" without mention of fetal malnutrition, unspecified [weight]
C0158851|ICD9CM|AB|764.00|Light-for-dates wtNOS
C0158852|ICD9CM|PT|764.01|"Light-for-dates" without mention of fetal malnutrition, less than 500 grams
C0158852|ICD9CM|AB|764.01|Light-for-dates <500g
C0158853|ICD9CM|PT|764.02|"Light-for-dates" without mention of fetal malnutrition, 500-749 grams
C0158853|ICD9CM|AB|764.02|Lt-for-dates 500-749g
C0158854|ICD9CM|PT|764.03|"Light-for-dates" without mention of fetal malnutrition, 750-999 grams
C0158854|ICD9CM|AB|764.03|Lt-for-dates 750-999g
C0158855|ICD9CM|PT|764.04|"Light-for-dates" without mention of fetal malnutrition, 1,000- 1,249 grams
C0158855|ICD9CM|AB|764.04|Lt-for-dates 1000-1249g
C0158856|ICD9CM|PT|764.05|"Light-for-dates"without mention of fetal malnutrition, 1,250- 1,499 grams
C0158856|ICD9CM|AB|764.05|Lt-for-dates 1250-1499g
C0158857|ICD9CM|PT|764.06|"Light-for-dates" without mention of fetal malnutrition, 1,500- 1,749 grams
C0158857|ICD9CM|AB|764.06|Lt-for-dates 1500-1749g
C0158858|ICD9CM|PT|764.07|"Light-for-dates" without mention of fetal malnutrition, 1,750- 1,999 grams
C0158858|ICD9CM|AB|764.07|Lt-for-dates 1750-1999g
C0158859|ICD9CM|PT|764.08|"Light-for-dates" without mention of fetal malnutrition, 2,000- 2,499 grams
C0158859|ICD9CM|AB|764.08|Lt-for-dates 2000-2499g
C0158860|ICD9CM|PT|764.09|"Light-for-dates" without mention of fetal malnutrition, 2,500 grams and over
C0158860|ICD9CM|AB|764.09|Lt-for-dates 2500+g
C0158861|ICD9CM|HT|764.1|"Light-for-dates" with signs of fetal malnutrition
C0158862|ICD9CM|PT|764.10|"Light-for-dates" with signs of fetal malnutrition, unspecified [weight]
C0158862|ICD9CM|AB|764.10|Lt-for-date w/mal wtNOS
C0158863|ICD9CM|PT|764.11|"Light-for-dates" with signs of fetal malnutrition, less than 500 grams
C0158863|ICD9CM|AB|764.11|Lt-for-date w/mal <500g
C0158864|ICD9CM|PT|764.12|"Light-for-dates"with signs of fetal malnutrition, 500-749 grams
C0158864|ICD9CM|AB|764.12|Lt-date w/mal 500-749g
C0158865|ICD9CM|PT|764.13|"Light-for-dates" with signs of fetal malnutrition, 750-999 grams
C0158865|ICD9CM|AB|764.13|Lt-date w/mal 750-999g
C0158866|ICD9CM|PT|764.14|"Light-for-dates" with signs of fetal malnutrition, 1,000-1,249 grams
C0158866|ICD9CM|AB|764.14|Lt-date w/mal 1000-1249g
C0158867|ICD9CM|PT|764.15|"Light-for-dates" with signs of fetal malnutrition, 1,250-1,499 grams
C0158867|ICD9CM|AB|764.15|Lt-date w/mal 1250-1499g
C0158868|ICD9CM|PT|764.16|"Light-for-dates" with signs of fetal malnutrition, 1,500-1,749 grams
C0158868|ICD9CM|AB|764.16|Lt-date w/mal 1500-1749g
C0158869|ICD9CM|PT|764.17|"Light-for-dates" with signs of fetal malnutrition, 1,750-1,999 grams
C0158869|ICD9CM|AB|764.17|Lt-date w/mal 1750-1999g
C0158870|ICD9CM|PT|764.18|"Light-for-dates"with signs of fetal malnutrition, 2,000-2,499 grams
C0158870|ICD9CM|AB|764.18|Lt-date w/mal 2000-2499g
C0158871|ICD9CM|PT|764.19|"Light-for-dates"with signs of fetal malnutrition, 2,500 grams and over
C0158871|ICD9CM|AB|764.19|Lt-for-date w/mal 2500+g
C0158872|ICD9CM|PT|764.20|Fetal malnutrition without mention of "light-for-dates", unspecified [weight]
C0158872|ICD9CM|AB|764.20|Fetal malnutrition wtNOS
C0158873|ICD9CM|PT|764.21|Fetal malnutrition without mention of "light-for-dates", less than 500 grams
C0158873|ICD9CM|AB|764.21|Fetal malnutrition <500g
C0158874|ICD9CM|PT|764.22|Fetal malnutrition without mention of "light-for-dates", 500-749 grams
C0158874|ICD9CM|AB|764.22|Fetal malnutr 500-749g
C0158875|ICD9CM|PT|764.23|Fetal malnutrition without mention of "light-for-dates", 750-999 grams
C0158875|ICD9CM|AB|764.23|Fetal mal 750-999g
C0158876|ICD9CM|PT|764.24|Fetal malnutrition without mention of "light-for-dates", 1,000-1,249 grams
C0158876|ICD9CM|AB|764.24|Fetal mal 1000-1249g
C0158877|ICD9CM|PT|764.25|Fetal malnutrition without mention of "light-for-dates", 1,250-1,499 grams
C0158877|ICD9CM|AB|764.25|Fetal mal 1250-1499g
C0158878|ICD9CM|PT|764.26|Fetal malnutrition without mention of "light-for-dates", 1,500-1,749 grams
C0158878|ICD9CM|AB|764.26|Fetal mal 1500-1749g
C0158879|ICD9CM|PT|764.27|Fetal malnutrition without mention of "light-for-dates", 1,750-1,999 grams
C0158879|ICD9CM|AB|764.27|Fetal malnutr 1750-1999g
C0158880|ICD9CM|PT|764.28|Fetal malnutrition without mention of "light-for-dates", 2,000-2,499 grams
C0158880|ICD9CM|AB|764.28|Fetal malnutr 2000-2499g
C0158881|ICD9CM|PT|764.29|Fetal malnutrition without mention of "light-for-dates", 2,500 grams and over
C0158881|ICD9CM|AB|764.29|Fetal malnutr 2500+g
C0158883|ICD9CM|PT|764.91|Fetal growth retardation, unspecified, less than 500 grams
C0158883|ICD9CM|AB|764.91|Fet growth retard <500g
C0158884|ICD9CM|PT|764.92|Fetal growth retardation, unspecified, 500-749 grams
C0158884|ICD9CM|AB|764.92|Fet growth ret 500-749g
C0158885|ICD9CM|PT|764.93|Fetal growth retardation, unspecified, 750-999 grams
C0158885|ICD9CM|AB|764.93|Fet growth ret 750-999g
C0158886|ICD9CM|PT|764.94|Fetal growth retardation, unspecified, 1,000-1,249 grams
C0158886|ICD9CM|AB|764.94|Fet grwth ret 1000-1249g
C0158887|ICD9CM|PT|764.95|Fetal growth retardation, unspecified, 1,250-1,499 grams
C0158887|ICD9CM|AB|764.95|Fet grwth ret 1250-1499g
C0158888|ICD9CM|PT|764.96|Fetal growth retardation, unspecified, 1,500-1,749 grams
C0158888|ICD9CM|AB|764.96|Fet grwth ret 1500-1749g
C0158889|ICD9CM|PT|764.97|Fetal growth retardation, unspecified, 1,750-1,999 grams
C0158889|ICD9CM|AB|764.97|Fet grwth ret 1750-1999g
C0158890|ICD9CM|PT|764.98|Fetal growth retardation, unspecified, 2,000-2,499 grams
C0158890|ICD9CM|AB|764.98|Fet grwth ret 2000-2499g
C0158891|ICD9CM|PT|764.99|Fetal growth retardation, unspecified, 2,500 grams and over
C0158891|ICD9CM|AB|764.99|Fet growth ret 2500+g
C0158892|ICD9CM|HT|765|Disorders relating to short gestation and unspecified low birthweight
C0158894|ICD9CM|PT|765.00|Extreme immaturity, unspecified [weight]
C0158894|ICD9CM|AB|765.00|Extreme immatur wtNOS
C0158895|ICD9CM|PT|765.01|Extreme immaturity, less than 500 grams
C0158895|ICD9CM|AB|765.01|Extreme immatur <500g
C0158896|ICD9CM|PT|765.02|Extreme immaturity, 500-749 grams
C0158896|ICD9CM|AB|765.02|Extreme immatur 500-749g
C0158897|ICD9CM|PT|765.03|Extreme immaturity, 750-999 grams
C0158897|ICD9CM|AB|765.03|Extreme immatur 750-999g
C0158898|ICD9CM|PT|765.04|Extreme immaturity, 1,000-1,249 grams
C0158898|ICD9CM|AB|765.04|Extreme immat 1000-1249g
C0158899|ICD9CM|PT|765.05|Extreme immaturity, 1,250-1,499 grams
C0158899|ICD9CM|AB|765.05|Extreme immat 1250-1499g
C0158900|ICD9CM|PT|765.06|Extreme immaturity, 1,500-1,749 grams
C0158900|ICD9CM|AB|765.06|Extreme immat 1500-1749g
C0158901|ICD9CM|PT|765.07|Extreme immaturity, 1,750-1,999 grams
C0158901|ICD9CM|AB|765.07|Extreme immat 1750-1999g
C0158902|ICD9CM|PT|765.08|Extreme immaturity, 2,000-2,499 grams
C0158902|ICD9CM|AB|765.08|Extreme immat 2000-2499g
C0158903|ICD9CM|PT|765.09|Extreme immaturity, 2,500 grams and over
C0158903|ICD9CM|AB|765.09|Extreme immat 2500+g
C0158905|ICD9CM|PT|765.11|Other preterm infants, less than 500 grams
C0158905|ICD9CM|AB|765.11|Preterm NEC <500g
C0158906|ICD9CM|PT|765.12|Other preterm infants, 500-749 grams
C0158906|ICD9CM|AB|765.12|Preterm NEC 500-749g
C0158907|ICD9CM|PT|765.13|Other preterm infants, 750-999 grams
C0158907|ICD9CM|AB|765.13|Preterm NEC 750-999g
C0158908|ICD9CM|PT|765.14|Other preterm infants, 1,000-1,249 grams
C0158908|ICD9CM|AB|765.14|Preterm NEC 1000-1249g
C0158909|ICD9CM|PT|765.15|Other preterm infants, 1,250-1,499 grams
C0158909|ICD9CM|AB|765.15|Preterm NEC 1250-1499g
C0158910|ICD9CM|PT|765.16|Other preterm infants, 1,500-1,749 grams
C0158910|ICD9CM|AB|765.16|Preterm NEC 1500-1749g
C0158911|ICD9CM|PT|765.17|Other preterm infants, 1,750-1,999 grams
C0158911|ICD9CM|AB|765.17|Preterm NEC 1750-1999g
C0158912|ICD9CM|PT|765.18|Other preterm infants, 2,000-2,499 grams
C0158912|ICD9CM|AB|765.18|Preterm NEC 2000-2499g
C0158913|ICD9CM|PT|765.19|Other preterm infants, 2,500 grams and over
C0158913|ICD9CM|AB|765.19|Preterm NEC 2500+g
C0158914|ICD9CM|HT|766|Disorders relating to long gestation and high birthweight
C0158917|ICD9CM|HT|766.2|Late infant, not "heavy-for-dates"
C0158925|ICD9CM|PT|767.7|Other cranial and peripheral nerve injuries due to birth trauma
C0158925|ICD9CM|AB|767.7|Nerve inj NEC at birth
C0158928|ICD9CM|PT|768.1|Fetal death from asphyxia or anoxia during labor
C0158928|ICD9CM|AB|768.1|Fet death-anoxia dur lab
C0158929|ICD9CM|PT|768.2|Fetal distress before onset of labor, in liveborn infant
C0158929|ICD9CM|AB|768.2|Fet distress befor labor
C0158931|ICD9CM|AB|768.5|Severe birth asphyxia
C0158931|ICD9CM|PT|768.5|Severe birth asphyxia
C0158934|ICD9CM|HT|770|Other respiratory conditions of fetus and newborn
C0158935|ICD9CM|AB|770.0|Congenital pneumonia
C0158935|ICD9CM|PT|770.0|Congenital pneumonia
C0158936|ICD9CM|PT|770.2|Interstitial emphysema and related conditions
C0158936|ICD9CM|AB|770.2|NB interstit emphysema
C0158939|ICD9CM|PT|770.5|Other and unspecified atelectasis
C0158939|ICD9CM|AB|770.5|NB atelectasis NEC/NOS
C0158940|ICD9CM|PT|770.6|Transitory tachypnea of newborn
C0158940|ICD9CM|AB|770.6|NB transitory tachypnea
C0158942|ICD9CM|HT|770.8|Other newborn respiratory problems
C0158944|ICD9CM|HT|771|Infections specific to the perinatal period
C0158945|ICD9CM|PT|771.1|Congenital cytomegalovirus infection
C0158945|ICD9CM|AB|771.1|Cong cytomegalovirus inf
C0158946|ICD9CM|PT|771.2|Other congenital infections specific to the perinatal period
C0158946|ICD9CM|AB|771.2|Congenital infec NEC
C0158947|ICD9CM|PT|771.4|Omphalitis of the newborn
C0158947|ICD9CM|AB|771.4|Omphalitis of newborn
C0158948|ICD9CM|PT|771.5|Neonatal infective mastitis
C0158948|ICD9CM|AB|771.5|Neonatal infec mastitis
C0158950|ICD9CM|PT|771.89|Other infections specific to the perinatal period
C0158950|ICD9CM|HT|771.8|Other infection specific to the perinatal period
C0158950|ICD9CM|AB|771.89|Perinatal infection NEC
C0158951|ICD9CM|PT|772.0|Fetal blood loss
C0158951|ICD9CM|AB|772.0|NB fetal blood loss NEC
C0158956|ICD9CM|PT|772.4|Gastrointestinal hemorrhage of fetus or newborn
C0158956|ICD9CM|AB|772.4|NB GI hemorrhage
C0158957|ICD9CM|PT|772.5|Adrenal hemorrhage of fetus or newborn
C0158957|ICD9CM|AB|772.5|NB adrenal hemorrhage
C0158959|ICD9CM|PT|772.8|Other specified hemorrhage of fetus or newborn
C0158959|ICD9CM|AB|772.8|Neonatal hemorrhage NEC
C0158962|ICD9CM|PT|773.0|Hemolytic disease of fetus or newborn due to Rh isoimmunization
C0158962|ICD9CM|AB|773.0|NB hemolyt dis:rh isoimm
C0158967|ICD9CM|PT|773.5|Late anemia of fetus or newborn due to isoimmunization
C0158967|ICD9CM|AB|773.5|NB late anemia:isoimmun
C0158968|ICD9CM|HT|774|Other perinatal jaundice
C0158969|ICD9CM|PT|774.0|Perinatal jaundice from hereditary hemolytic anemias
C0158969|ICD9CM|AB|774.0|Perinat jaund-hered anem
C0158971|ICD9CM|PT|774.2|Neonatal jaundice associated with preterm delivery
C0158971|ICD9CM|AB|774.2|Neonat jaund preterm del
C0158972|ICD9CM|HT|774.3|Neonatal jaundice due to delayed conjugation from other causes
C0158974|ICD9CM|PT|774.31|Neonatal jaundice due to delayed conjugation in diseases classified elsewhere
C0158974|ICD9CM|AB|774.31|Neonat jaund in oth dis
C0158975|ICD9CM|PT|774.39|Other neonatal jaundice due to delayed conjugation from other causes
C0158975|ICD9CM|AB|774.39|Delay conjugat jaund NEC
C0158976|ICD9CM|PT|774.4|Perinatal jaundice due to hepatocellular damage
C0158976|ICD9CM|AB|774.4|Fetal/neonatal hepatitis
C0158977|ICD9CM|PT|774.5|Perinatal jaundice from other causes
C0158977|ICD9CM|AB|774.5|Perinatal jaundice NEC
C0158978|ICD9CM|PT|774.7|Kernicterus of fetus or newborn not due to isoimmunization
C0158978|ICD9CM|AB|774.7|NB kernicterus
C0158979|ICD9CM|HT|775|Endocrine and metabolic disturbances specific to the fetus and newborn
C0158981|ICD9CM|PT|775.1|Neonatal diabetes mellitus
C0158981|ICD9CM|AB|775.1|Neonat diabetes mellitus
C0158982|ICD9CM|PT|775.2|Neonatal myasthenia gravis
C0158982|ICD9CM|AB|775.2|Neonat myasthenia gravis
C0158983|ICD9CM|AB|775.3|Neonatal thyrotoxicosis
C0158983|ICD9CM|PT|775.3|Neonatal thyrotoxicosis
C0158984|ICD9CM|PT|775.4|Hypocalcemia and hypomagnesemia of newborn
C0158984|ICD9CM|AB|775.4|Hypocalcem/hypomagnes NB
C0158986|ICD9CM|AB|775.6|Neonatal hypoglycemia
C0158986|ICD9CM|PT|775.6|Neonatal hypoglycemia
C0158987|ICD9CM|PT|775.7|Late metabolic acidosis of newborn
C0158987|ICD9CM|AB|775.7|Late metab acidosis NB
C0158989|ICD9CM|PT|775.9|Unspecified endocrine and metabolic disturbances specific to the fetus and newborn
C0158989|ICD9CM|AB|775.9|Transient met dis NB NOS
C0158991|ICD9CM|PT|776.1|Transient neonatal thrombocytopenia
C0158991|ICD9CM|AB|776.1|Neonatal thrombocytopen
C0158992|ICD9CM|PT|776.2|Disseminated intravascular coagulation in newborn
C0158992|ICD9CM|AB|776.2|Dissem intravasc coag NB
C0158993|ICD9CM|PT|776.3|Other transient neonatal disorders of coagulation
C0158993|ICD9CM|AB|776.3|Oth neonatal coag dis
C0158995|ICD9CM|AB|776.5|Congenital anemia
C0158995|ICD9CM|PT|776.5|Congenital anemia
C0158996|ICD9CM|AB|776.6|Anemia of prematurity
C0158996|ICD9CM|PT|776.6|Anemia of prematurity
C0158997|ICD9CM|PT|776.7|Transient neonatal neutropenia
C0158997|ICD9CM|AB|776.7|Neonatal neutropenia
C0158998|ICD9CM|PT|776.8|Other specified transient hematological disorders of fetus or newborn
C0158998|ICD9CM|AB|776.8|Transient hemat dis NEC
C0158999|ICD9CM|PT|776.9|Unspecified hematological disorder specific to newborn
C0158999|ICD9CM|AB|776.9|NB hematological dis NOS
C0159000|ICD9CM|HT|777|Perinatal disorders of digestive system
C0159000|ICD9CM|PT|777.9|Unspecified perinatal disorder of digestive system
C0159000|ICD9CM|AB|777.9|Perinat GI sys dis NOS
C0159004|ICD9CM|PT|777.4|Transitory ileus of newborn
C0159004|ICD9CM|AB|777.4|Transitory ileus of NB
C0159006|ICD9CM|PT|777.6|Perinatal intestinal perforation
C0159006|ICD9CM|AB|777.6|Perinatal intest perfor
C0159007|ICD9CM|PT|777.8|Other specified perinatal disorders of digestive system
C0159007|ICD9CM|AB|777.8|Perinat GI sys dis NEC
C0159009|ICD9CM|HT|778|Conditions involving the integument and temperature regulation of fetus and newborn
C0159011|ICD9CM|PT|778.2|Cold injury syndrome of newborn
C0159011|ICD9CM|AB|778.2|NB cold injury syndrome
C0159012|ICD9CM|PT|778.3|Other hypothermia of newborn
C0159012|ICD9CM|AB|778.3|NB hypothermia NEC
C0159013|ICD9CM|PT|778.4|Other disturbances of temperature regulation of newborn
C0159013|ICD9CM|AB|778.4|NB temp regulat dis NEC
C0159014|ICD9CM|PT|778.5|Other and unspecified edema of newborn
C0159014|ICD9CM|AB|778.5|Edema of newborn NEC/NOS
C0159015|ICD9CM|AB|778.6|Congenital hydrocele
C0159015|ICD9CM|PT|778.6|Congenital hydrocele
C0159018|ICD9CM|PT|778.9|Unspecified condition involving the integument and temperature regulation of fetus and newborn
C0159018|ICD9CM|AB|778.9|NB integument cond NOS
C0159019|ICD9CM|HT|779|Other and ill-defined conditions originating in the perinatal period
C0159020|ICD9CM|AB|779.0|Convulsions in newborn
C0159020|ICD9CM|PT|779.0|Convulsions in newborn
C0159021|ICD9CM|PT|779.1|Other and unspecified cerebral irritability in newborn
C0159021|ICD9CM|AB|779.1|NB cereb irrit NEC/NOS
C0159022|ICD9CM|PT|779.2|Cerebral depression, coma, and other abnormal cerebral signs in fetus or newborn
C0159022|ICD9CM|AB|779.2|Cns dysfunction syn NB
C0159023|ICD9CM|PT|779.31|Feeding problems in newborn
C0159023|ICD9CM|AB|779.31|NB feeding problems
C0159027|ICD9CM|HT|779.8|Other specified conditions originating in the perinatal period
C0159027|ICD9CM|PT|779.89|Other specified conditions originating in the perinatal period
C0159027|ICD9CM|AB|779.89|Perinatal condition NEC
C0159028|ICD9CM|HT|780|General symptoms
C0159033|ICD9CM|HT|781|Symptoms involving nervous and musculoskeletal systems
C0159034|ICD9CM|AB|781.4|Transient limb paralysis
C0159034|ICD9CM|PT|781.4|Transient paralysis of limb
C0159036|ICD9CM|HT|781.9|Other symptoms involving nervous and musculoskeletal systems
C0159036|ICD9CM|PT|781.99|Other symptoms involving nervous and musculoskeletal systems
C0159036|ICD9CM|AB|781.99|Nerve/musculskel sym NEC
C0159037|ICD9CM|PT|782.9|Other symptoms involving skin and integumentary tissues
C0159037|ICD9CM|HT|782|Symptoms involving skin and other integumentary tissue
C0159037|ICD9CM|AB|782.9|Integument tiss symp NEC
C0159038|ICD9CM|HT|782.6|Pallor and flushing
C0159039|ICD9CM|AB|782.7|Spontaneous ecchymoses
C0159039|ICD9CM|PT|782.7|Spontaneous ecchymoses
C0159040|ICD9CM|AB|782.8|Changes in skin texture
C0159040|ICD9CM|PT|782.8|Changes in skin texture
C0159043|ICD9CM|PT|783.9|Other symptoms concerning nutrition, metabolism, and development
C0159043|ICD9CM|AB|783.9|Nutr/metab/devel sym NEC
C0159045|ICD9CM|PT|784.2|Swelling, mass, or lump in head and neck
C0159045|ICD9CM|AB|784.2|Swelling in head & neck
C0159047|ICD9CM|AB|784.60|Symbolic dysfunction NOS
C0159047|ICD9CM|PT|784.60|Symbolic dysfunction, unspecified
C0159049|ICD9CM|HT|785|Symptoms involving cardiovascular system
C0159050|ICD9CM|PT|785.3|Other abnormal heart sounds
C0159050|ICD9CM|AB|785.3|Abnorm heart sounds NEC
C0159051|ICD9CM|HT|785.5|Shock without mention of trauma
C0159053|ICD9CM|HT|786.0|Dyspnea and respiratory abnormalities
C0159054|ICD9CM|AB|786.4|Abnormal sputum
C0159054|ICD9CM|PT|786.4|Abnormal sputum
C0159055|ICD9CM|PT|786.6|Swelling, mass, or lump in chest
C0159055|ICD9CM|AB|786.6|Chest swelling/mass/lump
C0159056|ICD9CM|AB|786.7|Abnormal chest sounds
C0159056|ICD9CM|PT|786.7|Abnormal chest sounds
C0159057|ICD9CM|PT|786.9|Other symptoms involving respiratory system and chest
C0159057|ICD9CM|AB|786.9|Resp sys/chest symp NEC
C0159058|ICD9CM|HT|787|Symptoms involving digestive system
C0159059|ICD9CM|AB|787.4|Visible peristalsis
C0159059|ICD9CM|PT|787.4|Visible peristalsis
C0159060|ICD9CM|AB|787.5|Abnormal bowel sounds
C0159060|ICD9CM|PT|787.5|Abnormal bowel sounds
C0159061|ICD9CM|HT|787.9|Other symptoms involving digestive system
C0159061|ICD9CM|PT|787.99|Other symptoms involving digestive system
C0159061|ICD9CM|AB|787.99|Digestve syst symptm NEC
C0159063|ICD9CM|HT|788.6|Other abnormality of urination
C0159063|ICD9CM|PT|788.69|Other abnormality of urination
C0159063|ICD9CM|AB|788.69|Oth abnormalt urination
C0159064|ICD9CM|HT|788.9|Other symptoms involving urinary system
C0159064|ICD9CM|PT|788.99|Other symptoms involving urinary system
C0159064|ICD9CM|AB|788.99|Oth symptm urinary systm
C0159065|ICD9CM|HT|789|Other symptoms involving abdomen and pelvis
C0159065|ICD9CM|PT|789.9|Other symptoms involving abdomen and pelvis
C0159065|ICD9CM|AB|789.9|Abdomen/pelvis symp NEC
C0159066|ICD9CM|HT|789.4|Abdominal rigidity
C0159066|ICD9CM|PT|789.40|Abdominal rigidity, unspecified site
C0159066|ICD9CM|AB|789.40|Abdmnal rgdt unspcf site
C0159070|ICD9CM|PT|790.3|Excessive blood level of alcohol
C0159070|ICD9CM|AB|790.3|Excess blood-alcohol lev
C0159071|ICD9CM|PT|790.4|Nonspecific elevation of levels of transaminase or lactic acid dehydrogenase [LDH]
C0159071|ICD9CM|AB|790.4|Elev transaminase/ldh
C0159072|ICD9CM|PT|790.5|Other nonspecific abnormal serum enzyme levels
C0159072|ICD9CM|AB|790.5|Abn serum enzy level NEC
C0159073|ICD9CM|HT|790.9|Other nonspecific findings on examination of blood
C0159073|ICD9CM|PT|790.99|Other nonspecific findings on examination of blood
C0159073|ICD9CM|AB|790.99|Oth nspcf finding blood
C0159075|ICD9CM|AB|791.1|Chyluria
C0159075|ICD9CM|PT|791.1|Chyluria
C0159076|ICD9CM|AB|791.4|Biliuria
C0159076|ICD9CM|PT|791.4|Biliuria
C0159077|ICD9CM|PT|791.7|Other cells and casts in urine
C0159077|ICD9CM|AB|791.7|Oth cells/casts in urine
C0159078|ICD9CM|PT|791.9|Other nonspecific findings on examination of urine
C0159078|ICD9CM|AB|791.9|Abn urine findings NEC
C0159079|ICD9CM|PT|792.9|Other nonspecific abnormal findings in body substances
C0159079|ICD9CM|HT|792|Nonspecific abnormal findings in other body substances
C0159079|ICD9CM|AB|792.9|Abn find-body subst NEC
C0159084|ICD9CM|PT|792.4|Nonspecific abnormal findings in saliva
C0159084|ICD9CM|AB|792.4|Abn findings-saliva
C0159085|ICD9CM|HT|793|Nonspecific (abnormal) findings on radiological and other examination of body structure
C0159088|ICD9CM|PT|793.2|Nonspecific (abnormal) findings on radiological and other examination of other intrathoracic organs
C0159088|ICD9CM|AB|793.2|Nonsp abn intrathor NEC
C0159089|ICD9CM|PT|793.3|Nonspecific (abnormal) findings on radiological and other examination of biliary tract
C0159089|ICD9CM|AB|793.3|Nonsp abn fd-bilry tract
C0159090|ICD9CM|PT|793.4|Nonspecific (abnormal) findings on radiological and other examination of gastrointestinal tract
C0159090|ICD9CM|AB|793.4|Nonsp abn find-gi tract
C0159092|ICD9CM|PT|793.6|Nonspecific (abnormal) findings on radiological and other examination of abdominal area, including retroperitoneum
C0159092|ICD9CM|AB|793.6|Nonsp abn fnd-abdom area
C0159093|ICD9CM|PT|793.7|Nonspecific (abnormal) findings on radiological and other examination of musculoskeletal system
C0159093|ICD9CM|AB|793.7|Nonsp abn find-ms system
C0159094|ICD9CM|HT|793.8|Nonspecific abnormal findings on radiological and other examination of breast
C0159099|ICD9CM|PT|794.02|Nonspecific abnormal electroencephalogram [EEG]
C0159099|ICD9CM|AB|794.02|Abn electroencephalogram
C0159100|ICD9CM|PT|794.09|Other nonspecific abnormal results of function study of brain and central nervous system
C0159100|ICD9CM|AB|794.09|Abn cns funct study NEC
C0159102|ICD9CM|PT|794.10|Nonspecific abnormal response to nerve stimulation, unspecified
C0159102|ICD9CM|AB|794.10|Abn stimul response NOS
C0159104|ICD9CM|PT|794.12|Nonspecific abnormal electro-oculogram [EOG]
C0159104|ICD9CM|AB|794.12|Abnorm electro-oculogram
C0159106|ICD9CM|PT|794.14|Nonspecific abnormal oculomotor studies
C0159106|ICD9CM|AB|794.14|Abn oculomotor studies
C0159107|ICD9CM|PT|794.15|Nonspecific abnormal auditory function studies
C0159107|ICD9CM|AB|794.15|Abn auditory funct study
C0159110|ICD9CM|PT|794.19|Other nonspecific abnormal results of function study of peripheral nervous system and special senses
C0159110|ICD9CM|AB|794.19|Abn periph nerv stud NEC
C0159117|ICD9CM|PT|794.6|Nonspecific abnormal results of other endocrine function study
C0159117|ICD9CM|AB|794.6|Abn endocrine study NEC
C0159118|ICD9CM|PT|794.7|Nonspecific abnormal results of function study of basal metabolism
C0159118|ICD9CM|AB|794.7|Abn basal metabol study
C0159120|ICD9CM|PT|794.9|Nonspecific abnormal results of other specified function study
C0159120|ICD9CM|AB|794.9|Abn function study NEC
C0159125|ICD9CM|HT|795.3|Nonspecific positive culture findings
C0159126|ICD9CM|PT|795.4|Other nonspecific abnormal histological findings
C0159126|ICD9CM|AB|795.4|Abn histologic find NEC
C0159128|ICD9CM|PT|795.6|False positive serological test for syphilis
C0159128|ICD9CM|AB|795.6|False pos sero test-syph
C0159131|ICD9CM|HT|796|Other nonspecific abnormal findings
C0159131|ICD9CM|PT|796.9|Other nonspecific abnormal findings
C0159131|ICD9CM|AB|796.9|Abnormal findings NEC
C0159132|ICD9CM|PT|796.0|Nonspecific abnormal toxicological findings
C0159132|ICD9CM|AB|796.0|Abn toxicologic finding
C0159135|ICD9CM|PT|796.4|Other abnormal clinical findings
C0159135|ICD9CM|AB|796.4|Abn clinical finding NEC
C0159138|ICD9CM|HT|799|Other ill-defined and unknown causes of morbidity and mortality
C0159139|ICD9CM|HT|800|Fracture of vault of skull
C0159140|ICD9CM|HT|800.0|Closed fracture of vault of skull without mention of intracranial injury
C0159141|ICD9CM|PT|800.00|Closed fracture of vault of skull without mention of intracranial injury, unspecified state of consciousness
C0159141|ICD9CM|AB|800.00|Closed skull vault fx
C0159142|ICD9CM|PT|800.01|Closed fracture of vault of skull without mention of intracranial injury, with no loss of consciousness
C0159142|ICD9CM|AB|800.01|Cl skull vlt fx w/o coma
C0159143|ICD9CM|PT|800.02|Closed fracture of vault of skull without mention of intracranial injury, with brief [less than one hour] loss of consciousness
C0159143|ICD9CM|AB|800.02|Cl skull vlt fx-brf coma
C0159144|ICD9CM|PT|800.03|Closed fracture of vault of skull without mention of intracranial injury, with moderate [1-24 hours] loss of consciousness
C0159144|ICD9CM|AB|800.03|Cl skull vlt fx-mod coma
C0159145|ICD9CM|PT|800.04|Closed fracture of vault of skull without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159145|ICD9CM|AB|800.04|Cl skl vlt fx-proln coma
C0159146|ICD9CM|PT|800.05|Closed fracture of vault of skull without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159146|ICD9CM|AB|800.05|Cl skul vlt fx-deep coma
C0159147|ICD9CM|PT|800.06|Closed fracture of vault of skull without mention of intracranial injury, with loss of consciousness of unspecified duration
C0159147|ICD9CM|AB|800.06|Cl skull vlt fx-coma NOS
C0159148|ICD9CM|PT|800.09|Closed fracture of vault of skull without mention of intracranial injury, with concussion, unspecified
C0159148|ICD9CM|AB|800.09|Cl skl vlt fx-concus NOS
C0159149|ICD9CM|HT|800.1|Closed fracture of vault of skull with cerebral laceration and contusion
C0159150|ICD9CM|PT|800.10|Closed fracture of vault of skull with cerebral laceration and contusion, unspecified state of consciousness
C0159150|ICD9CM|AB|800.10|Cl skl vlt fx/cerebr lac
C0159151|ICD9CM|PT|800.11|Closed fracture of vault of skull with cerebral laceration and contusion, with no loss of consciousness
C0159151|ICD9CM|AB|800.11|Cl skull vlt fx w/o coma
C0159152|ICD9CM|PT|800.12|Closed fracture of vault of skull with cerebral laceration and contusion, with brief [less than one hour] loss of consciousness
C0159152|ICD9CM|AB|800.12|Cl skull vlt fx-brf coma
C0159153|ICD9CM|PT|800.13|Closed fracture of vault of skull with cerebral laceration and contusion, with moderate [1-24 hours] loss of consciousness
C0159153|ICD9CM|AB|800.13|Cl skull vlt fx-mod coma
C0159154|ICD9CM|PT|800.14|Closed fracture of vault of skull with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159154|ICD9CM|AB|800.14|Cl skl vlt fx-proln coma
C0159155|ICD9CM|PT|800.15|Closed fracture of vault of skull with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159155|ICD9CM|AB|800.15|Cl skul vlt fx-deep coma
C0159156|ICD9CM|PT|800.16|Closed fracture of vault of skull with cerebral laceration and contusion, with loss of consciousness of unspecified duration
C0159156|ICD9CM|AB|800.16|Cl skull vlt fx-coma NOS
C0159158|ICD9CM|HT|800.2|Closed fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage
C0159159|ICD9CM|PT|800.20|Closed fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, unspecified state of consciousness
C0159159|ICD9CM|AB|800.20|Cl skl vlt fx/mening hem
C0159160|ICD9CM|PT|800.21|Closed fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with no loss of consciousness
C0159160|ICD9CM|AB|800.21|Cl skull vlt fx w/o coma
C0159161|ICD9CM|PT|800.22|Closed fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with brief [less than one hour] loss of consciousness
C0159161|ICD9CM|AB|800.22|Cl skull vlt fx-brf coma
C0159162|ICD9CM|PT|800.23|Closed fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159162|ICD9CM|AB|800.23|Cl skull vlt fx-mod coma
C0159163|ICD9CM|PT|800.24|Closed fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159163|ICD9CM|AB|800.24|Cl skl vlt fx-proln coma
C0159164|ICD9CM|PT|800.25|Closed fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159164|ICD9CM|AB|800.25|Cl skul vlt fx-deep coma
C0159165|ICD9CM|PT|800.26|Closed fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with loss of consciousness of unspecified duration
C0159165|ICD9CM|AB|800.26|Cl skull vlt fx-coma NOS
C0159167|ICD9CM|HT|800.3|Closed fracture of vault of skull with other and unspecified intracranial hemorrhage
C0159168|ICD9CM|PT|800.30|Closed fracture of vault of skull with other and unspecified intracranial hemorrhage, unspecified state of consciousness
C0159168|ICD9CM|AB|800.30|Cl skull vlt fx/hem NEC
C0159169|ICD9CM|PT|800.31|Closed fracture of vault of skull with other and unspecified intracranial hemorrhage, with no loss of consciousness
C0159169|ICD9CM|AB|800.31|Cl skull vlt fx w/o coma
C0159170|ICD9CM|PT|800.32|Closed fracture of vault of skull with other and unspecified intracranial hemorrhage, with brief [less than one hour] loss of consciousness
C0159170|ICD9CM|AB|800.32|Cl skull vlt fx-brf coma
C0159171|ICD9CM|PT|800.33|Closed fracture of vault of skull with other and unspecified intracranial hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159171|ICD9CM|AB|800.33|Cl skull vlt fx-mod coma
C0159172|ICD9CM|PT|800.34|Closed fracture of vault of skull with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159172|ICD9CM|AB|800.34|Cl skl vlt fx-proln coma
C0159173|ICD9CM|PT|800.35|Closed fracture of vault of skull with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159173|ICD9CM|AB|800.35|Cl skul vlt fx-deep coma
C0159174|ICD9CM|PT|800.36|Closed fracture of vault of skull with other and unspecified intracranial hemorrhage, with loss of consciousness of unspecified duration
C0159174|ICD9CM|AB|800.36|Cl skull vlt fx-coma NOS
C0159176|ICD9CM|HT|800.4|Closed fracture of vault of skull with intracranial injury of other and unspecified nature
C0159177|ICD9CM|PT|800.40|Closed fracture of vault of skull with intracranial injury of other and unspecified nature, unspecified state of consciousness
C0159177|ICD9CM|AB|800.40|Cl skl vlt fx/br inj NEC
C0159178|ICD9CM|PT|800.41|Closed fracture of vault of skull with intracranial injury of other and unspecified nature, with no loss of consciousness
C0159178|ICD9CM|AB|800.41|Cl skull vlt fx w/o coma
C0159179|ICD9CM|PT|800.42|Closed fracture of vault of skull with intracranial injury of other and unspecified nature, with brief [less than one hour] loss of consciousness
C0159179|ICD9CM|AB|800.42|Cl skull vlt fx-brf coma
C0159180|ICD9CM|PT|800.43|Closed fracture of vault of skull with intracranial injury of other and unspecified nature, with moderate [1-24 hours] loss of consciousness
C0159180|ICD9CM|AB|800.43|Cl skull vlt fx-mod coma
C0159181|ICD9CM|PT|800.44|Closed fracture of vault of skull with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159181|ICD9CM|AB|800.44|Cl skl vlt fx-proln coma
C0159182|ICD9CM|PT|800.45|Closed fracture of vault of skull with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159182|ICD9CM|AB|800.45|Cl skul vlt fx-deep coma
C0159183|ICD9CM|PT|800.46|Closed fracture of vault of skull with intracranial injury of other and unspecified nature, with loss of consciousness of unspecified duration
C0159183|ICD9CM|AB|800.46|Cl skull vlt fx-coma NOS
C0159184|ICD9CM|PT|800.49|Closed fracture of vault of skull with intracranial injury of other and unspecified nature, with concussion, unspecified
C0159184|ICD9CM|AB|800.49|Cl skl vlt fx-concus NOS
C0159185|ICD9CM|HT|800.5|Open fracture of vault of skull without mention of intracranial injury
C0159186|ICD9CM|PT|800.50|Open fracture of vault of skull without mention of intracranial injury, unspecified state of consciousness
C0159186|ICD9CM|AB|800.50|Opn skull vault fracture
C0159187|ICD9CM|PT|800.51|Open fracture of vault of skull without mention of intracranial injury, with no loss of consciousness
C0159187|ICD9CM|AB|800.51|Opn skul vlt fx w/o coma
C0159188|ICD9CM|PT|800.52|Open fracture of vault of skull without mention of intracranial injury, with brief [less than one hour] loss of consciousness
C0159188|ICD9CM|AB|800.52|Opn skul vlt fx-brf coma
C0159189|ICD9CM|PT|800.53|Open fracture of vault of skull without mention of intracranial injury, with moderate [1-24 hours] loss of consciousness
C0159189|ICD9CM|AB|800.53|Opn skul vlt fx-mod coma
C0159190|ICD9CM|PT|800.54|Open fracture of vault of skull without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159190|ICD9CM|AB|800.54|Opn skl vlt fx-proln com
C0159191|ICD9CM|PT|800.55|Open fracture of vault of skull without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159191|ICD9CM|AB|800.55|Opn skl vlt fx-deep coma
C0159192|ICD9CM|PT|800.56|Open fracture of vault of skull without mention of intracranial injury, with loss of consciousness of unspecified duration
C0159192|ICD9CM|AB|800.56|Opn skul vlt fx-coma NOS
C0159193|ICD9CM|PT|800.59|Open fracture of vault of skull without mention of intracranial injury, with concussion, unspecified
C0159193|ICD9CM|AB|800.59|Op skl vlt fx-concus NOS
C0159194|ICD9CM|HT|800.6|Open fracture of vault of skull with cerebral laceration and contusion
C0159195|ICD9CM|PT|800.60|Open fracture of vault of skull with cerebral laceration and contusion, unspecified state of consciousness
C0159195|ICD9CM|AB|800.60|Opn skl vlt fx/cereb lac
C0159196|ICD9CM|PT|800.61|Open fracture of vault of skull with cerebral laceration and contusion, with no loss of consciousness
C0159196|ICD9CM|AB|800.61|Opn skul vlt fx w/o coma
C0159197|ICD9CM|PT|800.62|Open fracture of vault of skull with cerebral laceration and contusion, with brief [less than one hour] loss of consciousness
C0159197|ICD9CM|AB|800.62|Opn skul vlt fx-brf coma
C0159198|ICD9CM|PT|800.63|Open fracture of vault of skull with cerebral laceration and contusion, with moderate [1-24 hours] loss of consciousness
C0159198|ICD9CM|AB|800.63|Opn skul vlt fx-mod coma
C0159199|ICD9CM|PT|800.64|Open fracture of vault of skull with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159199|ICD9CM|AB|800.64|Opn skl vlt fx-proln com
C0159200|ICD9CM|PT|800.65|Open fracture of vault of skull with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159200|ICD9CM|AB|800.65|Opn skl vlt fx-deep coma
C0159201|ICD9CM|PT|800.66|Open fracture of vault of skull with cerebral laceration and contusion, with loss of consciousness of unspecified duration
C0159201|ICD9CM|AB|800.66|Opn skul vlt fx-coma NOS
C0159203|ICD9CM|HT|800.7|Open fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage
C0159204|ICD9CM|PT|800.70|Open fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, unspecified state of consciousness
C0159204|ICD9CM|AB|800.70|Opn skl vlt fx/menin hem
C0159205|ICD9CM|PT|800.71|Open fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with no loss of consciousness
C0159205|ICD9CM|AB|800.71|Opn skul vlt fx w/o coma
C0159206|ICD9CM|PT|800.72|Open fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with brief [less than one hour] loss of consciousness
C0159206|ICD9CM|AB|800.72|Opn skul vlt fx-brf coma
C0159207|ICD9CM|PT|800.73|Open fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159207|ICD9CM|AB|800.73|Opn skul vlt fx-mod coma
C0159208|ICD9CM|PT|800.74|Open fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159208|ICD9CM|AB|800.74|Opn skl vlt fx-proln com
C0159209|ICD9CM|PT|800.75|Open fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159209|ICD9CM|AB|800.75|Opn skl vlt fx-deep coma
C0159210|ICD9CM|PT|800.76|Open fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with loss of consciousness of unspecified duration
C0159210|ICD9CM|AB|800.76|Opn skul vlt fx-coma NOS
C0159212|ICD9CM|HT|800.8|Open fracture of vault of skull with other and unspecified intracranial hemorrhage
C0159213|ICD9CM|PT|800.80|Open fracture of vault of skull with other and unspecified intracranial hemorrhage, unspecified state of consciousness
C0159213|ICD9CM|AB|800.80|Opn skull vlt fx/hem NEC
C0159214|ICD9CM|PT|800.81|Open fracture of vault of skull with other and unspecified intracranial hemorrhage, with no loss of consciousness
C0159214|ICD9CM|AB|800.81|Opn skul vlt fx w/o coma
C0159215|ICD9CM|PT|800.82|Open fracture of vault of skull with other and unspecified intracranial hemorrhage, with brief [less than one hour] loss of consciousness
C0159215|ICD9CM|AB|800.82|Opn skul vlt fx-brf coma
C0159216|ICD9CM|PT|800.83|Open fracture of vault of skull with other and unspecified intracranial hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159216|ICD9CM|AB|800.83|Opn skul vlt fx-mod coma
C0159217|ICD9CM|PT|800.84|Open fracture of vault of skull with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159217|ICD9CM|AB|800.84|Opn skl vlt fx-proln com
C0159218|ICD9CM|PT|800.85|Open fracture of vault of skull with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159218|ICD9CM|AB|800.85|Opn skl vlt fx-deep coma
C0159219|ICD9CM|PT|800.86|Open fracture of vault of skull with other and unspecified intracranial hemorrhage, with loss of consciousness of unspecified duration
C0159219|ICD9CM|AB|800.86|Opn skul vlt fx-coma NOS
C0159221|ICD9CM|HT|800.9|Open fracture of vault of skull with intracranial injury of other and unspecified nature
C0159222|ICD9CM|PT|800.90|Open fracture of vault of skull with intracranial injury of other and unspecified nature, unspecified state of consciousness
C0159222|ICD9CM|AB|800.90|Op skl vlt fx/br inj NEC
C0159223|ICD9CM|PT|800.91|Open fracture of vault of skull with intracranial injury of other and unspecified nature, with no loss of consciousness
C0159223|ICD9CM|AB|800.91|Opn skul vlt fx w/o coma
C0159224|ICD9CM|PT|800.92|Open fracture of vault of skull with intracranial injury of other and unspecified nature, with brief [less than one hour] loss of consciousness
C0159224|ICD9CM|AB|800.92|Opn skul vlt fx-brf coma
C0159225|ICD9CM|PT|800.93|Open fracture of vault of skull with intracranial injury of other and unspecified nature, with moderate [1-24 hours] loss of consciousness
C0159225|ICD9CM|AB|800.93|Opn skul vlt fx-mod coma
C0159226|ICD9CM|PT|800.94|Open fracture of vault of skull with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159226|ICD9CM|AB|800.94|Opn skl vlt fx-proln com
C0159227|ICD9CM|PT|800.95|Open fracture of vault of skull with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159227|ICD9CM|AB|800.95|Op skul vlt fx-deep coma
C0159228|ICD9CM|PT|800.96|Open fracture of vault of skull with intracranial injury of other and unspecified nature, with loss of consciousness of unspecified duration
C0159228|ICD9CM|AB|800.96|Opn skul vlt fx-coma NOS
C0159229|ICD9CM|PT|800.99|Open fracture of vault of skull with intracranial injury of other and unspecified nature, with concussion, unspecified
C0159229|ICD9CM|AB|800.99|Op skl vlt fx-concus NOS
C0159232|ICD9CM|PT|801.00|Closed fracture of base of skull without mention of intra cranial injury, unspecified state of consciousness
C0159232|ICD9CM|AB|801.00|Clos skull base fracture
C0159233|ICD9CM|PT|801.01|Closed fracture of base of skull without mention of intra cranial injury, with no loss of consciousness
C0159233|ICD9CM|AB|801.01|Cl skul base fx w/o coma
C0159234|ICD9CM|PT|801.02|Closed fracture of base of skull without mention of intra cranial injury, with brief [less than one hour] loss of consciousness
C0159234|ICD9CM|AB|801.02|Cl skul base fx-brf coma
C0159235|ICD9CM|PT|801.03|Closed fracture of base of skull without mention of intra cranial injury, with moderate [1-24 hours] loss of consciousness
C0159235|ICD9CM|AB|801.03|Cl skul base fx-mod coma
C0159236|ICD9CM|PT|801.04|Closed fracture of base of skull without mention of intra cranial injury, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159236|ICD9CM|AB|801.04|Cl skl base fx-prol coma
C0159237|ICD9CM|PT|801.05|Closed fracture of base of skull without mention of intra cranial injury, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159237|ICD9CM|AB|801.05|Cl skl base fx-deep coma
C0159238|ICD9CM|PT|801.06|Closed fracture of base of skull without mention of intra cranial injury, with loss of consciousness of unspecified duration
C0159238|ICD9CM|AB|801.06|Cl skul base fx-coma NOS
C0159239|ICD9CM|PT|801.09|Closed fracture of base of skull without mention of intra cranial injury, with concussion, unspecified
C0159239|ICD9CM|AB|801.09|Cl skull base fx-concuss
C0159240|ICD9CM|HT|801.1|Closed fracture of base of skull with cerebral laceration and contusion
C0159241|ICD9CM|PT|801.10|Closed fracture of base of skull with cerebral laceration and contusion, unspecified state of consciousness
C0159241|ICD9CM|AB|801.10|Cl skl base fx/cereb lac
C0159242|ICD9CM|PT|801.11|Closed fracture of base of skull with cerebral laceration and contusion, with no loss of consciousness
C0159242|ICD9CM|AB|801.11|Cl skul base fx w/o coma
C0159243|ICD9CM|PT|801.12|Closed fracture of base of skull with cerebral laceration and contusion, with brief [less than one hour] loss of consciousness
C0159243|ICD9CM|AB|801.12|Cl skul base fx-brf coma
C0159244|ICD9CM|PT|801.13|Closed fracture of base of skull with cerebral laceration and contusion, with moderate [1-24 hours] loss of consciousness
C0159244|ICD9CM|AB|801.13|Cl skul base fx-mod coma
C0159245|ICD9CM|PT|801.14|Closed fracture of base of skull with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159245|ICD9CM|AB|801.14|Cl skl base fx-prol coma
C0159246|ICD9CM|PT|801.15|Closed fracture of base of skull with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159246|ICD9CM|AB|801.15|Cl skl base fx-deep coma
C0159247|ICD9CM|PT|801.16|Closed fracture of base of skull with cerebral laceration and contusion, with loss of consciousness of unspecified duration
C0159247|ICD9CM|AB|801.16|Cl skul base fx-coma NOS
C0159249|ICD9CM|HT|801.2|Closed fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage
C0159250|ICD9CM|PT|801.20|Closed fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, unspecified state of consciousness
C0159250|ICD9CM|AB|801.20|Cl skl base fx/menin hem
C0159251|ICD9CM|PT|801.21|Closed fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with no loss of consciousness
C0159251|ICD9CM|AB|801.21|Cl skul base fx w/o coma
C0159252|ICD9CM|PT|801.22|Closed fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with brief [less than one hour] loss of consciousness
C0159252|ICD9CM|AB|801.22|Cl skul base fx/brf coma
C0159253|ICD9CM|PT|801.23|Closed fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159253|ICD9CM|AB|801.23|Cl skul base fx-mod coma
C0159254|ICD9CM|PT|801.24|Closed fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159254|ICD9CM|AB|801.24|Cl skl base fx-prol coma
C0159255|ICD9CM|PT|801.25|Closed fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159255|ICD9CM|AB|801.25|Cl skl base fx-deep coma
C0159256|ICD9CM|PT|801.26|Closed fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with loss of consciousness of unspecified duration
C0159256|ICD9CM|AB|801.26|Cl skul base fx-coma NOS
C0159258|ICD9CM|HT|801.3|Closed fracture of base of skull with other and unspecified intracranial hemorrhage
C0159259|ICD9CM|PT|801.30|Closed fracture of base of skull with other and unspecified intracranial hemorrhage, unspecified state of consciousness
C0159259|ICD9CM|AB|801.30|Cl skull base fx/hem NEC
C0159260|ICD9CM|PT|801.31|Closed fracture of base of skull with other and unspecified intracranial hemorrhage, with no loss of consciousness
C0159260|ICD9CM|AB|801.31|Cl skul base fx w/o coma
C0159261|ICD9CM|PT|801.32|Closed fracture of base of skull with other and unspecified intracranial hemorrhage, with brief [less than one hour] loss of consciousness
C0159261|ICD9CM|AB|801.32|Cl skul base fx-brf coma
C0159262|ICD9CM|PT|801.33|Closed fracture of base of skull with other and unspecified intracranial hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159262|ICD9CM|AB|801.33|Cl skul base fx-mod coma
C0159263|ICD9CM|PT|801.34|Closed fracture of base of skull with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159263|ICD9CM|AB|801.34|Cl skl base fx-prol coma
C0159264|ICD9CM|PT|801.35|Closed fracture of base of skull with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159264|ICD9CM|AB|801.35|Cl skl base fx-deep coma
C0159265|ICD9CM|PT|801.36|Closed fracture of base of skull with other and unspecified intracranial hemorrhage, with loss of consciousness of unspecified duration
C0159265|ICD9CM|AB|801.36|Cl skul base fx-coma NOS
C0159267|ICD9CM|HT|801.4|Closed fracture of base of skull with intracranial injury of other and unspecified nature
C0159268|ICD9CM|PT|801.40|Closed fracture of base of skull with intracranial injury of other and unspecified nature, unspecified state of consciousness
C0159268|ICD9CM|AB|801.40|Cl sk base fx/br inj NEC
C0159269|ICD9CM|PT|801.41|Closed fracture of base of skull with intracranial injury of other and unspecified nature, with no loss of consciousness
C0159269|ICD9CM|AB|801.41|Cl skul base fx w/o coma
C0159270|ICD9CM|PT|801.42|Closed fracture of base of skull with intracranial injury of other and unspecified nature, with brief [less than one hour] loss of consciousness
C0159270|ICD9CM|AB|801.42|Cl skul base fx-brf coma
C0159271|ICD9CM|PT|801.43|Closed fracture of base of skull with intracranial injury of other and unspecified nature, with moderate [1-24 hours] loss of consciousness
C0159271|ICD9CM|AB|801.43|Cl skul base fx-mod coma
C0159272|ICD9CM|PT|801.44|Closed fracture of base of skull with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours) loss of consciousness and return to pre-existing conscious level
C0159272|ICD9CM|AB|801.44|Cl skl base fx-prol coma
C0159273|ICD9CM|PT|801.45|Closed fracture of base of skull with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159273|ICD9CM|AB|801.45|Cl skl base fx-deep coma
C0159274|ICD9CM|PT|801.46|Closed fracture of base of skull with intracranial injury of other and unspecified nature, with loss of consciousness of unspecified duration
C0159274|ICD9CM|AB|801.46|Cl skul base fx-coma NOS
C0159275|ICD9CM|PT|801.49|Closed fracture of base of skull with intracranial injury of other and unspecified nature, with concussion, unspecified
C0159275|ICD9CM|AB|801.49|Cl skull base fx-concuss
C0159276|ICD9CM|HT|801.5|Open fracture of base of skull without mention of intracranial injury
C0159277|ICD9CM|PT|801.50|Open fracture of base of skull without mention of intracranial injury, unspecified state of consciousness
C0159277|ICD9CM|AB|801.50|Open skull base fracture
C0159278|ICD9CM|PT|801.51|Open fracture of base of skull without mention of intracranial injury, with no loss of consciousness
C0159278|ICD9CM|AB|801.51|Opn skl base fx w/o coma
C0159279|ICD9CM|PT|801.52|Open fracture of base of skull without mention of intracranial injury, with brief [less than one hour] loss of consciousness
C0159279|ICD9CM|AB|801.52|Opn skl base fx-brf coma
C0159280|ICD9CM|PT|801.53|Open fracture of base of skull without mention of intracranial injury, with moderate [1-24 hours] loss of consciousness
C0159280|ICD9CM|AB|801.53|Opn skl base fx-mod coma
C0159281|ICD9CM|PT|801.54|Open fracture of base of skull without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159281|ICD9CM|AB|801.54|Op skl base fx-prol coma
C0159282|ICD9CM|PT|801.55|Open fracture of base of skull without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159282|ICD9CM|AB|801.55|Op skl base fx-deep coma
C0159283|ICD9CM|PT|801.56|Open fracture of base of skull without mention of intracranial injury, with loss of consciousness of unspecified duration
C0159283|ICD9CM|AB|801.56|Opn skl base fx-coma NOS
C0159284|ICD9CM|PT|801.59|Open fracture of base of skull without mention of intracranial injury, with concussion, unspecified
C0159284|ICD9CM|AB|801.59|Opn skul base fx-concuss
C0159285|ICD9CM|HT|801.6|Open fracture of base of skull with cerebral laceration and contusion
C0159286|ICD9CM|PT|801.60|Open fracture of base of skull with cerebral laceration and contusion, unspecified state of consciousness
C0159286|ICD9CM|AB|801.60|Op skl base fx/cereb lac
C0159287|ICD9CM|PT|801.61|Open fracture of base of skull with cerebral laceration and contusion, with no loss of consciousness
C0159287|ICD9CM|AB|801.61|Opn skl base fx w/o coma
C0159288|ICD9CM|PT|801.62|Open fracture of base of skull with cerebral laceration and contusion, with brief [less than one hour] loss of consciousness
C0159288|ICD9CM|AB|801.62|Opn skl base fx-brf coma
C0159289|ICD9CM|PT|801.63|Open fracture of base of skull with cerebral laceration and contusion, with moderate [1-24 hours] loss of consciousness
C0159289|ICD9CM|AB|801.63|Opn skl base fx-mod coma
C0159290|ICD9CM|PT|801.64|Open fracture of base of skull with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159290|ICD9CM|AB|801.64|Op skl base fx-prol coma
C0159291|ICD9CM|PT|801.65|Open fracture of base of skull with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159291|ICD9CM|AB|801.65|Op skl base fx-deep coma
C0159292|ICD9CM|PT|801.66|Open fracture of base of skull with cerebral laceration and contusion, with loss of consciousness of unspecified duration
C0159292|ICD9CM|AB|801.66|Opn skl base fx-coma NOS
C0159294|ICD9CM|HT|801.7|Open fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage
C0159295|ICD9CM|PT|801.70|Open fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, unspecified state of consciousness
C0159295|ICD9CM|AB|801.70|Op skl base fx/menin hem
C0159296|ICD9CM|PT|801.71|Open fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with no loss of consciousness
C0159296|ICD9CM|AB|801.71|Opn skl base fx w/o coma
C0159297|ICD9CM|PT|801.72|Open fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with brief [less than one hour] loss of consciousness
C0159297|ICD9CM|AB|801.72|Opn skl base fx-brf coma
C0159298|ICD9CM|PT|801.73|Open fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159298|ICD9CM|AB|801.73|Opn skl base fx-mod coma
C0159299|ICD9CM|PT|801.74|Open fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159299|ICD9CM|AB|801.74|Op skl base fx-prol coma
C0159300|ICD9CM|PT|801.75|Open fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159300|ICD9CM|AB|801.75|Op skl base fx-deep coma
C0159301|ICD9CM|PT|801.76|Open fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with loss of consciousness of unspecified duration
C0159301|ICD9CM|AB|801.76|Opn skl base fx-coma NOS
C0159303|ICD9CM|HT|801.8|Open fracture of base of skull with other and unspecified intracranial hemorrhage
C0159304|ICD9CM|PT|801.80|Open fracture of base of skull with other and unspecified intracranial hemorrhage, unspecified state of consciousness
C0159304|ICD9CM|AB|801.80|Opn skul base fx/hem NEC
C0159305|ICD9CM|PT|801.81|Open fracture of base of skull with other and unspecified intracranial hemorrhage, with no loss of consciousness
C0159305|ICD9CM|AB|801.81|Opn skl base fx w/o coma
C0159306|ICD9CM|PT|801.82|Open fracture of base of skull with other and unspecified intracranial hemorrhage, with brief [less than one hour] loss of consciousness
C0159306|ICD9CM|AB|801.82|Opn skl base fx-brf coma
C0159307|ICD9CM|PT|801.83|Open fracture of base of skull with other and unspecified intracranial hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159307|ICD9CM|AB|801.83|Opn skl base fx-mod coma
C0159308|ICD9CM|PT|801.84|Open fracture of base of skull with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159308|ICD9CM|AB|801.84|Op skl base fx-prol coma
C0159309|ICD9CM|PT|801.85|Open fracture of base of skull with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159309|ICD9CM|AB|801.85|Op skl base fx-deep coma
C0159310|ICD9CM|PT|801.86|Open fracture of base of skull with other and unspecified intracranial hemorrhage, with loss of consciousness of unspecified duration
C0159310|ICD9CM|AB|801.86|Opn skl base fx-coma NOS
C0159312|ICD9CM|HT|801.9|Open fracture of base of skull with intracranial injury of other and unspecified nature
C0159313|ICD9CM|PT|801.90|Open fracture of base of skull with intracranial injury of other and unspecified nature, unspecified state of consciousness
C0159313|ICD9CM|AB|801.90|Op sk base fx/br inj NEC
C0159314|ICD9CM|PT|801.91|Open fracture of base of skull with intracranial injury of other and unspecified nature, with no loss of consciousness
C0159314|ICD9CM|AB|801.91|Op skul base fx w/o coma
C0159315|ICD9CM|PT|801.92|Open fracture of base of skull with intracranial injury of other and unspecified nature, with brief [less than one hour] loss of consciousness
C0159315|ICD9CM|AB|801.92|Opn skl base fx-brf coma
C0159316|ICD9CM|PT|801.93|Open fracture of base of skull with intracranial injury of other and unspecified nature, with moderate [1-24 hours] loss of consciousness
C0159316|ICD9CM|AB|801.93|Opn skl base fx-mod coma
C0159317|ICD9CM|PT|801.94|Open fracture of base of skull with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159317|ICD9CM|AB|801.94|Op skl base fx-prol coma
C0159318|ICD9CM|PT|801.95|Open fracture of base of skull with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159318|ICD9CM|AB|801.95|Op skl base fx-deep coma
C0159319|ICD9CM|PT|801.96|Open fracture of base of skull with intracranial injury of other and unspecified nature, with loss of consciousness of unspecified duration
C0159319|ICD9CM|AB|801.96|Opn skl base fx-coma NOS
C0159320|ICD9CM|PT|801.99|Open fracture of base of skull with intracranial injury of other and unspecified nature, with concussion, unspecified
C0159320|ICD9CM|AB|801.99|Opn skul base fx-concuss
C0159321|ICD9CM|HT|802|Fracture of face bones
C0159322|ICD9CM|PT|802.0|Closed fracture of nasal bones
C0159322|ICD9CM|AB|802.0|Nasal bone fx-closed
C0159323|ICD9CM|PT|802.1|Open fracture of nasal bones
C0159323|ICD9CM|AB|802.1|Nasal bone fx-open
C0159324|ICD9CM|HT|802.2|Mandible closed fracture
C0159324|ICD9CM|PT|802.20|Closed fracture of mandible, unspecified site
C0159324|ICD9CM|AB|802.20|Mandible fx NOS-closed
C0159325|ICD9CM|PT|802.21|Closed fracture of mandible, condylar process
C0159325|ICD9CM|AB|802.21|Fx condyl proc mandib-cl
C0159327|ICD9CM|PT|802.23|Closed fracture of mandible, coronoid process
C0159327|ICD9CM|AB|802.23|Fx coron proc mandib-cl
C0159330|ICD9CM|PT|802.26|Closed fracture of mandible, symphysis of body
C0159330|ICD9CM|AB|802.26|Fx symphy mandib body-cl
C0159331|ICD9CM|PT|802.27|Closed fracture of mandible, alveolar border of body
C0159331|ICD9CM|AB|802.27|Fx alveolar bord mand-cl
C0159333|ICD9CM|PT|802.29|Closed fracture of mandible, multiple sites
C0159333|ICD9CM|AB|802.29|Mult fx mandible-closed
C0159334|ICD9CM|HT|802.3|Mandible open fracture
C0159334|ICD9CM|PT|802.30|Open fracture of mandible, unspecified site
C0159334|ICD9CM|AB|802.30|Mandible fx NOS-open
C0159336|ICD9CM|PT|802.31|Open fracture of mandible, condylar process
C0159336|ICD9CM|AB|802.31|Fx condyl proc mand-open
C0159338|ICD9CM|PT|802.33|Open fracture of mandible, coronoid process
C0159338|ICD9CM|AB|802.33|Fx coron proc mandib-opn
C0159341|ICD9CM|PT|802.36|Open fracture of mandible, symphysis of body
C0159341|ICD9CM|AB|802.36|Fx symphy mandib bdy-opn
C0159342|ICD9CM|PT|802.37|Open fracture of mandible, alveolar border of body
C0159342|ICD9CM|AB|802.37|Fx alv bord mand bdy-opn
C0159344|ICD9CM|PT|802.39|Open fracture of mandible, multiple sites
C0159344|ICD9CM|AB|802.39|Mult fx mandible-open
C0159345|ICD9CM|PT|802.5|Open fracture of malar and maxillary bones
C0159345|ICD9CM|AB|802.5|Fx malar/maxillary-open
C0159348|ICD9CM|PT|802.8|Closed fracture of other facial bones
C0159348|ICD9CM|AB|802.8|Fx facial bone NEC-close
C0159349|ICD9CM|PT|802.9|Open fracture of other facial bones
C0159349|ICD9CM|AB|802.9|Fx facial bone NEC-open
C0159350|ICD9CM|HT|803|Other and unqualified skull fractures
C0159351|ICD9CM|PT|803.00|Other closed skull fracture without mention of intracranial injury, unspecified state of consciousness
C0159351|ICD9CM|AB|803.00|Close skull fracture NEC
C0159352|ICD9CM|PT|803.01|Other closed skull fracture without mention of intracranial injury, with no loss of consciousness
C0159352|ICD9CM|AB|803.01|Cl skull fx NEC w/o coma
C0159353|ICD9CM|PT|803.02|Other closed skull fracture without mention of intracranial injury, with brief [less than one hour] loss of consciousness
C0159353|ICD9CM|AB|803.02|Cl skull fx NEC-brf coma
C0159354|ICD9CM|PT|803.03|Other closed skull fracture without mention of intracranial injury, with moderate [1-24 hours] loss of consciousness
C0159354|ICD9CM|AB|803.03|Cl skull fx NEC-mod coma
C0159355|ICD9CM|PT|803.04|Other closed skull fracture without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159355|ICD9CM|AB|803.04|Cl skl fx NEC-proln coma
C0159356|ICD9CM|PT|803.05|Other closed skull fracture without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159356|ICD9CM|AB|803.05|Cl skul fx NEC-deep coma
C0159357|ICD9CM|PT|803.06|Other closed skull fracture without mention of intracranial injury, with loss of consciousness of unspecified duration
C0159357|ICD9CM|AB|803.06|Cl skull fx NEC-coma NOS
C0159358|ICD9CM|PT|803.09|Other closed skull fracture without mention of intracranial injury, with concussion, unspecified
C0159358|ICD9CM|AB|803.09|Cl skull fx NEC-concuss
C0159359|ICD9CM|HT|803.1|Other closed skull fracture with cerebral laceration and contusion
C0159360|ICD9CM|PT|803.10|Other closed skull fracture with cerebral laceration and contusion, unspecified state of consciousness
C0159360|ICD9CM|AB|803.10|Cl skl fx NEC/cerebr lac
C0159361|ICD9CM|PT|803.11|Other closed skull fracture with cerebral laceration and contusion, with no loss of consciousness
C0159361|ICD9CM|AB|803.11|Cl skull fx NEC w/o coma
C0159362|ICD9CM|PT|803.12|Other closed skull fracture with cerebral laceration and contusion, with brief [less than one hour] loss of consciousness
C0159362|ICD9CM|AB|803.12|Cl skull fx NEC-brf coma
C0159363|ICD9CM|PT|803.13|Other closed skull fracture with cerebral laceration and contusion, with moderate [1-24 hours] loss of consciousness
C0159363|ICD9CM|AB|803.13|Cl skull fx NEC-mod coma
C0159364|ICD9CM|PT|803.14|Other closed skull fracture with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159364|ICD9CM|AB|803.14|Cl skl fx NEC-proln coma
C0159365|ICD9CM|PT|803.15|Other closed skull fracture with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159365|ICD9CM|AB|803.15|Cl skul fx NEC-deep coma
C0159366|ICD9CM|PT|803.16|Other closed skull fracture with cerebral laceration and contusion, with loss of consciousness of unspecified duration
C0159366|ICD9CM|AB|803.16|Cl skull fx NEC-coma NOS
C0159368|ICD9CM|HT|803.2|Other closed skull fracture with subarachnoid, subdural, and extradural hemorrhage
C0159369|ICD9CM|PT|803.20|Other closed skull fracture with subarachnoid, subdural, and extradural hemorrhage, unspecified state of consciousness
C0159369|ICD9CM|AB|803.20|Cl skl fx NEC/mening hem
C0159370|ICD9CM|PT|803.21|Other closed skull fracture with subarachnoid, subdural, and extradural hemorrhage, with no loss of consciousness
C0159370|ICD9CM|AB|803.21|Cl skull fx NEC w/o coma
C0159371|ICD9CM|PT|803.22|Other closed skull fracture with subarachnoid, subdural, and extradural hemorrhage, with brief [less than one hour] loss of consciousness
C0159371|ICD9CM|AB|803.22|Cl skull fx NEC-brf coma
C0159372|ICD9CM|PT|803.23|Other closed skull fracture with subarachnoid, subdural, and extradural hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159372|ICD9CM|AB|803.23|Cl skull fx NEC-mod coma
C0159373|ICD9CM|PT|803.24|Other closed skull fracture with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159373|ICD9CM|AB|803.24|Cl skl fx NEC-proln coma
C0159374|ICD9CM|PT|803.25|Other closed skull fracture with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159374|ICD9CM|AB|803.25|Cl skul fx NEC-deep coma
C0159375|ICD9CM|PT|803.26|Other closed skull fracture with subarachnoid, subdural, and extradural hemorrhage, with loss of consciousness of unspecified duration
C0159375|ICD9CM|AB|803.26|Cl skull fx NEC-coma NOS
C0159377|ICD9CM|HT|803.3|Closed skull fracture with other and unspecified intracranial hemorrhage
C0159378|ICD9CM|PT|803.30|Other closed skull fracture with other and unspecified intracranial hemorrhage, unspecified state of unconsciousness
C0159378|ICD9CM|AB|803.30|Cl skull fx NEC/hem NEC
C0159379|ICD9CM|PT|803.31|Other closed skull fracture with other and unspecified intracranial hemorrhage, with no loss of consciousness
C0159379|ICD9CM|AB|803.31|Cl skull fx NEC w/o coma
C0159380|ICD9CM|PT|803.32|Other closed skull fracture with other and unspecified intracranial hemorrhage, with brief [less than one hour] loss of consciousness
C0159380|ICD9CM|AB|803.32|Cl skull fx NEC-brf coma
C0159381|ICD9CM|PT|803.33|Other closed skull fracture with other and unspecified intracranial hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159381|ICD9CM|AB|803.33|Cl skull fx NEC-mod coma
C0159382|ICD9CM|PT|803.34|Other closed skull fracture with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159382|ICD9CM|AB|803.34|Cl skl fx NEC-proln coma
C0159383|ICD9CM|PT|803.35|Other closed skull fracture with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159383|ICD9CM|AB|803.35|Cl skul fx NEC-deep coma
C0159384|ICD9CM|PT|803.36|Other closed skull fracture with other and unspecified intracranial hemorrhage, with loss of consciousness of unspecified duration
C0159384|ICD9CM|AB|803.36|Cl skull fx NEC-coma NOS
C0159386|ICD9CM|HT|803.4|Other closed skull fracture with intracranial injury of other and unspecified nature
C0159387|ICD9CM|PT|803.40|Other closed skull fracture with intracranial injury of other and unspecified nature, unspecified state of consciousness
C0159387|ICD9CM|AB|803.40|Cl skl fx NEC/br inj NEC
C0159388|ICD9CM|PT|803.41|Other closed skull fracture with intracranial injury of other and unspecified nature, with no loss of consciousness
C0159388|ICD9CM|AB|803.41|Cl skull fx NEC w/o coma
C0159389|ICD9CM|PT|803.42|Other closed skull fracture with intracranial injury of other and unspecified nature, with brief [less than one hour] loss of consciousness
C0159389|ICD9CM|AB|803.42|Cl skull fx NEC-brf coma
C0159390|ICD9CM|PT|803.43|Other closed skull fracture with intracranial injury of other and unspecified nature, with moderate [1-24 hours] loss of consciousness
C0159390|ICD9CM|AB|803.43|Cl skull fx NEC-mod coma
C0159391|ICD9CM|PT|803.44|Other closed skull fracture with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159391|ICD9CM|AB|803.44|Cl skl fx NEC-proln coma
C0159392|ICD9CM|PT|803.45|Other closed skull fracture with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159392|ICD9CM|AB|803.45|Cl skul fx NEC-deep coma
C0159393|ICD9CM|PT|803.46|Other closed skull fracture with intracranial injury of other and unspecified nature, with loss of consciousness of unspecified duration
C0159393|ICD9CM|AB|803.46|Cl skull fx NEC-coma NOS
C0159394|ICD9CM|PT|803.49|Other closed skull fracture with intracranial injury of other and unspecified nature, with concussion, unspecified
C0159394|ICD9CM|AB|803.49|Cl skull fx NEC-concuss
C0159395|ICD9CM|HT|803.5|Other open skull fracture without mention of intracranial injury
C0159396|ICD9CM|PT|803.50|Other open skull fracture without mention of injury, unspecified state of consciousness
C0159396|ICD9CM|AB|803.50|Open skull fracture NEC
C0159397|ICD9CM|PT|803.51|Other open skull fracture without mention of intracranial injury, with no loss of consciousness
C0159397|ICD9CM|AB|803.51|Opn skul fx NEC w/o coma
C0159398|ICD9CM|PT|803.52|Other open skull fracture without mention of intracranial injury, with brief [less than one hour] loss of consciousness
C0159398|ICD9CM|AB|803.52|Opn skul fx NEC-brf coma
C0159399|ICD9CM|PT|803.53|Other open skull fracture without mention of intracranial injury, with moderate [1-24 hours] loss of consciousness
C0159399|ICD9CM|AB|803.53|Opn skul fx NEC-mod coma
C0159400|ICD9CM|PT|803.54|Other open skull fracture without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159400|ICD9CM|AB|803.54|Opn skl fx NEC-prol coma
C0159401|ICD9CM|PT|803.55|Other open skull fracture without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159401|ICD9CM|AB|803.55|Opn skl fx NEC-deep coma
C0159402|ICD9CM|PT|803.56|Other open skull fracture without mention of intracranial injury, with loss of consciousness of unspecified duration
C0159402|ICD9CM|AB|803.56|Opn skul fx NEC-coma NOS
C0159403|ICD9CM|PT|803.59|Other open skull fracture without mention of intracranial injury, with concussion, unspecified
C0159403|ICD9CM|AB|803.59|Opn skull fx NEC-concuss
C0159404|ICD9CM|HT|803.6|Other open skull fracture with cerebral laceration and contusion
C0159405|ICD9CM|PT|803.60|Other open skull fracture with cerebral laceration and contusion, unspecified state of consciousness
C0159405|ICD9CM|AB|803.60|Opn skl fx NEC/cereb lac
C0159406|ICD9CM|PT|803.61|Other open skull fracture with cerebral laceration and contusion, with no loss of consciousness
C0159406|ICD9CM|AB|803.61|Opn skul fx NEC w/o coma
C0159407|ICD9CM|PT|803.62|Other open skull fracture with cerebral laceration and contusion, with brief [less than one hour] loss of consciousness
C0159407|ICD9CM|AB|803.62|Opn skul fx NEC-brf coma
C0159408|ICD9CM|PT|803.63|Other open skull fracture with cerebral laceration and contusion, with moderate [1-24 hours] loss of consciousness
C0159408|ICD9CM|AB|803.63|Opn skul fx NEC-mod coma
C0159409|ICD9CM|PT|803.64|Other open skull fracture with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159409|ICD9CM|AB|803.64|Opn skl fx NEC-proln com
C0159410|ICD9CM|PT|803.65|Other open skull fracture with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159410|ICD9CM|AB|803.65|Opn skl fx NEC-deep coma
C0159411|ICD9CM|PT|803.66|Other open skull fracture with cerebral laceration and contusion, with loss of consciousness of unspecified duration
C0159411|ICD9CM|AB|803.66|Opn skul fx NEC-coma NOS
C0159413|ICD9CM|HT|803.7|Other open skull fracture with subarachnoid, subdural, and extradural hemorrhage
C0159414|ICD9CM|PT|803.70|Other open skull fracture with subarachnoid, subdural, and extradural hemorrhage, unspecified state of consciousness
C0159414|ICD9CM|AB|803.70|Opn skl fx NEC/menin hem
C0159415|ICD9CM|PT|803.71|Other open skull fracture with subarachnoid, subdural, and extradural hemorrhage, with no loss of consciousness
C0159415|ICD9CM|AB|803.71|Opn skul fx NEC w/o coma
C0159416|ICD9CM|PT|803.72|Other open skull fracture with subarachnoid, subdural, and extradural hemorrhage, with brief [less than one hour] loss of consciousness
C0159416|ICD9CM|AB|803.72|Opn skul fx NEC-brf coma
C0159417|ICD9CM|PT|803.73|Other open skull fracture with subarachnoid, subdural, and extradural hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159417|ICD9CM|AB|803.73|Opn skul fx NEC-mod coma
C0159418|ICD9CM|PT|803.74|Other open skull fracture with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159418|ICD9CM|AB|803.74|Opn skl fx NEC-prol coma
C0159419|ICD9CM|PT|803.75|Other open skull fracture with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159419|ICD9CM|AB|803.75|Opn skl fx NEC-deep coma
C0159420|ICD9CM|PT|803.76|Other open skull fracture with subarachnoid, subdural, and extradural hemorrhage, with loss of consciousness of unspecified duration
C0159420|ICD9CM|AB|803.76|Opn skul fx NEC-coma NOS
C0159422|ICD9CM|HT|803.8|Other open skull fracture with other and unspecified intracranial hemorrhage
C0159423|ICD9CM|PT|803.80|Other open skull fracture with other and unspecified intracranial hemorrhage, unspecified state of consciousness
C0159423|ICD9CM|AB|803.80|Opn skull fx NEC/hem NEC
C0159424|ICD9CM|PT|803.81|Other open skull fracture with other and unspecified intracranial hemorrhage, with no loss of consciousness
C0159424|ICD9CM|AB|803.81|Opn skul fx NEC w/o coma
C0159425|ICD9CM|PT|803.82|Other open skull fracture with other and unspecified intracranial hemorrhage, with brief [less than one hour] loss of consciousness
C0159425|ICD9CM|AB|803.82|Opn skul fx NEC-brf coma
C0159426|ICD9CM|PT|803.83|Other open skull fracture with other and unspecified intracranial hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159426|ICD9CM|AB|803.83|Opn skul fx NEC-mod coma
C0159427|ICD9CM|PT|803.84|Other open skull fracture with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159427|ICD9CM|AB|803.84|Opn skl fx NEC-prol coma
C0159428|ICD9CM|PT|803.85|Other open skull fracture with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159428|ICD9CM|AB|803.85|Opn skl fx NEC-deep coma
C0159429|ICD9CM|PT|803.86|Other open skull fracture with other and unspecified intracranial hemorrhage, with loss of consciousness of unspecified duration
C0159429|ICD9CM|AB|803.86|Opn skul fx NEC-coma NOS
C0159431|ICD9CM|HT|803.9|Other open skull fracture with intracranial injury of other and unspecified nature
C0159432|ICD9CM|PT|803.90|Other open skull fracture with intracranial injury of other and unspecified nature, unspecified state of consciousness
C0159432|ICD9CM|AB|803.90|Op skl fx NEC/br inj NEC
C0159433|ICD9CM|PT|803.91|Other open skull fracture with intracranial injury of other and unspecified nature, with no loss of consciousness
C0159433|ICD9CM|AB|803.91|Opn skul fx NEC w/o coma
C0159434|ICD9CM|PT|803.92|Other open skull fracture with intracranial injury of other and unspecified nature, with brief [less than one hour] loss of consciousness
C0159434|ICD9CM|AB|803.92|Opn skul fx NEC-brf coma
C0159435|ICD9CM|PT|803.93|Other open skull fracture with intracranial injury of other and unspecified nature, with moderate [1-24 hours] loss of consciousness
C0159435|ICD9CM|AB|803.93|Opn skul fx NEC-mod coma
C0159436|ICD9CM|PT|803.94|Other open skull fracture with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159436|ICD9CM|AB|803.94|Opn skl fx NEC-prol coma
C0159437|ICD9CM|PT|803.95|Other open skull fracture with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159437|ICD9CM|AB|803.95|Opn skl fx NEC-deep coma
C0159438|ICD9CM|PT|803.96|Other open skull fracture with intracranial injury of other and unspecified nature, with loss of consciousness of unspecified duration
C0159438|ICD9CM|AB|803.96|Opn skul fx NEC-coma NOS
C0159439|ICD9CM|PT|803.99|Other open skull fracture with intracranial injury of other and unspecified nature, with concussion, unspecified
C0159439|ICD9CM|AB|803.99|Opn skull fx NEC-concuss
C0159440|ICD9CM|HT|804|Multiple fractures involving skull or face with other bones
C0159441|ICD9CM|HT|804.0|Closed fractures involving skull or face with other bones, without mention of intracranial injury
C0159442|ICD9CM|PT|804.00|Closed fractures involving skull or face with other bones, without mention of intracranial injury, unspecified state of consciousness
C0159442|ICD9CM|AB|804.00|Cl skul fx w oth bone fx
C0159443|ICD9CM|PT|804.01|Closed fractures involving skull or face with other bones, without mention of intracranial injury, with no loss of consciousness
C0159443|ICD9CM|AB|804.01|Cl skl w oth fx w/o coma
C0159444|ICD9CM|PT|804.02|Closed fractures involving skull or face with other bones, without mention of intracranial injury, with brief [less than one hour] loss of consciousness
C0159444|ICD9CM|AB|804.02|Cl skl w oth fx-brf coma
C0159445|ICD9CM|PT|804.03|Closed fractures involving skull or face with other bones, without mention of intracranial injury, with moderate [1-24 hours] loss of consciousness
C0159445|ICD9CM|AB|804.03|Cl skl w oth fx-mod coma
C0159446|ICD9CM|PT|804.04|Closed fractures involving skull or face with other bones, without mention or intracranial injury, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159446|ICD9CM|AB|804.04|Cl skl/oth fx-proln coma
C0159447|ICD9CM|PT|804.05|Closed fractures involving skull of face with other bones, without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159447|ICD9CM|AB|804.05|Cl skul/oth fx-deep coma
C0159448|ICD9CM|PT|804.06|Closed fractures involving skull of face with other bones, without mention of intracranial injury, with loss of consciousness of unspecified duration
C0159448|ICD9CM|AB|804.06|Cl skl w oth fx-coma NOS
C0159449|ICD9CM|PT|804.09|Closed fractures involving skull of face with other bones, without mention of intracranial injury, with concussion, unspecified
C0159449|ICD9CM|AB|804.09|Cl skul w oth fx-concuss
C0159450|ICD9CM|HT|804.1|Closed fractures involving skull or face with other bones, with cerebral laceration and contusion
C0159451|ICD9CM|PT|804.10|Closed fractures involving skull or face with other bones, with cerebral laceration and contusion, unspecified state of consciousness
C0159451|ICD9CM|AB|804.10|Cl sk w oth fx/cereb lac
C0159452|ICD9CM|PT|804.11|Closed fractures involving skull or face with other bones, with cerebral laceration and contusion, with no loss of consciousness
C0159452|ICD9CM|AB|804.11|Cl skl w oth fx w/o coma
C0159453|ICD9CM|PT|804.12|Closed fractures involving skull or face with other bones, with cerebral laceration and contusion, with brief [less than one hour] loss of consciousness
C0159453|ICD9CM|AB|804.12|Cl skl w oth fx-brf coma
C0159454|ICD9CM|PT|804.13|Closed fractures involving skull or face with other bones, with cerebral laceration and contusion, with moderate [1-24 hours] loss of consciousness
C0159454|ICD9CM|AB|804.13|Cl skl w oth fx-mod coma
C0159455|ICD9CM|PT|804.14|Closed fractures involving skull or face with other bones, with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159455|ICD9CM|AB|804.14|Cl skl/oth fx-proln coma
C0159456|ICD9CM|PT|804.15|Closed fractures involving skull or face with other bones, with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159456|ICD9CM|AB|804.15|Cl skul/oth fx-deep coma
C0159457|ICD9CM|PT|804.16|Closed fractures involving skull or face with other bones, with cerebral laceration and contusion, with loss of consciousness of unspecified duration
C0159457|ICD9CM|AB|804.16|Cl skl w oth fx-coma NOS
C0159459|ICD9CM|HT|804.2|Closed fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage
C0159460|ICD9CM|PT|804.20|Closed fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, unspecified state of consciousness
C0159460|ICD9CM|AB|804.20|Cl skl/oth fx/mening hem
C0159461|ICD9CM|PT|804.21|Closed fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with no loss of consciousness
C0159461|ICD9CM|AB|804.21|Cl skl w oth fx w/o coma
C0159462|ICD9CM|PT|804.22|Closed fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with brief [less than one hour] loss of consciousness
C0159462|ICD9CM|AB|804.22|Cl skl w oth fx-brf coma
C0159463|ICD9CM|PT|804.23|Closed fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159463|ICD9CM|AB|804.23|Cl skl w oth fx-mod coma
C0159464|ICD9CM|PT|804.24|Closed fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159464|ICD9CM|AB|804.24|Cl skl/oth fx-proln coma
C0159465|ICD9CM|PT|804.25|Closed fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159465|ICD9CM|AB|804.25|Cl skul/oth fx-deep coma
C0159466|ICD9CM|PT|804.26|Closed fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with loss of consciousness of unspecified duration
C0159466|ICD9CM|AB|804.26|Cl skl w oth fx-coma NOS
C0159468|ICD9CM|HT|804.3|Closed fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage
C0159469|ICD9CM|PT|804.30|Closed fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, unspecified state of consciousness
C0159469|ICD9CM|AB|804.30|Cl skul w oth fx/hem NEC
C0159470|ICD9CM|PT|804.31|Closed fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with no loss of consciousness
C0159470|ICD9CM|AB|804.31|Cl skl w oth fx w/o coma
C0159471|ICD9CM|PT|804.32|Closed fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with brief [less than one hour] loss of consciousness
C0159471|ICD9CM|AB|804.32|Cl skl w oth fx-brf coma
C0159472|ICD9CM|PT|804.33|Closed fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159472|ICD9CM|AB|804.33|Cl skl w oth fx-mod coma
C0159473|ICD9CM|PT|804.34|Closed fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre- existing conscious level
C0159473|ICD9CM|AB|804.34|Cl skl/oth fx-proln coma
C0159474|ICD9CM|PT|804.35|Closed fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159474|ICD9CM|AB|804.35|Cl skul/oth fx-deep coma
C0159475|ICD9CM|PT|804.36|Closed fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with loss of consciousness of unspecified duration
C0159475|ICD9CM|AB|804.36|Cl skl w oth fx-coma NOS
C0159477|ICD9CM|HT|804.4|Closed fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature
C0159478|ICD9CM|PT|804.40|Closed fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, unspecified state of consciousness
C0159478|ICD9CM|AB|804.40|Cl skl/oth fx/br inj NEC
C0159479|ICD9CM|PT|804.41|Closed fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with no loss of consciousness
C0159479|ICD9CM|AB|804.41|Cl skl w oth fx w/o coma
C0159480|ICD9CM|PT|804.42|Closed fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with brief [less than one hour] loss of consciousness
C0159480|ICD9CM|AB|804.42|Cl skl w oth fx-brf coma
C0159481|ICD9CM|PT|804.43|Closed fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with moderate [1-24 hours] loss of consciousness
C0159481|ICD9CM|AB|804.43|Cl skl w oth fx-mod coma
C0159482|ICD9CM|PT|804.44|Closed fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159482|ICD9CM|AB|804.44|Cl skl/oth fx-proln coma
C0159483|ICD9CM|PT|804.45|Closed fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159483|ICD9CM|AB|804.45|Cl skul/oth fx-deep coma
C0159484|ICD9CM|PT|804.46|Closed fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with loss of consciousness of unspecified duration
C0159484|ICD9CM|AB|804.46|Cl skl w oth fx-coma NOS
C0159485|ICD9CM|PT|804.49|Closed fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with concussion, unspecified
C0159485|ICD9CM|AB|804.49|Cl skul w oth fx-concuss
C0159486|ICD9CM|HT|804.5|Open fractures involving skull or face with other bones, without mention of intracranial injury
C0159487|ICD9CM|PT|804.50|Open fractures involving skull or face with other bones, without mention of intracranial injury, unspecified state of consciousness
C0159487|ICD9CM|AB|804.50|Opn skull fx/oth bone fx
C0159488|ICD9CM|PT|804.51|Open fractures involving skull or face with other bones, without mention of intracranial injury, with no loss of consciousness
C0159488|ICD9CM|AB|804.51|Opn skul/oth fx w/o coma
C0159489|ICD9CM|PT|804.52|Open fractures involving skull or face with other bones, without mention of intracranial injury, with brief [less than one hour] loss of consciousness
C0159489|ICD9CM|AB|804.52|Opn skul/oth fx-brf coma
C0159490|ICD9CM|PT|804.53|Open fractures involving skull or face with other bones, without mention of intracranial injury, with moderate [1-24 hours] loss of consciousness
C0159490|ICD9CM|AB|804.53|Opn skul/oth fx-mod coma
C0159491|ICD9CM|PT|804.54|Open fractures involving skull or face with other bones, without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159491|ICD9CM|AB|804.54|Opn skl/oth fx-prol coma
C0159492|ICD9CM|PT|804.55|Open fractures involving skull or face with other bones, without mention of intracranial injury, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159492|ICD9CM|AB|804.55|Opn skl/oth fx-deep coma
C0159493|ICD9CM|PT|804.56|Open fractures involving skull or face with other bones, without mention of intracranial injury, with loss of consciousness of unspecified duration
C0159493|ICD9CM|AB|804.56|Opn skul/oth fx-coma NOS
C0159494|ICD9CM|PT|804.59|Open fractures involving skull or face with other bones, without mention of intracranial injury, with concussion, unspecified
C0159494|ICD9CM|AB|804.59|Opn skull/oth fx-concuss
C0159495|ICD9CM|HT|804.6|Open fractures involving skull or face with other bones, with cerebral laceration and contusion
C0159496|ICD9CM|PT|804.60|Open fractures involving skull or face with other bones, with cerebral laceration and contusion, unspecified state of consciousness
C0159496|ICD9CM|AB|804.60|Opn skl/oth fx/cereb lac
C0159497|ICD9CM|PT|804.61|Open fractures involving skull or face with other bones, with cerebral laceration and contusion, with no loss of consciousness
C0159497|ICD9CM|AB|804.61|Opn skul/oth fx w/o coma
C0159498|ICD9CM|PT|804.62|Open fractures involving skull or face with other bones, with cerebral laceration and contusion, with brief [less than one hour] loss of consciousness
C0159498|ICD9CM|AB|804.62|Opn skul/oth fx-brf coma
C0159499|ICD9CM|PT|804.63|Open fractures involving skull or face with other bones, with cerebral laceration and contusion, with moderate [1-24 hours] loss of consciousness
C0159499|ICD9CM|AB|804.63|Opn skul/oth fx-mod coma
C0159500|ICD9CM|PT|804.64|Open fractures involving skull or face with other bones, with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159500|ICD9CM|AB|804.64|Opn skl/oth fx-prol coma
C0159501|ICD9CM|PT|804.65|Open fractures involving skull or face with other bones, with cerebral laceration and contusion, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159501|ICD9CM|AB|804.65|Opn skl/oth fx-deep coma
C0159502|ICD9CM|PT|804.66|Open fractures involving skull or face with other bones, with cerebral laceration and contusion, with loss of consciousness of unspecified duration
C0159502|ICD9CM|AB|804.66|Opn skul/oth fx-coma NOS
C0159504|ICD9CM|HT|804.7|Open fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage
C0159505|ICD9CM|PT|804.70|Open fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, unspecified state of consciousness
C0159505|ICD9CM|AB|804.70|Opn skl/oth fx/menin hem
C0159506|ICD9CM|PT|804.71|Open fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with no loss of consciousness
C0159506|ICD9CM|AB|804.71|Opn skul/oth fx w/o coma
C0159507|ICD9CM|PT|804.72|Open fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with brief [less than one hour] loss of consciousness
C0159507|ICD9CM|AB|804.72|Opn skul/oth fx-brf coma
C0159508|ICD9CM|PT|804.73|Open fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159508|ICD9CM|AB|804.73|Opn skul/oth fx-mod coma
C0159509|ICD9CM|PT|804.74|Open fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159509|ICD9CM|AB|804.74|Opn skl/oth fx-prol coma
C0159510|ICD9CM|PT|804.75|Open fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with prolonged [more than 24 hours] loss of consciousness, without return to pre-existing conscious level
C0159510|ICD9CM|AB|804.75|Opn skl/oth fx-deep coma
C0159511|ICD9CM|PT|804.76|Open fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with loss of consciousness of unspecified duration
C0159511|ICD9CM|AB|804.76|Opn skul/oth fx-coma NOS
C0159513|ICD9CM|HT|804.8|Open fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage
C0159514|ICD9CM|PT|804.80|Open fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, unspecified state of consciousness
C0159514|ICD9CM|AB|804.80|Opn skl w oth fx/hem NEC
C0159515|ICD9CM|PT|804.81|Open fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with no loss of consciousness
C0159515|ICD9CM|AB|804.81|Opn skul/oth fx w/o coma
C0159516|ICD9CM|PT|804.82|Open fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with brief [less than one hour] loss of consciousness
C0159516|ICD9CM|AB|804.82|Opn skul/oth fx-brf coma
C0159517|ICD9CM|PT|804.83|Open fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with moderate [1-24 hours] loss of consciousness
C0159517|ICD9CM|AB|804.83|Opn skul/oth fx-mod coma
C0159518|ICD9CM|PT|804.84|Open fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159518|ICD9CM|AB|804.84|Opn skl/oth fx-prol coma
C0159519|ICD9CM|PT|804.85|Open fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with prolonged [more than 24 hours] loss consciousness, without return to pre-existing conscious level
C0159519|ICD9CM|AB|804.85|Opn skl/oth fx-deep coma
C0159520|ICD9CM|PT|804.86|Open fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with loss of consciousness of unspecified duration
C0159520|ICD9CM|AB|804.86|Opn skul/oth fx-coma NOS
C0159522|ICD9CM|HT|804.9|Open fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature
C0159523|ICD9CM|PT|804.90|Open fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, unspecified state of consciousness
C0159523|ICD9CM|AB|804.90|Op skl/oth fx/br inj NEC
C0159524|ICD9CM|PT|804.91|Open fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with no loss of consciousness
C0159524|ICD9CM|AB|804.91|Opn skul/oth fx w/o coma
C0159525|ICD9CM|PT|804.92|Open fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with brief [less than one hour] loss of consciousness
C0159525|ICD9CM|AB|804.92|Opn skul/oth fx-brf coma
C0159526|ICD9CM|PT|804.93|Open fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with moderate [1-24 hours] loss of consciousness
C0159526|ICD9CM|AB|804.93|Opn skul/oth fx-mod coma
C0159527|ICD9CM|PT|804.94|Open fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0159527|ICD9CM|AB|804.94|Opn skl/oth fx-prol coma
C0159528|ICD9CM|PT|804.95|Open fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0159528|ICD9CM|AB|804.95|Opn skl/oth fx-deep coma
C0159529|ICD9CM|PT|804.96|Open fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with loss of consciousness of unspecified duration
C0159529|ICD9CM|AB|804.96|Opn skul/oth fx-coma NOS
C0159530|ICD9CM|PT|804.99|Open fractures involving skull or face with other bones, with intracranial injury of other and unspecified nature, with concussion, unspecified
C0159530|ICD9CM|AB|804.99|Opn skull/oth fx-concuss
C0159533|ICD9CM|PT|805.01|Closed fracture of first cervical vertebra
C0159533|ICD9CM|AB|805.01|Fx c1 vertebra-closed
C0159534|ICD9CM|PT|805.02|Closed fracture of second cervical vertebra
C0159534|ICD9CM|AB|805.02|Fx c2 vertebra-closed
C0159535|ICD9CM|PT|805.03|Closed fracture of third cervical vertebra
C0159535|ICD9CM|AB|805.03|Fx c3 vertebra-closed
C0159536|ICD9CM|PT|805.04|Closed fracture of fourth cervical vertebra
C0159536|ICD9CM|AB|805.04|Fx c4 vertebra-closed
C0159537|ICD9CM|PT|805.05|Closed fracture of fifth cervical vertebra
C0159537|ICD9CM|AB|805.05|Fx c5 vertebra-closed
C0159538|ICD9CM|PT|805.06|Closed fracture of sixth cervical vertebra
C0159538|ICD9CM|AB|805.06|Fx c6 vertebra-closed
C0159539|ICD9CM|PT|805.07|Closed fracture of seventh cervical vertebra
C0159539|ICD9CM|AB|805.07|Fx c7 vertebra-closed
C0159540|ICD9CM|PT|805.08|Closed fracture of multiple cervical vertebrae
C0159540|ICD9CM|AB|805.08|Fx mult cervical vert-cl
C0159543|ICD9CM|PT|805.11|Open fracture of first cervical vertebra
C0159543|ICD9CM|AB|805.11|Fx c1 vertebra-open
C0159544|ICD9CM|PT|805.12|Open fracture of second cervical vertebra
C0159544|ICD9CM|AB|805.12|Fx c2 vertebra-open
C0159545|ICD9CM|PT|805.13|Open fracture of third cervical vertebra
C0159545|ICD9CM|AB|805.13|Fx c3 vertebra-open
C0159546|ICD9CM|PT|805.14|Open fracture of fourth cervical vertebra
C0159546|ICD9CM|AB|805.14|Fx c4 vertebra-open
C0159547|ICD9CM|PT|805.15|Open fracture of fifth cervical vertebra
C0159547|ICD9CM|AB|805.15|Fx c5 vertebra-open
C0159548|ICD9CM|PT|805.16|Open fracture of sixth cervical vertebra
C0159548|ICD9CM|AB|805.16|Fx c6 vertebra-open
C0159549|ICD9CM|PT|805.17|Open fracture of seventh cervical vertebra
C0159549|ICD9CM|AB|805.17|Fx c7 vertebra-open
C0159550|ICD9CM|PT|805.18|Open fracture of multiple cervical vertebrae
C0159550|ICD9CM|AB|805.18|Fx mlt cervical vert-opn
C0159551|ICD9CM|PT|805.2|Closed fracture of dorsal [thoracic] vertebra without mention of spinal cord injury
C0159551|ICD9CM|AB|805.2|Fx dorsal vertebra-close
C0159552|ICD9CM|PT|805.3|Open fracture of dorsal [thoracic] vertebra without mention of spinal cord injury
C0159552|ICD9CM|AB|805.3|Fx dorsal vertebra-open
C0159555|ICD9CM|PT|805.6|Closed fracture of sacrum and coccyx without mention of spinal cord injury
C0159555|ICD9CM|AB|805.6|Fx sacrum/coccyx-closed
C0159556|ICD9CM|PT|805.7|Open fracture of sacrum and coccyx without mention of spinal cord injury
C0159556|ICD9CM|AB|805.7|Fx sacrum/coccyx-open
C0159557|ICD9CM|PT|805.9|Open fracture of unspecified vertebral column without mention of spinal cord injury
C0159557|ICD9CM|AB|805.9|Vertebral fx NOS-open
C0159560|ICD9CM|PT|806.00|Closed fracture of C1-C4 level with unspecified spinal cord injury
C0159560|ICD9CM|AB|806.00|C1-c4 fx-cl/cord inj NOS
C0159562|ICD9CM|PT|806.02|Closed fracture of C1-C4 level with anterior cord syndrome
C0159562|ICD9CM|AB|806.02|C1-c4 fx-cl/ant cord syn
C0159563|ICD9CM|PT|806.03|Closed fracture of C1-C4 level with central cord syndrome
C0159563|ICD9CM|AB|806.03|C1-c4 fx-cl/cen cord syn
C0159564|ICD9CM|PT|806.04|Closed fracture of C1-C4 level with other specified spinal cord injury
C0159564|ICD9CM|AB|806.04|C1-c4 fx-cl/cord inj NEC
C0159565|ICD9CM|PT|806.05|Closed fracture of C5-C7 level with unspecified spinal cord injury
C0159565|ICD9CM|AB|806.05|C5-c7 fx-cl/cord inj NOS
C0159567|ICD9CM|PT|806.07|Closed fracture of C5-C7 level with anterior cord syndrome
C0159567|ICD9CM|AB|806.07|C5-c7 fx-cl/ant cord syn
C0159568|ICD9CM|PT|806.08|Closed fracture of C5-C7 level with central cord syndrome
C0159568|ICD9CM|AB|806.08|C5-c7 fx-cl/cen cord syn
C0159569|ICD9CM|PT|806.09|Closed fracture of C5-C7 level with other specified spinal cord injury
C0159569|ICD9CM|AB|806.09|C5-c7 fx-cl/cord inj NEC
C0159571|ICD9CM|PT|806.10|Open fracture of C1-C4 level with unspecified spinal cord injury
C0159571|ICD9CM|AB|806.10|C1-c4 fx-op/cord inj NOS
C0159573|ICD9CM|PT|806.12|Open fracture of C1-C4 level with anterior cord syndrome
C0159573|ICD9CM|AB|806.12|C1-c4 fx-op/ant cord syn
C0159574|ICD9CM|PT|806.13|Open fracture of C1-C4 level with central cord syndrome
C0159574|ICD9CM|AB|806.13|C1-c4 fx-op/cen cord syn
C0159575|ICD9CM|PT|806.14|Open fracture of C1-C4 level with other specified spinal cord injury
C0159575|ICD9CM|AB|806.14|C1-c4 fx-op/cord inj NEC
C0159576|ICD9CM|PT|806.15|Open fracture of C5-C7 level with unspecified spinal cord injury
C0159576|ICD9CM|AB|806.15|C5-c7 fx-op/cord inj NOS
C0159578|ICD9CM|PT|806.17|Open fracture of C5-C7 level with anterior cord syndrome
C0159578|ICD9CM|AB|806.17|C5-c7 fx-op/ant cord syn
C0159579|ICD9CM|PT|806.18|Open fracture of C5-C7 level with central cord syndrome
C0159579|ICD9CM|AB|806.18|C5-c7 fx-op/cen cord syn
C0159580|ICD9CM|PT|806.19|Open fracture of C5-C7 level with other specified spinal cord injury
C0159580|ICD9CM|AB|806.19|C5-c7 fx-op/cord inj NEC
C0159582|ICD9CM|PT|806.20|Closed fracture of T1-T6 level with unspecified spinal cord injury
C0159582|ICD9CM|AB|806.20|T1-t6 fx-cl/cord inj NOS
C0159584|ICD9CM|PT|806.22|Closed fracture of T1-T6 level with anterior cord syndrome
C0159584|ICD9CM|AB|806.22|T1-t6 fx-cl/ant cord syn
C0159585|ICD9CM|PT|806.23|Closed fracture of T1-T6 level with central cord syndrome
C0159585|ICD9CM|AB|806.23|T1-t6 fx-cl/cen cord syn
C0159586|ICD9CM|PT|806.24|Closed fracture of T1-T6 level with other specified spinal cord injury
C0159586|ICD9CM|AB|806.24|T1-t6 fx-cl/cord inj NEC
C0159587|ICD9CM|PT|806.25|Closed fracture of T7-T12 level with unspecified spinal cord injury
C0159587|ICD9CM|AB|806.25|T7-t12 fx-cl/crd inj NOS
C0159589|ICD9CM|PT|806.27|Closed fracture of T7-T12 level with anterior cord syndrome
C0159589|ICD9CM|AB|806.27|T7-t12 fx-cl/ant crd syn
C0159590|ICD9CM|PT|806.28|Closed fracture of T7-T12 level with central cord syndrome
C0159590|ICD9CM|AB|806.28|T7-t12 fx-cl/cen crd syn
C0159591|ICD9CM|PT|806.29|Closed fracture of T7-T12 level with other specified spinal cord injury
C0159591|ICD9CM|AB|806.29|T7-t12 fx-cl/crd inj NEC
C0159593|ICD9CM|PT|806.30|Open fracture of T1-T6 level with unspecified spinal cord injury
C0159593|ICD9CM|AB|806.30|T1-t6 fx-op/cord inj NOS
C0159595|ICD9CM|PT|806.32|Open fracture of T1-T6 level with anterior cord syndrome
C0159595|ICD9CM|AB|806.32|T1-t6 fx-op/ant cord syn
C0159596|ICD9CM|PT|806.33|Open fracture of T1-T6 level with central cord syndrome
C0159596|ICD9CM|AB|806.33|T1-t6 fx-op/cen cord syn
C0159597|ICD9CM|PT|806.34|Open fracture of T1-T6 level with other specified spinal cord injury
C0159597|ICD9CM|AB|806.34|T1-t6 fx-op/cord inj NEC
C0159598|ICD9CM|PT|806.35|Open fracture of T7-T12 level with unspecified spinal cord injury
C0159598|ICD9CM|AB|806.35|T7-t12 fx-op/crd inj NOS
C0159600|ICD9CM|PT|806.37|Open fracture of T7-T12 level with anterior cord syndrome
C0159600|ICD9CM|AB|806.37|T7-t12 fx-op/ant crd syn
C0159601|ICD9CM|PT|806.38|Open fracture of T7-T12 level with central cord syndrome
C0159601|ICD9CM|AB|806.38|T7-t12 fx-op/cen crd syn
C0159602|ICD9CM|PT|806.39|Open fracture of T7-T12 level with other specified spinal cord injury
C0159602|ICD9CM|AB|806.39|T7-t12 fx-op/crd inj NEC
C0159606|ICD9CM|HT|806.6|Closed fracture of sacrum and coccyx with spinal cord injury
C0159606|ICD9CM|PT|806.60|Closed fracture of sacrum and coccyx with unspecified spinal cord injury
C0159606|ICD9CM|AB|806.60|Fx sacrum-cl/crd inj NOS
C0159607|ICD9CM|PT|806.61|Closed fracture of sacrum and coccyx with complete cauda equina lesion
C0159607|ICD9CM|AB|806.61|Fx sacr-cl/cauda equ les
C0159608|ICD9CM|PT|806.62|Closed fracture of sacrum and coccyx with other cauda equina injury
C0159608|ICD9CM|AB|806.62|Fx sacr-cl/cauda inj NEC
C0159609|ICD9CM|PT|806.69|Closed fracture of sacrum and coccyx with other spinal cord injury
C0159609|ICD9CM|AB|806.69|Fx sacrum-cl/crd inj NEC
C0159611|ICD9CM|HT|806.7|Open fracture of sacrum and coccyx with spinal cord injury
C0159611|ICD9CM|PT|806.70|Open fracture of sacrum and coccyx with unspecified spinal cord injury
C0159611|ICD9CM|AB|806.70|Fx sacrum-op/crd inj NOS
C0159612|ICD9CM|PT|806.71|Open fracture of sacrum and coccyx with complete cauda equina lesion
C0159612|ICD9CM|AB|806.71|Fx sacr-op/cauda equ les
C0159613|ICD9CM|PT|806.72|Open fracture of sacrum and coccyx with other cauda equina injury
C0159613|ICD9CM|AB|806.72|Fx sacr-op/cauda inj NEC
C0159614|ICD9CM|PT|806.79|Open fracture of sacrum and coccyx with other spinal cord injury
C0159614|ICD9CM|AB|806.79|Fx sacrum-op/crd inj NEC
C0159615|ICD9CM|PT|806.8|Closed fracture of unspecified vertebral column with spinal cord injury
C0159615|ICD9CM|AB|806.8|Vert fx NOS-cl w crd inj
C0159616|ICD9CM|PT|806.9|Open fracture of unspecified vertebral column with spinal cord injury
C0159616|ICD9CM|AB|806.9|Vert fx NOS-op w crd inj
C0159617|ICD9CM|HT|807|Fracture of rib(s), sternum, larynx, and trachea
C0159618|ICD9CM|PT|807.01|Closed fracture of one rib
C0159618|ICD9CM|AB|807.01|Fracture one rib-closed
C0159619|ICD9CM|PT|807.02|Closed fracture of two ribs
C0159619|ICD9CM|AB|807.02|Fracture two ribs-closed
C0159620|ICD9CM|PT|807.03|Closed fracture of three ribs
C0159620|ICD9CM|AB|807.03|Fracture three ribs-clos
C0159621|ICD9CM|PT|807.04|Closed fracture of four ribs
C0159621|ICD9CM|AB|807.04|Fracture four ribs-close
C0159622|ICD9CM|PT|807.05|Closed fracture of five ribs
C0159622|ICD9CM|AB|807.05|Fracture five ribs-close
C0159623|ICD9CM|PT|807.06|Closed fracture of six ribs
C0159623|ICD9CM|AB|807.06|Fracture six ribs-closed
C0159624|ICD9CM|PT|807.07|Closed fracture of seven ribs
C0159624|ICD9CM|AB|807.07|Fracture seven ribs-clos
C0159625|ICD9CM|PT|807.08|Closed fracture of eight or more ribs
C0159625|ICD9CM|AB|807.08|Fx eight/more rib-closed
C0159626|ICD9CM|PT|807.09|Closed fracture of multiple ribs, unspecified
C0159626|ICD9CM|AB|807.09|Fx mult ribs NOS-closed
C0159628|ICD9CM|PT|807.11|Open fracture of one rib
C0159628|ICD9CM|AB|807.11|Fracture one rib-open
C0159629|ICD9CM|PT|807.12|Open fracture of two ribs
C0159629|ICD9CM|AB|807.12|Fracture two ribs-open
C0159630|ICD9CM|PT|807.13|Open fracture of three ribs
C0159630|ICD9CM|AB|807.13|Fracture three ribs-open
C0159631|ICD9CM|PT|807.14|Open fracture of four ribs
C0159631|ICD9CM|AB|807.14|Fracture four ribs-open
C0159632|ICD9CM|PT|807.15|Open fracture of five ribs
C0159632|ICD9CM|AB|807.15|Fracture five ribs-open
C0159633|ICD9CM|PT|807.16|Open fracture of six ribs
C0159633|ICD9CM|AB|807.16|Fracture six ribs-open
C0159634|ICD9CM|PT|807.17|Open fracture of seven ribs
C0159634|ICD9CM|AB|807.17|Fracture seven ribs-open
C0159635|ICD9CM|PT|807.18|Open fracture of eight or more ribs
C0159635|ICD9CM|AB|807.18|Fx eight/more ribs-open
C0159636|ICD9CM|PT|807.19|Open fracture of multiple ribs, unspecified
C0159636|ICD9CM|AB|807.19|Fx mult ribs NOS-open
C0159637|ICD9CM|PT|807.2|Closed fracture of sternum
C0159637|ICD9CM|AB|807.2|Fracture of sternum-clos
C0159638|ICD9CM|PT|807.3|Open fracture of sternum
C0159638|ICD9CM|AB|807.3|Fracture of sternum-open
C0159639|ICD9CM|PT|807.5|Closed fracture of larynx and trachea
C0159639|ICD9CM|AB|807.5|Fx larynx/trachea-closed
C0159640|ICD9CM|PT|807.6|Open fracture of larynx and trachea
C0159640|ICD9CM|AB|807.6|Fx larynx/trachea-open
C0159641|ICD9CM|PT|808.0|Closed fracture of acetabulum
C0159641|ICD9CM|AB|808.0|Fracture acetabulum-clos
C0159642|ICD9CM|PT|808.1|Open fracture of acetabulum
C0159642|ICD9CM|AB|808.1|Fracture acetabulum-open
C0159643|ICD9CM|PT|808.2|Closed fracture of pubis
C0159643|ICD9CM|AB|808.2|Fracture of pubis-closed
C0159644|ICD9CM|PT|808.3|Open fracture of pubis
C0159644|ICD9CM|AB|808.3|Fracture of pubis-open
C0159645|ICD9CM|HT|808.4|Closed fracture of other specified part of pelvis
C0159645|ICD9CM|PT|808.49|Closed fracture of other specified part of pelvis
C0159645|ICD9CM|AB|808.49|Pelvic fracture NEC-clos
C0159646|ICD9CM|PT|808.41|Closed fracture of ilium
C0159646|ICD9CM|AB|808.41|Fracture of ilium-closed
C0159647|ICD9CM|PT|808.42|Closed fracture of ischium
C0159647|ICD9CM|AB|808.42|Fracture ischium-closed
C0159649|ICD9CM|HT|808.5|Open fracture of other specified part of pelvis
C0159649|ICD9CM|PT|808.59|Open fracture of other specified part of pelvis
C0159649|ICD9CM|AB|808.59|Pelvic fracture NEC-open
C0159651|ICD9CM|PT|808.52|Open fracture of ischium
C0159651|ICD9CM|AB|808.52|Fracture of ischium-open
C0159655|ICD9CM|HT|809|Ill-defined fractures of bones of trunk
C0159656|ICD9CM|PT|809.0|Fracture of bones of trunk, closed
C0159656|ICD9CM|AB|809.0|Fracture trunk bone-clos
C0159657|ICD9CM|PT|809.1|Fracture of bones of trunk, open
C0159657|ICD9CM|AB|809.1|Fracture trunk bone-open
C0159658|ICD9CM|HT|810|Fracture of clavicle
C0159659|ICD9CM|HT|810.0|Closed fracture of clavicle
C0159659|ICD9CM|PT|810.00|Closed fracture of clavicle, unspecified part
C0159659|ICD9CM|AB|810.00|Fx clavicle NOS-closed
C0159661|ICD9CM|PT|810.02|Closed fracture of shaft of clavicle
C0159661|ICD9CM|AB|810.02|Fx clavicle shaft-closed
C0159663|ICD9CM|HT|810.1|Open fracture of clavicle
C0159663|ICD9CM|PT|810.10|Open fracture of clavicle, unspecified part
C0159663|ICD9CM|AB|810.10|Fx clavicle NOS-open
C0159665|ICD9CM|PT|810.12|Open fracture of shaft of clavicle
C0159665|ICD9CM|AB|810.12|Fx clavicle shaft-open
C0159667|ICD9CM|HT|811|Fracture of scapula
C0159668|ICD9CM|PT|811.00|Closed fracture of scapula, unspecified part
C0159668|ICD9CM|HT|811.0|Closed fracture of scapula
C0159668|ICD9CM|AB|811.00|Fx scapula NOS-closed
C0159669|ICD9CM|PT|811.01|Closed fracture of acromial process of scapula
C0159669|ICD9CM|AB|811.01|Fx scapul, acrom proc-cl
C0159671|ICD9CM|PT|811.03|Closed fracture of glenoid cavity and neck of scapula
C0159671|ICD9CM|AB|811.03|Fx scap, glen cav/nck-cl
C0159672|ICD9CM|PT|811.09|Closed fracture of scapula, other
C0159672|ICD9CM|AB|811.09|Fx scapula NEC-closed
C0159673|ICD9CM|HT|811.1|Open fracture of scapula
C0159673|ICD9CM|PT|811.10|Open fracture of scapula, unspecified part
C0159673|ICD9CM|AB|811.10|Fx scapula NOS-open
C0159674|ICD9CM|PT|811.11|Open fracture of acromial process of scapula
C0159674|ICD9CM|AB|811.11|Fx scapul, acrom proc-op
C0159675|ICD9CM|PT|811.12|Open fracture of coracoid process
C0159675|ICD9CM|AB|811.12|Fx scapul, corac proc-op
C0159677|ICD9CM|PT|811.19|Open fracture of scapula, other
C0159677|ICD9CM|AB|811.19|Fx scapula NEC-open
C0159678|ICD9CM|HT|812.0|Fracture of upper end of humerus, closed
C0159679|ICD9CM|PT|812.00|Closed fracture of unspecified part of upper end of humerus
C0159679|ICD9CM|AB|812.00|Fx up end humerus NOS-cl
C0159680|ICD9CM|PT|812.01|Closed fracture of surgical neck of humerus
C0159680|ICD9CM|AB|812.01|Fx surg nck humerus-clos
C0159683|ICD9CM|PT|812.09|Other closed fracture of upper end of humerus
C0159683|ICD9CM|AB|812.09|Fx upper humerus NEC-cl
C0159684|ICD9CM|HT|812.1|Fracture of upper end of humerus, open
C0159685|ICD9CM|PT|812.10|Open fracture of unspecified part of upper end of humerus
C0159685|ICD9CM|AB|812.10|Fx upper humerus NOS-opn
C0159686|ICD9CM|PT|812.11|Open fracture of surgical neck of humerus
C0159686|ICD9CM|AB|812.11|Fx surg neck humerus-opn
C0159689|ICD9CM|PT|812.19|Other open fracture of upper end of humerus
C0159689|ICD9CM|AB|812.19|Fx upper humerus NEC-opn
C0159690|ICD9CM|HT|812.2|Closed fracture of shaft or unspecified part of humerus
C0159692|ICD9CM|PT|812.21|Closed fracture of shaft of humerus
C0159692|ICD9CM|AB|812.21|Fx humerus shaft-closed
C0159693|ICD9CM|HT|812.3|Fracture of shaft or unspecified part of humerus, open
C0159695|ICD9CM|PT|812.31|Open fracture of shaft of humerus
C0159695|ICD9CM|AB|812.31|Fx humerus shaft-open
C0159701|ICD9CM|PT|812.44|Closed fracture of unspecified condyle(s) of humerus
C0159701|ICD9CM|AB|812.44|Fx humer, condyl NOS-cl
C0159702|ICD9CM|PT|812.49|Other closed fracture of lower end of humerus
C0159702|ICD9CM|AB|812.49|Fx lower humerus NEC-cl
C0159708|ICD9CM|PT|812.54|Open fracture of unspecified condyle(s) of humerus
C0159708|ICD9CM|AB|812.54|Fx humer, condyl NOS-opn
C0159709|ICD9CM|PT|812.59|Other open fracture of lower end of humerus
C0159709|ICD9CM|AB|812.59|Fx lower humer NEC-open
C0159710|ICD9CM|HT|813|Fracture of radius and ulna
C0159713|ICD9CM|PT|813.01|Closed fracture of olecranon process of ulna
C0159713|ICD9CM|AB|813.01|Fx olecran proc ulna-cl
C0159715|ICD9CM|PT|813.04|Other and unspecified closed fractures of proximal end of ulna (alone)
C0159715|ICD9CM|AB|813.04|Fx upper ulna NEC/NOS-cl
C0159716|ICD9CM|PT|813.05|Closed fracture of head of radius
C0159716|ICD9CM|AB|813.05|Fx radius head-closed
C0159717|ICD9CM|PT|813.06|Closed fracture of neck of radius
C0159717|ICD9CM|AB|813.06|Fx radius neck-closed
C0159718|ICD9CM|PT|813.07|Other and unspecified closed fractures of proximal end of radius (alone)
C0159718|ICD9CM|AB|813.07|Fx up radius NEC/NOS-cl
C0159720|ICD9CM|HT|813.1|Fracture of upper end of radius and ulna, open
C0159720|ICD9CM|PT|813.18|Open fracture of radius with ulna, upper end (any part)
C0159720|ICD9CM|AB|813.18|Fx up radius w ulna-open
C0159722|ICD9CM|PT|813.11|Open fracture of olecranon process of ulna
C0159722|ICD9CM|AB|813.11|Fx olecran proc ulna-opn
C0159723|ICD9CM|PT|813.12|Open fracture of coronoid process of ulna
C0159723|ICD9CM|AB|813.12|Fx coronoid pro ulna-opn
C0159724|ICD9CM|PT|813.13|Open Monteggia's fracture
C0159724|ICD9CM|AB|813.13|Monteggia's fx-open
C0159725|ICD9CM|PT|813.14|Other and unspecified open fractures of proximal end of ulna (alone)
C0159725|ICD9CM|AB|813.14|Fx up ulna NEC/NOS-open
C0159726|ICD9CM|PT|813.15|Open fracture of head of radius
C0159726|ICD9CM|AB|813.15|Fx radius head-open
C0159727|ICD9CM|PT|813.16|Open fracture of neck of radius
C0159727|ICD9CM|AB|813.16|Fx radius neck-open
C0159728|ICD9CM|PT|813.17|Other and unspecified open fractures of proximal end of radius (alone)
C0159728|ICD9CM|AB|813.17|Fx up radius NEC/NOS-opn
C0159730|ICD9CM|HT|813.2|Fracture of shaft of radius and ulna, closed
C0159730|ICD9CM|PT|813.23|Closed fracture of shaft of radius with ulna
C0159730|ICD9CM|AB|813.23|Fx shaft rad w ulna-clos
C0159731|ICD9CM|PT|813.20|Closed fracture of shaft of radius or ulna, unspecified
C0159731|ICD9CM|AB|813.20|Fx shaft forearm NOS-cl
C0159733|ICD9CM|PT|813.22|Closed fracture of shaft of ulna (alone)
C0159733|ICD9CM|AB|813.22|Fx ulna shaft-closed
C0159734|ICD9CM|HT|813.3|Fracture of shaft of radius and ulna, open
C0159734|ICD9CM|PT|813.33|Open fracture of shaft of radius with ulna
C0159734|ICD9CM|AB|813.33|Fx shaft rad w ulna-open
C0159735|ICD9CM|PT|813.30|Open fracture of shaft of radius or ulna, unspecified
C0159735|ICD9CM|AB|813.30|Fx shaft forearm NOS-opn
C0159737|ICD9CM|PT|813.32|Open fracture of shaft of ulna (alone)
C0159737|ICD9CM|AB|813.32|Fx ulna shaft-open
C0159738|ICD9CM|HT|813.4|Fracture of lower end of radius and ulna, closed
C0159738|ICD9CM|PT|813.44|Closed fracture of lower end of radius with ulna
C0159738|ICD9CM|AB|813.44|Fx low radius w ulna-cl
C0159739|ICD9CM|PT|813.40|Closed fracture of lower end of forearm, unspecified
C0159739|ICD9CM|AB|813.40|Fx lower forearm NOS-cl
C0159740|ICD9CM|PT|813.42|Other closed fractures of distal end of radius (alone)
C0159740|ICD9CM|AB|813.42|Fx distal radius NEC-cl
C0159742|ICD9CM|HT|813.5|Fracture of lower end of radius and ulna, open
C0159742|ICD9CM|PT|813.54|Open fracture of lower end of radius with ulna
C0159742|ICD9CM|AB|813.54|Fx low radius w ulna-opn
C0159743|ICD9CM|PT|813.50|Open fracture of lower end of forearm, unspecified
C0159743|ICD9CM|AB|813.50|Fx lower forearm NOS-opn
C0159744|ICD9CM|PT|813.51|Open Colles' fracture
C0159744|ICD9CM|AB|813.51|Colles' fracture-open
C0159745|ICD9CM|PT|813.52|Other open fractures of distal end of radius (alone)
C0159745|ICD9CM|AB|813.52|Fx distal radius NEC-opn
C0159746|ICD9CM|PT|813.53|Open fracture of distal end of ulna (alone)
C0159746|ICD9CM|AB|813.53|Fx distal ulna-open
C0159747|ICD9CM|PT|813.83|Closed fracture of unspecified part of radius with ulna
C0159747|ICD9CM|HT|813.8|Fracture of unspecified part of radius with ulna, closed
C0159747|ICD9CM|AB|813.83|Fx radius w ulna NOS-cl
C0159748|ICD9CM|PT|813.80|Closed fracture of unspecified part of forearm
C0159748|ICD9CM|AB|813.80|Fx forearm NOS-closed
C0159749|ICD9CM|PT|813.93|Open fracture of unspecified part of radius with ulna
C0159749|ICD9CM|HT|813.9|Fracture of unspecified part of radius with ulna, open
C0159749|ICD9CM|AB|813.93|Fx radius w ulna NOS-opn
C0159750|ICD9CM|PT|813.90|Open fracture of unspecified part of forearm
C0159750|ICD9CM|AB|813.90|Fx forearm NOS-open
C0159751|ICD9CM|PT|813.91|Open fracture of unspecified part of radius (alone)
C0159751|ICD9CM|AB|813.91|Fracture radius NOS-open
C0159752|ICD9CM|PT|813.92|Open fracture of unspecified part of ulna (alone)
C0159752|ICD9CM|AB|813.92|Fracture ulna NOS-open
C0159758|ICD9CM|PT|814.04|Closed fracture of pisiform bone of wrist
C0159758|ICD9CM|AB|814.04|Fx pisiform-closed
C0159763|ICD9CM|PT|814.09|Closed fracture of other bone of wrist
C0159763|ICD9CM|AB|814.09|Fx carpal bone NEC-close
C0159765|ICD9CM|PT|814.10|Open fracture of carpal bone, unspecified
C0159765|ICD9CM|HT|814.1|Open fractures of carpal bones
C0159765|ICD9CM|AB|814.10|Fx carpal bone NOS-open
C0159769|ICD9CM|PT|814.14|Open fracture of pisiform bone of wrist
C0159769|ICD9CM|AB|814.14|Fx pisiform-open
C0159774|ICD9CM|PT|814.19|Open fracture of other bone of wrist
C0159774|ICD9CM|AB|814.19|Fx carpal bone NEC-open
C0159776|ICD9CM|HT|815.0|Closed fracture of metacarpal bones
C0159776|ICD9CM|PT|815.00|Closed fracture of metacarpal bone(s), site unspecified
C0159776|ICD9CM|AB|815.00|Fx metacarpal NOS-closed
C0159783|ICD9CM|HT|815.1|Open fracture of metacarpal bones
C0159783|ICD9CM|PT|815.10|Open fracture of metacarpal bone(s), site unspecified
C0159783|ICD9CM|AB|815.10|Fx metacarpal NOS-open
C0159790|ICD9CM|HT|816|Fracture of one or more phalanges of hand
C0159791|ICD9CM|HT|816.0|Closed fracture of one or more phalanges of hand
C0159791|ICD9CM|PT|816.00|Closed fracture of phalanx or phalanges of hand, unspecified
C0159791|ICD9CM|AB|816.00|Fx phalanx, hand NOS-cl
C0159793|ICD9CM|PT|816.01|Closed fracture of middle or proximal phalanx or phalanges of hand
C0159793|ICD9CM|AB|816.01|Fx mid/prx phal, hand-cl
C0159794|ICD9CM|PT|816.02|Closed fracture of distal phalanx or phalanges of hand
C0159794|ICD9CM|AB|816.02|Fx dist phalanx, hand-cl
C0159795|ICD9CM|PT|816.03|Closed fracture of multiple sites of phalanx or phalanges of hand
C0159795|ICD9CM|AB|816.03|Fx mult phalan, hand-cl
C0159796|ICD9CM|HT|816.1|Open fracture of one or more phalanges of hand
C0159796|ICD9CM|PT|816.10|Open fracture of phalanx or phalanges of hand, unspecified
C0159796|ICD9CM|AB|816.10|Fx phalanx, hand NOS-opn
C0159798|ICD9CM|PT|816.11|Open fracture of middle or proximal phalanx or phalanges of hand
C0159798|ICD9CM|AB|816.11|Fx mid/prx phal, hand-op
C0159799|ICD9CM|PT|816.12|Open fracture of distal phalanx or phalanges of hand
C0159799|ICD9CM|AB|816.12|Fx distal phal, hand-opn
C0159800|ICD9CM|PT|816.13|Open fracture of multiple sites of phalanx or phalanges of hand
C0159800|ICD9CM|AB|816.13|Fx mult phalan, hand-opn
C0159801|ICD9CM|HT|817|Multiple fractures of hand bones
C0159802|ICD9CM|PT|817.0|Multiple closed fractures of hand bones
C0159802|ICD9CM|AB|817.0|Multiple fx hand-closed
C0159803|ICD9CM|PT|817.1|Multiple open fractures of hand bones
C0159803|ICD9CM|AB|817.1|Multiple fx hand-open
C0159804|ICD9CM|HT|818|Ill-defined fractures of upper limb
C0159805|ICD9CM|PT|818.0|Ill-defined closed fractures of upper limb
C0159805|ICD9CM|AB|818.0|Fx arm mult/NOS-closed
C0159806|ICD9CM|PT|818.1|Ill-defined open fractures of upper limb
C0159806|ICD9CM|AB|818.1|Fx arm mult/NOS-open
C0159807|ICD9CM|HT|819|Multiple fractures involving both upper limbs, and upper limb with rib(s) and sternum
C0159808|ICD9CM|PT|819.0|Multiple closed fractures involving both upper limbs, and upper limb with rib(s) and sternum
C0159808|ICD9CM|AB|819.0|Fx arms w rib/sternum-cl
C0159809|ICD9CM|PT|819.1|Multiple open fractures involving both upper limbs, and upper limb with rib(s) and sternum
C0159809|ICD9CM|AB|819.1|Fx arms w rib/stern-open
C0159810|ICD9CM|HT|820.0|Transcervical fracture, closed
C0159811|ICD9CM|PT|820.00|Closed fracture of intracapsular section of neck of femur, unspecified
C0159811|ICD9CM|AB|820.00|Fx femur intrcaps NOS-cl
C0159812|ICD9CM|PT|820.01|Closed fracture of epiphysis (separation) (upper) of neck of femur
C0159812|ICD9CM|AB|820.01|Fx up femur epiphy-clos
C0159813|ICD9CM|PT|820.02|Closed fracture of midcervical section of neck of femur
C0159813|ICD9CM|AB|820.02|Fx femur, midcervic-clos
C0159814|ICD9CM|PT|820.03|Closed fracture of base of neck of femur
C0159814|ICD9CM|AB|820.03|Fx base femoral nck-clos
C0159815|ICD9CM|PT|820.09|Other closed transcervical fracture of neck of femur
C0159815|ICD9CM|AB|820.09|Fx femur intrcaps NEC-cl
C0159816|ICD9CM|HT|820.1|Transcervical fracture, open
C0159817|ICD9CM|PT|820.10|Open fracture of intracapsular section of neck of femur, unspecified
C0159817|ICD9CM|AB|820.10|Fx femur intrcap NOS-opn
C0159818|ICD9CM|PT|820.11|Open fracture of epiphysis (separation) (upper) of neck of femur
C0159818|ICD9CM|AB|820.11|Fx up femur epiphy-open
C0159819|ICD9CM|PT|820.12|Open fracture of midcervical section of neck of femur
C0159819|ICD9CM|AB|820.12|Fx femur, midcervic-open
C0159820|ICD9CM|PT|820.13|Open fracture of base of neck of femur
C0159820|ICD9CM|AB|820.13|Fx base femoral nck-open
C0159821|ICD9CM|PT|820.19|Other open transcervical fracture of neck of femur
C0159821|ICD9CM|AB|820.19|Fx femur intrcap NEC-opn
C0159822|ICD9CM|HT|820.2|Pertrochanteric fracture of femur, closed
C0159823|ICD9CM|PT|820.20|Closed fracture of trochanteric section of neck of femur
C0159823|ICD9CM|AB|820.20|Trochanteric fx NOS-clos
C0159824|ICD9CM|PT|820.21|Closed fracture of intertrochanteric section of neck of femur
C0159824|ICD9CM|AB|820.21|Intertrochanteric fx-cl
C0159826|ICD9CM|HT|820.3|Pertrochanteric fracture of femur, open
C0159827|ICD9CM|PT|820.30|Open fracture of trochanteric section of neck of femur, unspecified
C0159827|ICD9CM|AB|820.30|Trochanteric fx NOS-open
C0159828|ICD9CM|PT|820.31|Open fracture of intertrochanteric section of neck of femur
C0159828|ICD9CM|AB|820.31|Intertrochanteric fx-opn
C0159831|ICD9CM|HT|821|Fracture of other and unspecified parts of femur
C0159832|ICD9CM|HT|821.0|Fracture of shaft or unspecified part of femur, closed
C0159833|ICD9CM|PT|821.01|Closed fracture of shaft of femur
C0159833|ICD9CM|AB|821.01|Fx femur shaft-closed
C0159834|ICD9CM|HT|821.1|Fracture of shaft or unspecified part of femur, open
C0159835|ICD9CM|PT|821.10|Open fracture of unspecified part of femur
C0159835|ICD9CM|AB|821.10|Fx femur NOS-open
C0159836|ICD9CM|PT|821.11|Open fracture of shaft of femur
C0159836|ICD9CM|AB|821.11|Fx femur shaft-open
C0159837|ICD9CM|HT|821.2|Fracture of lower end of femur, closed
C0159838|ICD9CM|PT|821.20|Closed fracture of lower end of femur, unspecified part
C0159838|ICD9CM|AB|821.20|Fx low end femur NOS-cl
C0159840|ICD9CM|PT|821.22|Closed fracture of epiphysis, lower (separation) of femur
C0159840|ICD9CM|AB|821.22|Fx low femur epiphy-clos
C0159842|ICD9CM|PT|821.29|Other closed fracture of lower end of femur
C0159842|ICD9CM|AB|821.29|Fx low end femur NEC-cl
C0159843|ICD9CM|HT|821.3|Fracture of lower end of femur, open
C0159844|ICD9CM|PT|821.30|Open fracture of lower end of femur, unspecified part
C0159844|ICD9CM|AB|821.30|Fx low end femur NOS-opn
C0159846|ICD9CM|PT|821.32|Open fracture of epiphysis. Lower (separation) of femur
C0159846|ICD9CM|AB|821.32|Fx low femur epiphy-open
C0159848|ICD9CM|PT|821.39|Other open fracture of lower end of femur
C0159848|ICD9CM|AB|821.39|Fx low end femur NEC-opn
C0159849|ICD9CM|HT|822|Fracture of patella
C0159850|ICD9CM|PT|822.0|Closed fracture of patella
C0159850|ICD9CM|AB|822.0|Fracture patella-closed
C0159851|ICD9CM|PT|822.1|Open fracture of patella
C0159851|ICD9CM|AB|822.1|Fracture patella-open
C0159852|ICD9CM|HT|823|Fracture of tibia and fibula
C0159854|ICD9CM|PT|823.00|Closed fracture of upper end of tibia alone
C0159854|ICD9CM|AB|823.00|Fx upper end tibia-close
C0159858|ICD9CM|PT|823.10|Open fracture of upper end of tibia alone
C0159858|ICD9CM|AB|823.10|Fx upper end tibia-open
C0159862|ICD9CM|PT|823.20|Closed fracture of shaft of tibia alone
C0159862|ICD9CM|AB|823.20|Fx shaft tibia-closed
C0159863|ICD9CM|PT|823.21|Closed fracture of shaft of fibula alone
C0159863|ICD9CM|AB|823.21|Fx shaft fibula-closed
C0159864|ICD9CM|HT|823.2|Fracture of shaft of tibia and fibula, closed
C0159864|ICD9CM|PT|823.22|Closed fracture of shaft of fibula with tibia
C0159864|ICD9CM|AB|823.22|Fx shaft fib w tib-clos
C0159866|ICD9CM|PT|823.30|Open fracture of shaft of tibia alone
C0159866|ICD9CM|AB|823.30|Fx tibia shaft-open
C0159867|ICD9CM|PT|823.31|Open fracture of shaft of fibula alone
C0159867|ICD9CM|AB|823.31|Fx fibula shaft-open
C0159868|ICD9CM|HT|823.3|Fracture of shaft of tibia and fibula, open
C0159868|ICD9CM|PT|823.32|Open fracture of shaft of fibula with tibia
C0159868|ICD9CM|AB|823.32|Fx shaft tibia w fib-opn
C0159870|ICD9CM|PT|823.80|Closed fracture of unspecified part of tibia alone
C0159870|ICD9CM|AB|823.80|Fx tibia NOS-closed
C0159871|ICD9CM|PT|823.81|Closed fracture of unspecified part of fibula alone
C0159871|ICD9CM|AB|823.81|Fx fibula NOS-closed
C0159874|ICD9CM|PT|823.90|Open fracture of unspecified part of tibia alone
C0159874|ICD9CM|AB|823.90|Fx tibia NOS-open
C0159875|ICD9CM|PT|823.91|Open fracture of unspecified part of fibula alone
C0159875|ICD9CM|AB|823.91|Fx fibula NOS-open
C0159876|ICD9CM|PT|823.92|Open fracture of unspecified part of fibula with tibia
C0159876|ICD9CM|HT|823.9|Fracture of unspecified part of tibia and fibula, open
C0159876|ICD9CM|AB|823.92|Fx tibia w fib NOS-open
C0159877|ICD9CM|HT|824|Fracture of ankle
C0159882|ICD9CM|PT|824.5|Bimalleolar fracture, open
C0159882|ICD9CM|AB|824.5|Fx bimalleolar-open
C0159883|ICD9CM|PT|824.6|Trimalleolar fracture, closed
C0159883|ICD9CM|AB|824.6|Fx trimalleolar-closed
C0159884|ICD9CM|PT|824.7|Trimalleolar fracture, open
C0159884|ICD9CM|AB|824.7|Fx trimalleolar-open
C0159888|ICD9CM|PT|825.0|Fracture of calcaneus, closed
C0159888|ICD9CM|AB|825.0|Fracture calcaneus-close
C0159889|ICD9CM|PT|825.1|Fracture of calcaneus, open
C0159889|ICD9CM|AB|825.1|Fracture calcaneus-open
C0159890|ICD9CM|PT|825.29|Other closed fracture of tarsal and metatarsal bones
C0159890|ICD9CM|HT|825.2|Fracture of other tarsal and metatarsal bones, closed
C0159890|ICD9CM|AB|825.29|Fx foot bone NEC-closed
C0159892|ICD9CM|PT|825.21|Closed fracture of astragalus
C0159892|ICD9CM|AB|825.21|Fx astragalus-closed
C0159899|ICD9CM|PT|825.31|Open fracture of astragalus
C0159899|ICD9CM|AB|825.31|Fx astragalus-open
C0159904|ICD9CM|PT|825.39|Other open fracture of tarsal and metatarsal bones
C0159904|ICD9CM|HT|825.3|Fracture of other tarsal and metatarsal bones, open
C0159904|ICD9CM|AB|825.39|Fx foot bone NEC-open
C0159905|ICD9CM|HT|826|Fracture of one or more phalanges of foot
C0159906|ICD9CM|PT|826.0|Closed fracture of one or more phalanges of foot
C0159906|ICD9CM|AB|826.0|Fx phalanx, foot-closed
C0159907|ICD9CM|PT|826.1|Open fracture of one or more phalanges of foot
C0159907|ICD9CM|AB|826.1|Fx phalanx, foot-open
C0159908|ICD9CM|HT|827|Other, multiple, and ill-defined fractures of lower limb
C0159909|ICD9CM|PT|827.0|Other, multiple and ill-defined fractures of lower limb, closed
C0159909|ICD9CM|AB|827.0|Fx lower limb NEC-closed
C0159910|ICD9CM|PT|827.1|Other, multiple and ill-defined fractures of lower limb, open
C0159910|ICD9CM|AB|827.1|Fx lower limb NEC-open
C0159911|ICD9CM|HT|828|Multiple fractures involving both lower limbs, lower with upper limb, and lower limb(s) with rib(s) and sternum
C0159912|ICD9CM|PT|828.0|Closed multiple fractures involving both lower limbs, lower with upper limb, and lower limb(s) with rib(s) and sternum
C0159912|ICD9CM|AB|828.0|Fx legs w arm/rib-closed
C0159913|ICD9CM|PT|828.1|Open multiple fractures involving both lower limbs, lower with upper limb, and lower limb(s) with rib(s) and sternum
C0159913|ICD9CM|AB|828.1|Fx legs w arm/rib-open
C0159914|ICD9CM|HT|830|Dislocation of jaw
C0159915|ICD9CM|PT|830.0|Closed dislocation of jaw
C0159915|ICD9CM|AB|830.0|Dislocation jaw-closed
C0159916|ICD9CM|PT|830.1|Open dislocation of jaw
C0159916|ICD9CM|AB|830.1|Dislocation jaw-open
C0159917|ICD9CM|PT|831.01|Closed anterior dislocation of humerus
C0159917|ICD9CM|AB|831.01|Ant disloc humerus-close
C0159918|ICD9CM|PT|831.02|Closed posterior dislocation of humerus
C0159918|ICD9CM|AB|831.02|Post disloc humerus-clos
C0159919|ICD9CM|PT|831.03|Closed inferior dislocation of humerus
C0159919|ICD9CM|AB|831.03|Infer disloc humerus-cl
C0159920|ICD9CM|PT|831.04|Closed dislocation of acromioclavicular (joint)
C0159920|ICD9CM|AB|831.04|Disloc acromioclavic-cl
C0159921|ICD9CM|PT|831.09|Closed dislocation of shoulder, other
C0159921|ICD9CM|AB|831.09|Disloc shoulder NEC-clos
C0159926|ICD9CM|PT|831.14|Open dislocation of acromioclavicular (joint)
C0159926|ICD9CM|AB|831.14|Disloc acromioclavic-opn
C0159927|ICD9CM|PT|831.19|Open dislocation of shoulder, other
C0159927|ICD9CM|AB|831.19|Disloc shoulder NEC-open
C0159930|ICD9CM|PT|832.01|Closed anterior dislocation of elbow
C0159930|ICD9CM|AB|832.01|Ant disloc elbow-closed
C0159931|ICD9CM|PT|832.02|Closed posterior dislocation of elbow
C0159931|ICD9CM|AB|832.02|Post disloc elbow-closed
C0159932|ICD9CM|PT|832.03|Closed medial dislocation of elbow
C0159932|ICD9CM|AB|832.03|Med disloc elbow-closed
C0159933|ICD9CM|PT|832.04|Closed lateral dislocation of elbow
C0159933|ICD9CM|AB|832.04|Lat disloc elbow-closed
C0159934|ICD9CM|PT|832.09|Closed dislocation of elbow, other
C0159934|ICD9CM|AB|832.09|Dislocat elbow NEC-close
C0159940|ICD9CM|PT|832.19|Open dislocation of elbow, other
C0159940|ICD9CM|AB|832.19|Dislocat elbow NEC-open
C0159942|ICD9CM|HT|833.0|Closed dislocation of wrist
C0159942|ICD9CM|PT|833.00|Closed dislocation of wrist, unspecified part
C0159942|ICD9CM|AB|833.00|Disloc wrist NOS-closed
C0159943|ICD9CM|PT|833.01|Closed dislocation of radioulnar (joint), distal
C0159943|ICD9CM|AB|833.01|Disloc dist radiouln-cl
C0159944|ICD9CM|PT|833.02|Closed dislocation of radiocarpal (joint)
C0159944|ICD9CM|AB|833.02|Disloc radiocarpal-clos
C0159945|ICD9CM|PT|833.03|Closed dislocation of midcarpal (joint)
C0159945|ICD9CM|AB|833.03|Disloca midcarpal-closed
C0159946|ICD9CM|PT|833.04|Closed dislocation of carpometacarpal (joint)
C0159946|ICD9CM|AB|833.04|Disloc carpometacarp-cl
C0159947|ICD9CM|PT|833.05|Closed dislocation of metacarpal (bone), proximal end
C0159947|ICD9CM|AB|833.05|Disloc metacarpal-closed
C0159948|ICD9CM|PT|833.09|Closed dislocation of wrist, other
C0159948|ICD9CM|AB|833.09|Disloc wrist NEC-closed
C0159950|ICD9CM|PT|833.11|Open dislocation of radioulnar (joint), distal
C0159950|ICD9CM|AB|833.11|Disloc dist radiouln-opn
C0159951|ICD9CM|PT|833.12|Open dislocation of radiocarpal (joint)
C0159951|ICD9CM|AB|833.12|Disloc radiocarpal-open
C0159952|ICD9CM|PT|833.13|Open dislocation of midcarpal (joint)
C0159952|ICD9CM|AB|833.13|Dislocat midcarpal-open
C0159953|ICD9CM|PT|833.14|Open dislocation of carpometacarpal (joint)
C0159953|ICD9CM|AB|833.14|Disloc carpometacarp-opn
C0159955|ICD9CM|PT|833.19|Open dislocation of wrist, other
C0159955|ICD9CM|AB|833.19|Dislocat wrist NEC-open
C0159956|ICD9CM|HT|834|Dislocation of finger
C0159957|ICD9CM|HT|834.0|Closed dislocation of finger
C0159960|ICD9CM|HT|834.1|Open dislocation of finger
C0159961|ICD9CM|PT|834.11|Open dislocation of metacarpophalangeal (joint)
C0159961|ICD9CM|AB|834.11|Disl metacarpophalan-opn
C0159962|ICD9CM|PT|834.12|Open dislocation interphalangeal (joint), hand
C0159962|ICD9CM|AB|834.12|Disl interphaln hand-opn
C0159963|ICD9CM|PT|835.01|Closed posterior dislocation of hip
C0159963|ICD9CM|AB|835.01|Posterior disloc hip-cl
C0159964|ICD9CM|PT|835.02|Closed obturator dislocation of hip
C0159964|ICD9CM|AB|835.02|Obturator disloc hip-cl
C0159965|ICD9CM|PT|835.03|Other closed anterior dislocation of hip
C0159965|ICD9CM|AB|835.03|Ant disloc hip NEC-clos
C0159968|ICD9CM|PT|835.12|Open obturator dislocation of hip
C0159968|ICD9CM|AB|835.12|Obturator disloc hip-opn
C0159969|ICD9CM|PT|835.13|Other open anterior dislocation of hip
C0159969|ICD9CM|AB|835.13|Ant disloc hip NEC-open
C0159970|ICD9CM|HT|836|Dislocation of knee
C0159973|ICD9CM|PT|836.2|Other tear of cartilage or meniscus of knee, current
C0159973|ICD9CM|AB|836.2|Tear meniscus NEC-curren
C0159975|ICD9CM|PT|836.4|Dislocation of patella, open
C0159975|ICD9CM|AB|836.4|Dislocation patella-open
C0159976|ICD9CM|HT|836.5|Other dislocation of knee, closed
C0159976|ICD9CM|PT|836.59|Other dislocation of knee, closed
C0159976|ICD9CM|AB|836.59|Dislocat knee NEC-closed
C0159978|ICD9CM|PT|836.51|Anterior dislocation of tibia, proximal end, closed
C0159978|ICD9CM|AB|836.51|Ant disloc prox tibia-cl
C0159979|ICD9CM|PT|836.52|Posterior dislocation of tibia, proximal end, closed
C0159979|ICD9CM|AB|836.52|Post disl prox tibia-cl
C0159980|ICD9CM|PT|836.53|Medial dislocation of tibia, proximal end, closed
C0159980|ICD9CM|AB|836.53|Med disloc prox tibia-cl
C0159981|ICD9CM|PT|836.54|Lateral dislocation of tibia, proximal end, closed
C0159981|ICD9CM|AB|836.54|Lat disloc prox tibia-cl
C0159982|ICD9CM|HT|836.6|Other dislocation of knee, open
C0159982|ICD9CM|PT|836.69|Other dislocation of knee, open
C0159982|ICD9CM|AB|836.69|Dislocat knee NEC-open
C0159984|ICD9CM|PT|836.61|Anterior dislocation of tibia, proximal end, open
C0159984|ICD9CM|AB|836.61|Ant disl prox tibia-open
C0159985|ICD9CM|PT|836.62|Posterior dislocation of tibia, proximal end, open
C0159985|ICD9CM|AB|836.62|Post disl prox tibia-opn
C0159986|ICD9CM|PT|836.63|Medial dislocation of tibia, proximal end, open
C0159986|ICD9CM|AB|836.63|Med disl prox tibia-open
C0159987|ICD9CM|PT|836.64|Lateral dislocation of tibia, proximal end, open
C0159987|ICD9CM|AB|836.64|Lat disl prox tibia-open
C0159990|ICD9CM|PT|837.1|Open dislocation of ankle
C0159990|ICD9CM|AB|837.1|Dislocation ankle-open
C0159993|ICD9CM|PT|838.01|Closed dislocation of tarsal (bone), joint unspecified
C0159993|ICD9CM|AB|838.01|Disloc tarsal NOS-closed
C0159994|ICD9CM|PT|838.02|Closed dislocation of midtarsal (joint)
C0159994|ICD9CM|AB|838.02|Disloc midtarsal-closed
C0159995|ICD9CM|PT|838.03|Closed dislocation of tarsometatarsal (joint)
C0159995|ICD9CM|AB|838.03|Disloc tarsometatars-cl
C0159996|ICD9CM|PT|838.04|Closed dislocation of metatarsal (bone), joint unspecified
C0159996|ICD9CM|AB|838.04|Disloc metatarsal NOS-cl
C0159997|ICD9CM|PT|838.05|Closed dislocation of metatarsophalangeal (joint)
C0159997|ICD9CM|AB|838.05|Disl metatarsophalang-cl
C0159998|ICD9CM|PT|838.06|Closed dislocation of interphalangeal (joint), foot
C0159998|ICD9CM|AB|838.06|Disl interphalan foot-cl
C0159999|ICD9CM|PT|838.09|Closed dislocation of foot, other
C0159999|ICD9CM|AB|838.09|Dislocat foot NEC-closed
C0160001|ICD9CM|PT|838.11|Open dislocation of tarsal (bone), joint unspecified
C0160001|ICD9CM|AB|838.11|Disloc tarsal NOS-open
C0160004|ICD9CM|PT|838.14|Open dislocation of metatarsal (bone), joint unspecified
C0160004|ICD9CM|AB|838.14|Disl metatarsal NOS-open
C0160005|ICD9CM|PT|838.15|Open dislocation of metatarsophalangeal (joint)
C0160005|ICD9CM|AB|838.15|Disloc metatarsophal-opn
C0160006|ICD9CM|PT|838.16|Open dislocation of interphalangeal (joint), foot
C0160006|ICD9CM|AB|838.16|Dis interphalan foot-opn
C0160007|ICD9CM|PT|838.19|Open dislocation of foot, other
C0160007|ICD9CM|AB|838.19|Dislocat foot NEC-open
C0160008|ICD9CM|HT|839.0|Closed dislocation, cervical vertebra
C0160008|ICD9CM|PT|839.00|Closed dislocation, cervical vertebra, unspecified
C0160008|ICD9CM|AB|839.00|Disloc cerv vert NOS-cl
C0160009|ICD9CM|PT|839.01|Closed dislocation, first cervical vertebra
C0160009|ICD9CM|AB|839.01|Disloc 1st cerv vert-cl
C0160010|ICD9CM|PT|839.02|Closed dislocation, second cervical vertebra
C0160010|ICD9CM|AB|839.02|Disloc 2nd cerv vert-cl
C0160011|ICD9CM|PT|839.03|Closed dislocation, third cervical vertebra
C0160011|ICD9CM|AB|839.03|Disloc 3rd cerv vert-cl
C0160012|ICD9CM|PT|839.04|Closed dislocation, fourth cervical vertebra
C0160012|ICD9CM|AB|839.04|Disloc 4th cerv vert-cl
C0160013|ICD9CM|PT|839.05|Closed dislocation, fifth cervical vertebra
C0160013|ICD9CM|AB|839.05|Disloc 5th cerv vert-cl
C0160014|ICD9CM|PT|839.06|Closed dislocation, sixth cervical vertebra
C0160014|ICD9CM|AB|839.06|Disloc 6th cerv vert-cl
C0160015|ICD9CM|PT|839.07|Closed dislocation, seventh cervical vertebra
C0160015|ICD9CM|AB|839.07|Disloc 7th cerv vert-cl
C0160016|ICD9CM|PT|839.08|Closed dislocation, multiple cervical vertebrae
C0160016|ICD9CM|AB|839.08|Disloc mult cerv vert-cl
C0160017|ICD9CM|HT|839.1|Open dislocation, cervical vertebra
C0160017|ICD9CM|PT|839.10|Open dislocation, cervical vertebra, unspecified
C0160017|ICD9CM|AB|839.10|Disloc cerv vert NOS-opn
C0160018|ICD9CM|PT|839.11|Open dislocation, first cervical vertebra
C0160018|ICD9CM|AB|839.11|Disloc lst cerv vert-opn
C0160019|ICD9CM|PT|839.12|Open dislocation, second cervical vertebra
C0160019|ICD9CM|AB|839.12|Disloc 2nd cerv vert-opn
C0160020|ICD9CM|PT|839.13|Open dislocation, third cervical vertebra
C0160020|ICD9CM|AB|839.13|Disloc 3rd cerv vert-opn
C0160021|ICD9CM|PT|839.14|Open dislocation, fourth cervical vertebra
C0160021|ICD9CM|AB|839.14|Disloc 4th cerv vert-opn
C0160022|ICD9CM|PT|839.15|Open dislocation, fifth cervical vertebra
C0160022|ICD9CM|AB|839.15|Disloc 5th cerv vert-opn
C0160023|ICD9CM|PT|839.16|Open dislocation, sixth cervical vertebra
C0160023|ICD9CM|AB|839.16|Disloc 6th cerv vert-opn
C0160024|ICD9CM|PT|839.17|Open dislocation, seventh cervical vertebra
C0160024|ICD9CM|AB|839.17|Disloc 7th cerv vert-opn
C0160025|ICD9CM|PT|839.18|Open dislocation, multiple cervical vertebrae
C0160025|ICD9CM|AB|839.18|Disloc mlt cerv vert-opn
C0160026|ICD9CM|HT|839.2|Closed dislocation, thoracic and lumbar vertebra
C0160027|ICD9CM|PT|839.20|Closed dislocation, lumbar vertebra
C0160027|ICD9CM|AB|839.20|Dislocat lumbar vert-cl
C0160028|ICD9CM|PT|839.21|Closed dislocation, thoracic vertebra
C0160028|ICD9CM|AB|839.21|Disloc thoracic vert-cl
C0160029|ICD9CM|HT|839.3|Open dislocation, thoracic and lumbar vertebra
C0160030|ICD9CM|PT|839.30|Open dislocation, lumbar vertebra
C0160030|ICD9CM|AB|839.30|Dislocat lumbar vert-opn
C0160031|ICD9CM|PT|839.31|Open dislocation, thoracic vertebra
C0160031|ICD9CM|AB|839.31|Disloc thoracic vert-opn
C0160032|ICD9CM|PT|839.49|Closed dislocation, vertebra, other
C0160032|ICD9CM|HT|839.4|Closed dislocation, other vertebra
C0160032|ICD9CM|AB|839.49|Dislocat vertebra NEC-cl
C0160033|ICD9CM|PT|839.40|Closed dislocation, vertebra, unspecified site
C0160033|ICD9CM|AB|839.40|Dislocat vertebra NOS-cl
C0160034|ICD9CM|PT|839.41|Closed dislocation, coccyx
C0160034|ICD9CM|AB|839.41|Dislocat coccyx-closed
C0160035|ICD9CM|PT|839.42|Closed dislocation, sacrum
C0160035|ICD9CM|AB|839.42|Dislocat sacrum-closed
C0160036|ICD9CM|HT|839.5|Open dislocation, other vertebra
C0160036|ICD9CM|PT|839.59|Open dislocation, vertebra,other
C0160036|ICD9CM|AB|839.59|Disloc vertebra NEC-open
C0160037|ICD9CM|PT|839.50|Open dislocation, vertebra, unspecified site
C0160037|ICD9CM|AB|839.50|Disloc vertebra NOS-open
C0160038|ICD9CM|PT|839.51|Open dislocation, coccyx
C0160038|ICD9CM|AB|839.51|Dislocat coccyx-open
C0160039|ICD9CM|PT|839.52|Open dislocation, sacrum
C0160039|ICD9CM|AB|839.52|Dislocat sacrum-open
C0160040|ICD9CM|HT|839.6|Closed dislocation, other location
C0160040|ICD9CM|PT|839.69|Closed dislocation, other location
C0160040|ICD9CM|AB|839.69|Dislocat site NEC-closed
C0160041|ICD9CM|PT|839.61|Closed dislocation, sternum
C0160041|ICD9CM|AB|839.61|Dislocat sternum-closed
C0160042|ICD9CM|HT|839.7|Open dislocation, other location
C0160042|ICD9CM|PT|839.79|Open dislocation, other location
C0160042|ICD9CM|AB|839.79|Dislocat site NEC-open
C0160043|ICD9CM|PT|839.71|Open dislocation, sternum
C0160043|ICD9CM|AB|839.71|Dislocation sternum-open
C0160044|ICD9CM|PT|839.9|Open dislocation, multiple and ill-defined sites
C0160044|ICD9CM|AB|839.9|Dislocation NEC-open
C0160045|ICD9CM|HT|840|Sprains and strains of shoulder and upper arm
C0160047|ICD9CM|PT|840.1|Coracoclavicular (ligament) sprain
C0160047|ICD9CM|AB|840.1|Sprain coracoclavicular
C0160051|ICD9CM|PT|840.5|Subscapularis (muscle) sprain
C0160051|ICD9CM|AB|840.5|Sprain subscapularis
C0160053|ICD9CM|PT|840.8|Sprains and strains of other specified sites of shoulder and upper arm
C0160053|ICD9CM|AB|840.8|Sprain shoulder/arm NEC
C0160054|ICD9CM|PT|840.9|Sprains and strains of unspecified site of shoulder and upper arm
C0160054|ICD9CM|AB|840.9|Sprain shoulder/arm NOS
C0160055|ICD9CM|HT|841|Sprains and strains of elbow and forearm
C0160056|ICD9CM|PT|841.0|Radial collateral ligament sprain
C0160056|ICD9CM|AB|841.0|Sprain radial collat lig
C0160058|ICD9CM|PT|841.2|Radiohumeral (joint) sprain
C0160058|ICD9CM|AB|841.2|Sprain radiohumeral
C0160060|ICD9CM|PT|841.8|Sprains and strains of other specified sites of elbow and forearm
C0160060|ICD9CM|AB|841.8|Sprain elbow/forearm NEC
C0160061|ICD9CM|PT|841.9|Sprains and strains of unspecified site of elbow and forearm
C0160061|ICD9CM|AB|841.9|Sprain elbow/forearm NOS
C0160062|ICD9CM|HT|842|Sprains and strains of wrist and hand
C0160063|ICD9CM|HT|842.0|Wrist sprain
C0160063|ICD9CM|AB|842.00|Sprain of wrist NOS
C0160063|ICD9CM|PT|842.00|Sprain of wrist, unspecified site
C0160067|ICD9CM|PT|842.09|Other sprains and strains of wrist
C0160067|ICD9CM|AB|842.09|Sprain of wrist NEC
C0160068|ICD9CM|HT|842.1|Hand sprain
C0160068|ICD9CM|AB|842.10|Sprain of hand NOS
C0160068|ICD9CM|PT|842.10|Sprain of hand, unspecified site
C0160070|ICD9CM|PT|842.11|Sprain of carpometacarpal (joint) of hand
C0160070|ICD9CM|AB|842.11|Sprain carpometacarpal
C0160071|ICD9CM|PT|842.12|Sprain of metacarpophalangeal (joint) of hand
C0160071|ICD9CM|AB|842.12|Sprain metacarpophalang
C0160072|ICD9CM|PT|842.13|Sprain of interphalangeal (joint) of hand
C0160072|ICD9CM|AB|842.13|Sprain interphalangeal
C0160073|ICD9CM|PT|842.19|Other sprains and strains of hand
C0160073|ICD9CM|AB|842.19|Sprain of hand NEC
C0160074|ICD9CM|HT|843|Sprains and strains of hip and thigh
C0160075|ICD9CM|PT|843.0|Iliofemoral (ligament) sprain
C0160075|ICD9CM|AB|843.0|Sprain iliofemoral
C0160077|ICD9CM|PT|843.8|Sprains and strains of other specified sites of hip and thigh
C0160077|ICD9CM|AB|843.8|Sprain hip & thigh NEC
C0160078|ICD9CM|PT|843.9|Sprains and strains of unspecified site of hip and thigh
C0160078|ICD9CM|AB|843.9|Sprain hip & thigh NOS
C0160079|ICD9CM|HT|844|Sprains and strains of knee and leg
C0160080|ICD9CM|PT|844.0|Sprain of lateral collateral ligament of knee
C0160080|ICD9CM|AB|844.0|Sprain lateral coll lig
C0160081|ICD9CM|PT|844.1|Sprain of medial collateral ligament of knee
C0160081|ICD9CM|AB|844.1|Sprain medial collat lig
C0160082|ICD9CM|PT|844.2|Sprain of cruciate ligament of knee
C0160082|ICD9CM|AB|844.2|Sprain cruciate lig knee
C0160084|ICD9CM|PT|844.8|Sprains and strains of other specified sites of knee and leg
C0160084|ICD9CM|AB|844.8|Sprain of knee & leg NEC
C0160085|ICD9CM|PT|844.9|Sprains and strains of unspecified site of knee and leg
C0160085|ICD9CM|AB|844.9|Sprain of knee & leg NOS
C0160086|ICD9CM|HT|845|Sprains and strains of ankle and foot
C0160087|ICD9CM|HT|845.0|Ankle sprain
C0160087|ICD9CM|AB|845.00|Sprain of ankle NOS
C0160087|ICD9CM|PT|845.00|Sprain of ankle, unspecified site
C0160089|ICD9CM|PT|845.01|Sprain of deltoid (ligament), ankle
C0160089|ICD9CM|AB|845.01|Sprain of ankle deltoid
C0160090|ICD9CM|PT|845.02|Sprain of calcaneofibular (ligament) of ankle
C0160090|ICD9CM|AB|845.02|Sprain calcaneofibular
C0160091|ICD9CM|PT|845.03|Sprain of tibiofibular (ligament), distal of ankle
C0160091|ICD9CM|AB|845.03|Sprain distal tibiofibul
C0160092|ICD9CM|PT|845.09|Other sprains and strains of ankle
C0160092|ICD9CM|AB|845.09|Sprain of ankle NEC
C0160093|ICD9CM|HT|845.1|Foot sprain
C0160094|ICD9CM|PT|845.10|Sprain of foot, unspecified site
C0160094|ICD9CM|AB|845.10|Sprain of foot NOS
C0160096|ICD9CM|AB|845.12|Sprain metatarsophalang
C0160096|ICD9CM|PT|845.12|Sprain of metatarsophalangeal (joint) of foot
C0160097|ICD9CM|PT|845.13|Sprain of interphalangeal (joint), toe
C0160097|ICD9CM|AB|845.13|Sprain interphalang toe
C0160098|ICD9CM|PT|845.19|Other sprain of foot
C0160098|ICD9CM|AB|845.19|Sprain of foot NEC
C0160099|ICD9CM|HT|846|Sprains and strains of sacroiliac region
C0160102|ICD9CM|PT|846.2|Sprain of sacrospinatus (ligament)
C0160102|ICD9CM|AB|846.2|Sprain sacrospinatus
C0160103|ICD9CM|PT|846.3|Sprain of sacrotuberous (ligament)
C0160103|ICD9CM|AB|846.3|Sprain sacrotuberous
C0160104|ICD9CM|PT|846.8|Sprain of other specified sites of sacroiliac region
C0160104|ICD9CM|AB|846.8|Sprain sacroiliac NEC
C0160105|ICD9CM|PT|846.9|Sprain of unspecified site of sacroiliac region
C0160105|ICD9CM|AB|846.9|Sprain sacroiliac NOS
C0160106|ICD9CM|HT|847|Sprains and strains of other and unspecified parts of back
C0160107|ICD9CM|PT|847.1|Sprain of thoracic
C0160107|ICD9CM|AB|847.1|Sprain thoracic region
C0160108|ICD9CM|PT|847.2|Sprain of lumbar
C0160108|ICD9CM|AB|847.2|Sprain lumbar region
C0160109|ICD9CM|AB|847.3|Sprain of sacrum
C0160109|ICD9CM|PT|847.3|Sprain of sacrum
C0160110|ICD9CM|AB|847.4|Sprain of coccyx
C0160110|ICD9CM|PT|847.4|Sprain of coccyx
C0160111|ICD9CM|PT|847.9|Sprain of unspecified site of back
C0160111|ICD9CM|AB|847.9|Sprain of back NOS
C0160112|ICD9CM|PT|848.0|Sprain of septal cartilage of nose
C0160112|ICD9CM|AB|848.0|Sprain of nasal septum
C0160113|ICD9CM|AB|848.1|Sprain of jaw
C0160113|ICD9CM|PT|848.1|Sprain of jaw
C0160114|ICD9CM|AB|848.2|Sprain of thyroid region
C0160114|ICD9CM|PT|848.2|Sprain of thyroid region
C0160115|ICD9CM|AB|848.3|Sprain of ribs
C0160115|ICD9CM|PT|848.3|Sprain of ribs
C0160118|ICD9CM|PT|848.42|Sprain of chondrosternal (joint)
C0160118|ICD9CM|AB|848.42|Sprain chondrosternal
C0160119|ICD9CM|PT|848.49|Sprain of sternum, other
C0160119|ICD9CM|AB|848.49|Sprain of sternum NEC
C0160121|ICD9CM|PT|850.0|Concussion with no loss of consciousness
C0160121|ICD9CM|AB|850.0|Concussion w/o coma
C0160122|ICD9CM|HT|850.1|Concussion with brief loss of consciousness
C0160123|ICD9CM|PT|850.2|Concussion with moderate loss of consciousness
C0160123|ICD9CM|AB|850.2|Concussion-moderate coma
C0160124|ICD9CM|PT|850.3|Concussion with prolonged loss of consciousness and return to pre-existing conscious level
C0160124|ICD9CM|AB|850.3|Concussion-prolong coma
C0160125|ICD9CM|PT|850.4|Concussion with prolonged loss of consciousness, without return to pre-existing conscious level
C0160125|ICD9CM|AB|850.4|Concussion-deep coma
C0160126|ICD9CM|PT|850.5|Concussion with loss of consciousness of unspecified duration
C0160126|ICD9CM|AB|850.5|Concussion w coma NOS
C0160127|ICD9CM|HT|851|Cerebral laceration and contusion
C0160128|ICD9CM|HT|851.0|Cortex (cerebral) contusion without mention of open intracranial wound
C0160131|ICD9CM|PT|851.02|Cortex (cerebral) contusion without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160131|ICD9CM|AB|851.02|Cortex contus-brief coma
C0160133|ICD9CM|PT|851.04|Cortex (cerebral) contusion without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160133|ICD9CM|AB|851.04|Cortx contus-prolng coma
C0160134|ICD9CM|PT|851.05|Cortex (cerebral) contusion without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160134|ICD9CM|AB|851.05|Cortex contus-deep coma
C0160137|ICD9CM|HT|851.1|Cortex (cerebral) contusion with open intracranial wound
C0160138|ICD9CM|PT|851.10|Cortex (cerebral) contusion with open intracranial wound, unspecified state of consciousness
C0160138|ICD9CM|AB|851.10|Cortex contusion/opn wnd
C0160140|ICD9CM|PT|851.12|Cortex (cerebral) contusion with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160140|ICD9CM|AB|851.12|Opn cort contus-brf coma
C0160141|ICD9CM|PT|851.13|Cortex (cerebral) contusion with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160141|ICD9CM|AB|851.13|Opn cort contus-mod coma
C0160142|ICD9CM|PT|851.14|Cortex (cerebral) contusion with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160142|ICD9CM|AB|851.14|Opn cort contu-prol coma
C0160143|ICD9CM|PT|851.15|Cortex (cerebral) contusion with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160143|ICD9CM|AB|851.15|Opn cort contu-deep coma
C0160149|ICD9CM|PT|851.22|Cortex (cerebral) laceration without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160149|ICD9CM|AB|851.22|Cortex lacera-brief coma
C0160150|ICD9CM|PT|851.23|Cortex (cerebral) laceration without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160150|ICD9CM|AB|851.23|Cortex lacerat-mod coma
C0160151|ICD9CM|PT|851.24|Cortex (cerebral) laceration without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160151|ICD9CM|AB|851.24|Cortex lacerat-prol coma
C0160152|ICD9CM|PT|851.25|Cortex (cerebral) laceration without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160152|ICD9CM|AB|851.25|Cortex lacerat-deep coma
C0160158|ICD9CM|PT|851.32|Cortex (cerebral) laceration with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160158|ICD9CM|AB|851.32|Opn cortx lac-brief coma
C0160159|ICD9CM|PT|851.33|Cortex (cerebral) laceration with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160159|ICD9CM|AB|851.33|Opn cortx lacer-mod coma
C0160160|ICD9CM|PT|851.34|Cortex (cerebral) laceration with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160160|ICD9CM|AB|851.34|Opn cortx lac-proln coma
C0160164|ICD9CM|HT|851.4|Cerebellar or brain stem contusion without mention of open intracranial wound
C0160165|ICD9CM|PT|851.40|Cerebellar or brain stem contusion without mention of open intracranial wound, unspecified state of consciousness
C0160165|ICD9CM|AB|851.40|Cerebel/brain stm contus
C0160166|ICD9CM|PT|851.41|Cerebellar or brain stem contusion without mention of open intracranial wound, with no loss of consciousness
C0160166|ICD9CM|AB|851.41|Cerebell contus w/o coma
C0160167|ICD9CM|PT|851.42|Cerebellar or brain stem contusion without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160167|ICD9CM|AB|851.42|Cerebell contus-brf coma
C0160168|ICD9CM|PT|851.43|Cerebellar or brain stem contusion without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160168|ICD9CM|AB|851.43|Cerebell contus-mod coma
C0160169|ICD9CM|PT|851.44|Cerebellar or brain stem contusion without mention of open intracranial wound, with prolonged [more than 24 hours] loss consciousness and return to pre-existing conscious level
C0160169|ICD9CM|AB|851.44|Cerebel contus-prol coma
C0160170|ICD9CM|PT|851.45|Cerebellar or brain stem contusion without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160170|ICD9CM|AB|851.45|Cerebel contus-deep coma
C0160171|ICD9CM|PT|851.46|Cerebellar or brain stem contusion without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0160171|ICD9CM|AB|851.46|Cerebell contus-coma NOS
C0160173|ICD9CM|HT|851.5|Cerebellar or brain stem contusion with open intracranial wound
C0160174|ICD9CM|PT|851.50|Cerebellar or brain stem contusion with open intracranial wound, unspecified state of consciousness
C0160174|ICD9CM|AB|851.50|Cerebel contus w opn wnd
C0160175|ICD9CM|PT|851.51|Cerebellar or brain stem contusion with open intracranial wound, with no loss of consciousness
C0160175|ICD9CM|AB|851.51|Opn cerebe cont w/o coma
C0160176|ICD9CM|PT|851.52|Cerebellar or brain stem contusion with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160176|ICD9CM|AB|851.52|Opn cerebe cont-brf coma
C0160177|ICD9CM|PT|851.53|Cerebellar or brain stem contusion with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160177|ICD9CM|AB|851.53|Opn cerebe cont-mod coma
C0160178|ICD9CM|PT|851.54|Cerebellar or brain stem contusion with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160178|ICD9CM|AB|851.54|Opn cerebe cont-prol com
C0160179|ICD9CM|PT|851.55|Cerebellar or brain stem contusion with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160179|ICD9CM|AB|851.55|Opn cerebe cont-deep com
C0160180|ICD9CM|PT|851.56|Cerebellar or brain stem contusion with open intracranial wound, with loss of consciousness of unspecified duration
C0160180|ICD9CM|AB|851.56|Opn cerebe cont-coma NOS
C0160182|ICD9CM|HT|851.6|Cerebellar or brain stem laceration without mention of open intracranial wound
C0160183|ICD9CM|PT|851.60|Cerebellar or brain stem laceration without mention of open intracranial wound, unspecified state of consciousness
C0160183|ICD9CM|AB|851.60|Cerebel/brain stem lacer
C0160184|ICD9CM|PT|851.61|Cerebellar or brain stem laceration without mention of open intracranial wound, with no loss of consciousness
C0160184|ICD9CM|AB|851.61|Cerebel lacerat w/o coma
C0160185|ICD9CM|PT|851.62|Cerebellar or brain stem laceration without mention of open intracranial wound, with brief [less than 1 hour] loss of consciousness
C0160185|ICD9CM|AB|851.62|Cerebel lacer-brief coma
C0160186|ICD9CM|PT|851.63|Cerebellar or brain stem laceration without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160186|ICD9CM|AB|851.63|Cerebel lacerat-mod coma
C0160187|ICD9CM|PT|851.64|Cerebellar or brain stem laceration without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160187|ICD9CM|AB|851.64|Cerebel lacer-proln coma
C0160188|ICD9CM|PT|851.65|Cerebellar or brain stem laceration without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160188|ICD9CM|AB|851.65|Cerebell lacer-deep coma
C0160189|ICD9CM|PT|851.66|Cerebellar or brain stem laceration without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0160189|ICD9CM|AB|851.66|Cerebel lacerat-coma NOS
C0160191|ICD9CM|HT|851.7|Cerebellar or brain stem laceration with open intracranial wound
C0160192|ICD9CM|PT|851.70|Cerebellar or brain stem laceration with open intracranial wound, unspecified state of consciousness
C0160192|ICD9CM|AB|851.70|Cerebel lacer w open wnd
C0160193|ICD9CM|PT|851.71|Cerebellar or brain stem laceration with open intracranial wound, with no loss of consciousness
C0160193|ICD9CM|AB|851.71|Opn cerebel lac w/o coma
C0160194|ICD9CM|PT|851.72|Cerebellar or brain stem laceration with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160194|ICD9CM|AB|851.72|Opn cerebel lac-brf coma
C0160195|ICD9CM|PT|851.73|Cerebellar or brain stem laceration with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160195|ICD9CM|AB|851.73|Opn cerebel lac-mod coma
C0160196|ICD9CM|PT|851.74|Cerebellar or brain stem laceration with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160196|ICD9CM|AB|851.74|Opn cerebe lac-prol coma
C0160197|ICD9CM|PT|851.75|Cerebellar or brain stem laceration with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160197|ICD9CM|AB|851.75|Opn cerebe lac-deep coma
C0160198|ICD9CM|PT|851.76|Cerebellar or brain stem laceration with open intracranial wound, with loss of consciousness of unspecified duration
C0160198|ICD9CM|AB|851.76|Opn cerebel lac-coma NOS
C0160200|ICD9CM|HT|851.8|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound
C0160201|ICD9CM|PT|851.80|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, unspecified state of consciousness
C0160201|ICD9CM|AB|851.80|Brain laceration NEC
C0160202|ICD9CM|PT|851.81|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with no loss of consciousness
C0160202|ICD9CM|AB|851.81|Brain lacer NEC w/o coma
C0160203|ICD9CM|PT|851.82|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160203|ICD9CM|AB|851.82|Brain lac NEC-brief coma
C0160204|ICD9CM|PT|851.83|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160204|ICD9CM|AB|851.83|Brain lacer NEC-mod coma
C0160205|ICD9CM|PT|851.84|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre- existing conscious level
C0160205|ICD9CM|AB|851.84|Brain lac NEC-proln coma
C0160206|ICD9CM|PT|851.85|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160206|ICD9CM|AB|851.85|Brain lac NEC-deep coma
C0160207|ICD9CM|PT|851.86|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0160207|ICD9CM|AB|851.86|Brain lacer NEC-coma NOS
C0160209|ICD9CM|HT|851.9|Other and unspecified cerebral laceration and contusion, with open intracranial wound
C0160210|ICD9CM|PT|851.90|Other and unspecified cerebral laceration and contusion, with open intracranial wound, unspecified state of consciousness
C0160210|ICD9CM|AB|851.90|Brain lac NEC w open wnd
C0160211|ICD9CM|PT|851.91|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with no loss of consciousness
C0160211|ICD9CM|AB|851.91|Opn brain lacer w/o coma
C0160212|ICD9CM|PT|851.92|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160212|ICD9CM|AB|851.92|Opn brain lac-brief coma
C0160213|ICD9CM|PT|851.93|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160213|ICD9CM|AB|851.93|Opn brain lacer-mod coma
C0160214|ICD9CM|PT|851.94|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160214|ICD9CM|AB|851.94|Opn brain lac-proln coma
C0160215|ICD9CM|PT|851.95|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160215|ICD9CM|AB|851.95|Open brain lac-deep coma
C0160216|ICD9CM|PT|851.96|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with loss of consciousness of unspecified duration
C0160216|ICD9CM|AB|851.96|Opn brain lacer-coma NOS
C0160218|ICD9CM|HT|852|Subarachnoid, subdural, and extradural hemorrhage, following injury
C0160219|ICD9CM|HT|852.0|Subarachnoid hemorrhage following injury without mention of open intracranial wound
C0160220|ICD9CM|PT|852.00|Subarachnoid hemorrhage following injury without mention of open intracranial wound, unspecified state of consciousness
C0160220|ICD9CM|AB|852.00|Traum subarachnoid hem
C0160221|ICD9CM|PT|852.01|Subarachnoid hemorrhage following injury without mention of open intracranial wound, with no loss of consciousness
C0160221|ICD9CM|AB|852.01|Subarachnoid hem-no coma
C0160222|ICD9CM|PT|852.02|Subarachnoid hemorrhage following injury without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160222|ICD9CM|AB|852.02|Subarach hem-brief coma
C0160223|ICD9CM|PT|852.03|Subarachnoid hemorrhage following injury without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160223|ICD9CM|AB|852.03|Subarach hem-mod coma
C0160224|ICD9CM|PT|852.04|Subarachnoid hemorrhage following injury without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160224|ICD9CM|AB|852.04|Subarach hem-prolng coma
C0160225|ICD9CM|PT|852.05|Subarachnoid hemorrhage following injury without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160225|ICD9CM|AB|852.05|Subarach hem-deep coma
C0160226|ICD9CM|PT|852.06|Subarachnoid hemorrhage following injury without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0160226|ICD9CM|AB|852.06|Subarach hem-coma NOS
C0160227|ICD9CM|PT|852.09|Subarachnoid hemorrhage following injury without mention of open intracranial wound, with concussion, unspecified
C0160227|ICD9CM|AB|852.09|Subarach hem-concussion
C0160228|ICD9CM|HT|852.1|Subarachnoid hemorrhage following injury with open intracranial wound
C0160229|ICD9CM|PT|852.10|Subarachnoid hemorrhage following injury with open intracranial wound, unspecified state of consciousness
C0160229|ICD9CM|AB|852.10|Subarach hem w opn wound
C0160230|ICD9CM|PT|852.11|Subarachnoid hemorrhage following injury with open intracranial wound, with no loss of consciousness
C0160230|ICD9CM|AB|852.11|Opn subarach hem-no coma
C0160231|ICD9CM|PT|852.12|Subarachnoid hemorrhage following injury with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160231|ICD9CM|AB|852.12|Op subarach hem-brf coma
C0160232|ICD9CM|PT|852.13|Subarachnoid hemorrhage following injury with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160232|ICD9CM|AB|852.13|Op subarach hem-mod coma
C0160233|ICD9CM|PT|852.14|Subarachnoid hemorrhage following injury with open intracranial wound, with prolonged [more than 24 hours) loss of consciousness and return to pre-existing conscious level
C0160233|ICD9CM|AB|852.14|Op subarach hem-prol com
C0160234|ICD9CM|PT|852.15|Subarachnoid hemorrhage following injury with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160234|ICD9CM|AB|852.15|Op subarach hem-deep com
C0160235|ICD9CM|PT|852.16|Subarachnoid hemorrhage following injury with open intracranial wound, with loss of consciousness of unspecified duration
C0160235|ICD9CM|AB|852.16|Op subarach hem-coma NOS
C0160237|ICD9CM|HT|852.2|Subdural hemorrhage following injury without mention of open intracranial wound
C0160238|ICD9CM|PT|852.20|Subdural hemorrhage following injury without mention of open intracranial wound, unspecified state of consciousness
C0160238|ICD9CM|AB|852.20|Traumatic subdural hem
C0160239|ICD9CM|PT|852.21|Subdural hemorrhage following injury without mention of open intracranial wound, with no loss of consciousness
C0160239|ICD9CM|AB|852.21|Subdural hem w/o coma
C0160240|ICD9CM|PT|852.22|Subdural hemorrhage following injury without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160240|ICD9CM|AB|852.22|Subdural hem-brief coma
C0160241|ICD9CM|PT|852.23|Subdural hemorrhage following injury without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160241|ICD9CM|AB|852.23|Subdural hemorr-mod coma
C0160242|ICD9CM|PT|852.24|Subdural hemorrhage following injury without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160242|ICD9CM|AB|852.24|Subdural hem-prolng coma
C0160243|ICD9CM|PT|852.25|Subdural hemorrhage following injury without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160243|ICD9CM|AB|852.25|Subdural hem-deep coma
C0160244|ICD9CM|PT|852.26|Subdural hemorrhage following injury without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0160244|ICD9CM|AB|852.26|Subdural hemorr-coma NOS
C0160245|ICD9CM|PT|852.29|Subdural hemorrhage following injury without mention of open intracranial wound, with concussion, unspecified
C0160245|ICD9CM|AB|852.29|Subdural hem-concussion
C0160246|ICD9CM|HT|852.3|Subdural hemorrhage following injury, with open intracranial wound
C0160247|ICD9CM|PT|852.30|Subdural hemorrhage following injury with open intracranial wound, unspecified state of consciousness
C0160247|ICD9CM|AB|852.30|Subdural hem w opn wound
C0160248|ICD9CM|PT|852.31|Subdural hemorrhage following injury with open intracranial wound, with no loss of consciousness
C0160248|ICD9CM|AB|852.31|Open subdur hem w/o coma
C0160249|ICD9CM|PT|852.32|Subdural hemorrhage following injury with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160249|ICD9CM|AB|852.32|Opn subdur hem-brf coma
C0160250|ICD9CM|PT|852.33|Subdural hemorrhage following injury with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160250|ICD9CM|AB|852.33|Opn subdur hem-mod coma
C0160251|ICD9CM|PT|852.34|Subdural hemorrhage following injury with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160251|ICD9CM|AB|852.34|Opn subdur hem-prol coma
C0160252|ICD9CM|PT|852.35|Subdural hemorrhage following injury with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160252|ICD9CM|AB|852.35|Opn subdur hem-deep coma
C0160253|ICD9CM|PT|852.36|Subdural hemorrhage following injury with open intracranial wound, with loss of consciousness of unspecified duration
C0160253|ICD9CM|AB|852.36|Opn subdur hem-coma NOS
C0160255|ICD9CM|HT|852.4|Extradural hemorrhage following injury without mention of open intracranial wound
C0160258|ICD9CM|PT|852.42|Extradural hemorrhage following injury without mention of open intracranial wound, with brief [less than 1 hour] loss of consciousness
C0160258|ICD9CM|AB|852.42|Extradur hem-brief coma
C0160259|ICD9CM|PT|852.43|Extradural hemorrhage following injury without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160259|ICD9CM|AB|852.43|Extradural hem-mod coma
C0160260|ICD9CM|PT|852.44|Extradural hemorrhage following injury without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160260|ICD9CM|AB|852.44|Extradur hem-proln coma
C0160263|ICD9CM|PT|852.49|Extradural hemorrhage following injury without mention of open intracranial wound, with concussion, unspecified
C0160263|ICD9CM|AB|852.49|Extadural hem-concuss
C0160264|ICD9CM|HT|852.5|Extradural hemorrhage following injury with open intracranial wound
C0160265|ICD9CM|PT|852.50|Extradural hemorrhage following injury with open intracranial wound, unspecified state of consciousness
C0160265|ICD9CM|AB|852.50|Extradural hem w opn wnd
C0160266|ICD9CM|PT|852.51|Extradural hemorrhage following injury with open intracranial wound, with no loss of consciousness
C0160266|ICD9CM|AB|852.51|Extradural hemor-no coma
C0160267|ICD9CM|PT|852.52|Extradural hemorrhage following injury with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160267|ICD9CM|AB|852.52|Extradur hem-brief coma
C0160268|ICD9CM|PT|852.53|Extradural hemorrhage following injury with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160268|ICD9CM|AB|852.53|Extradural hem-mod coma
C0160269|ICD9CM|PT|852.54|Extradural hemorrhage following injury with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160269|ICD9CM|AB|852.54|Extradur hem-proln coma
C0160270|ICD9CM|PT|852.55|Extradural hemorrhage following injury with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160270|ICD9CM|AB|852.55|Extradur hem-deep coma
C0160271|ICD9CM|PT|852.56|Extradural hemorrhage following injury with open intracranial wound, with loss of consciousness of unspecified duration
C0160271|ICD9CM|AB|852.56|Extradural hem-coma NOS
C0160273|ICD9CM|HT|853|Other and unspecified intracranial hemorrhage following injury
C0160274|ICD9CM|HT|853.0|Other and unspecified intracranial hemorrhage following injury, without mention of open intracranial wound
C0160275|ICD9CM|PT|853.00|Other and unspecified intracranial hemorrhage following injury without mention of open intracranial wound, unspecified state of consciousness
C0160275|ICD9CM|AB|853.00|Traumatic brain hem NEC
C0160276|ICD9CM|PT|853.01|Other and unspecified intracranial hemorrhage following injury without mention of open intracranial wound, with no loss of consciousness
C0160276|ICD9CM|AB|853.01|Brain hem NEC w/o coma
C0160277|ICD9CM|PT|853.02|Other and unspecified intracranial hemorrhage following injury without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160277|ICD9CM|AB|853.02|Brain hem NEC-brief coma
C0160278|ICD9CM|PT|853.03|Other and unspecified intracranial hemorrhage following injury without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160278|ICD9CM|AB|853.03|Brain hem NEC-mod coma
C0160279|ICD9CM|PT|853.04|Other and unspecified intracranial hemorrhage following injury without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre- existing conscious level
C0160279|ICD9CM|AB|853.04|Brain hem NEC-proln coma
C0160280|ICD9CM|PT|853.05|Other and unspecified intracranial hemorrhage following injury without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160280|ICD9CM|AB|853.05|Brain hem NEC-deep coma
C0160281|ICD9CM|PT|853.06|Other and unspecified intracranial hemorrhage following injury without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0160281|ICD9CM|AB|853.06|Brain hem NEC-coma NOS
C0160283|ICD9CM|HT|853.1|Other and unspecified intracranial hemorrhage following injury with open intracranial wound
C0160284|ICD9CM|PT|853.10|Other and unspecified intracranial hemorrhage following injury with open intracranial wound, unspecified state of consciousness
C0160284|ICD9CM|AB|853.10|Brain hem NEC w opn wnd
C0160285|ICD9CM|PT|853.11|Other and unspecified intracranial hemorrhage following injury with open intracranial wound, with no loss of consciousness
C0160285|ICD9CM|AB|853.11|Brain hem opn w/o coma
C0160286|ICD9CM|PT|853.12|Other and unspecified intracranial hemorrhage following injury with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160286|ICD9CM|AB|853.12|Brain hem opn-brf coma
C0160287|ICD9CM|PT|853.13|Other and unspecified intracranial hemorrhage following injury with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160287|ICD9CM|AB|853.13|Brain hem open-mod coma
C0160288|ICD9CM|PT|853.14|Other and unspecified intracranial hemorrhage following injury with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160288|ICD9CM|AB|853.14|Brain hem opn-proln coma
C0160289|ICD9CM|PT|853.15|Other and unspecified intracranial hemorrhage following injury with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160289|ICD9CM|AB|853.15|Brain hem open-deep coma
C0160290|ICD9CM|PT|853.16|Other and unspecified intracranial hemorrhage following injury with open intracranial wound, with loss of consciousness of unspecified duration
C0160290|ICD9CM|AB|853.16|Brain hem open-coma NOS
C0160292|ICD9CM|HT|854|Intracranial injury of other and unspecified nature
C0160293|ICD9CM|PT|854.01|Intracranial injury of other and unspecified nature without mention of open intracranial wound, with no loss of consciousness
C0160293|ICD9CM|AB|854.01|Brain injury NEC-no coma
C0160294|ICD9CM|PT|854.02|Intracranial injury of other and unspecified nature without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160294|ICD9CM|AB|854.02|Brain inj NEC-brief coma
C0160295|ICD9CM|PT|854.03|Intracranial injury of other and unspecified nature without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160295|ICD9CM|AB|854.03|Brain inj NEC-mod coma
C0160296|ICD9CM|PT|854.04|Intracranial injury of other and unspecified nature without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160296|ICD9CM|AB|854.04|Brain inj NEC-proln coma
C0160297|ICD9CM|PT|854.05|Intracranial injury of other and unspecified nature without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160297|ICD9CM|AB|854.05|Brain inj NEC-deep coma
C0160298|ICD9CM|PT|854.06|Intracranial injury of other and unspecified nature without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0160298|ICD9CM|AB|854.06|Brain inj NEC-coma NOS
C0160299|ICD9CM|PT|854.09|Intracranial injury of other and unspecified nature without mention of open intracranial wound, with concussion, unspecified
C0160299|ICD9CM|AB|854.09|Brain inj NEC-concussion
C0160300|ICD9CM|HT|854.1|Intracranial injury of other and unspecified nature with open intracranial wound
C0160301|ICD9CM|PT|854.10|Intracranial injury of other and unspecified nature with open intracranial wound, unspecified state of consciousness
C0160301|ICD9CM|AB|854.10|Brain injury w opn wnd
C0160302|ICD9CM|PT|854.11|Intracranial injury of other and unspecified nature with open intracranial wound, with no loss of consciousness
C0160302|ICD9CM|AB|854.11|Opn brain inj w/o coma
C0160303|ICD9CM|PT|854.12|Intracranial injury of other and unspecified nature with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160303|ICD9CM|AB|854.12|Opn brain inj-brief coma
C0160304|ICD9CM|PT|854.13|Intracranial injury of other and unspecified nature with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160304|ICD9CM|AB|854.13|Opn brain inj-mod coma
C0160305|ICD9CM|PT|854.14|Intracranial injury of other and unspecified nature with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160305|ICD9CM|AB|854.14|Opn brain inj-proln coma
C0160306|ICD9CM|PT|854.15|Intracranial injury of other and unspecified nature with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160306|ICD9CM|AB|854.15|Opn brain inj-deep coma
C0160307|ICD9CM|PT|854.16|Intracranial injury of other and unspecified nature with open intracranial wound, with loss of consciousness of unspecified duration
C0160307|ICD9CM|AB|854.16|Open brain inj-coma NOS
C0160308|ICD9CM|PT|854.19|Intracranial injury of other and unspecified nature with open intracranial wound, with concussion, unspecified
C0160308|ICD9CM|AB|854.19|Opn brain inj-concussion
C0160312|ICD9CM|PT|860.2|Traumatic hemothorax without mention of open wound into thorax
C0160312|ICD9CM|AB|860.2|Traum hemothorax-closed
C0160316|ICD9CM|HT|861|Injury to heart and lung
C0160318|ICD9CM|PT|861.00|Unspecified injury of heart without mention of open wound into thorax
C0160318|ICD9CM|HT|861.0|Heart injury, without mention of open wound into thorax
C0160318|ICD9CM|AB|861.00|Heart injury NOS-closed
C0160319|ICD9CM|PT|861.01|Contusion of heart without mention of open wound into thorax
C0160319|ICD9CM|AB|861.01|Heart contusion-closed
C0160320|ICD9CM|PT|861.02|Laceration of heart without penetration of heart chambers or without mention of open wound into thorax
C0160320|ICD9CM|AB|861.02|Heart laceration-closed
C0160321|ICD9CM|PT|861.03|Laceration of heart with penetration of heart chambers without mention of open wound into thorax
C0160321|ICD9CM|AB|861.03|Heart chamber lacerat-cl
C0160323|ICD9CM|HT|861.1|Heart injury, with open wound into thorax
C0160323|ICD9CM|PT|861.10|Unspecified injury of heart with open wound into thorax
C0160323|ICD9CM|AB|861.10|Heart injury NOS-open
C0160324|ICD9CM|PT|861.11|Contusion of heart with open wound into thorax
C0160324|ICD9CM|AB|861.11|Heart contusion-open
C0160325|ICD9CM|PT|861.12|Laceration of heart without penetration of heart chambers, with open wound into thorax
C0160325|ICD9CM|AB|861.12|Heart laceration-open
C0160326|ICD9CM|PT|861.13|Laceration of heart with penetration of heart chambers with open wound into thorax
C0160326|ICD9CM|AB|861.13|Heart chamber lacer-opn
C0160328|ICD9CM|HT|861.2|Lung injury, without mention of open wound into thorax
C0160328|ICD9CM|AB|861.20|Lung injury NOS-closed
C0160328|ICD9CM|PT|861.20|Unspecified injury of lung without mention of open wound into thorax
C0160329|ICD9CM|AB|861.21|Lung contusion-closed
C0160329|ICD9CM|PT|861.21|Contusion of lung without mention of open wound into thorax
C0160330|ICD9CM|AB|861.22|Lung laceration-closed
C0160330|ICD9CM|PT|861.22|Laceration of lung without mention of open wound into thorax
C0160332|ICD9CM|HT|861.3|Lung injury, with open wound into thorax
C0160332|ICD9CM|PT|861.30|Unspecified injury of lung with open wound into thorax
C0160332|ICD9CM|AB|861.30|Lung injury NOS-open
C0160333|ICD9CM|PT|861.31|Contusion of lung with open wound into thorax
C0160333|ICD9CM|AB|861.31|Lung contusion-open
C0160334|ICD9CM|PT|861.32|Laceration of lung with open wound into thorax
C0160334|ICD9CM|AB|861.32|Lung laceration-open
C0160335|ICD9CM|HT|862|Injury to other and unspecified intrathoracic organs
C0160336|ICD9CM|PT|862.1|Injury to diaphragm, with open wound into cavity
C0160336|ICD9CM|AB|862.1|Diaphragm injury-open
C0160337|ICD9CM|HT|862.2|Injury to other specified intrathoracic organs without mention of open wound into cavity
C0160337|ICD9CM|PT|862.29|Injury to other specified intrathoracic organs without mention of open wound into cavity
C0160337|ICD9CM|AB|862.29|Intrathoracic inj NEC-cl
C0160338|ICD9CM|AB|862.21|Bronchus injury-closed
C0160338|ICD9CM|PT|862.21|Injury to bronchus without mention of open wound into cavity
C0160340|ICD9CM|HT|862.3|Injury to other specified intrathoracic organs with open wound into cavity
C0160340|ICD9CM|PT|862.39|Injury to other specified intrathoracic organs with open wound into cavity
C0160340|ICD9CM|AB|862.39|Intrathorac inj NEC-open
C0160341|ICD9CM|PT|862.31|Injury to bronchus with open wound into cavity
C0160341|ICD9CM|AB|862.31|Bronchus injury-open
C0160342|ICD9CM|PT|862.32|Injury to esophagus with open wound into cavity
C0160342|ICD9CM|AB|862.32|Esophagus injury-open
C0160343|ICD9CM|PT|862.8|Injury to multiple and unspecified intrathoracic organs, without mention of open wound into cavity
C0160343|ICD9CM|AB|862.8|Intrathoracic inj NOS-cl
C0160345|ICD9CM|HT|863|Injury to gastrointestinal tract
C0160346|ICD9CM|PT|863.0|Injury to stomach, without mention of open wound into cavity
C0160346|ICD9CM|AB|863.0|Stomach injury-closed
C0160347|ICD9CM|PT|863.1|Injury to stomach, with open wound into cavity
C0160347|ICD9CM|AB|863.1|Stomach injury-open
C0160348|ICD9CM|HT|863.2|Injury to small intestine without mention of open wound into cavity
C0160349|ICD9CM|PT|863.20|Injury to small intestine, unspecified site, without open wound into cavity
C0160349|ICD9CM|AB|863.20|Small intest inj NOS-cl
C0160350|ICD9CM|PT|863.21|Injury to duodenum, without open wound into cavity
C0160350|ICD9CM|AB|863.21|Duodenum injury-closed
C0160351|ICD9CM|PT|863.29|Other injury to small intestine, without mention of open wound into cavity
C0160351|ICD9CM|AB|863.29|Small intest inj NEC-cl
C0160352|ICD9CM|HT|863.3|Injury to small intestine with open wound into cavity
C0160353|ICD9CM|PT|863.30|Injury to small intestine, unspecified site, with open wound into cavity
C0160353|ICD9CM|AB|863.30|Small intest inj NOS-opn
C0160354|ICD9CM|PT|863.31|Injury to duodenum, with open wound into cavity
C0160354|ICD9CM|AB|863.31|Duodenum injury-open
C0160355|ICD9CM|PT|863.39|Other injury to small intestine, with open wound into cavity
C0160355|ICD9CM|AB|863.39|Small intest inj NEC-opn
C0160356|ICD9CM|HT|863.4|Injury to colon or rectum without mention of open wound into cavity
C0160357|ICD9CM|PT|863.40|Injury to colon, unspecified site, without mention of open wound into cavity
C0160357|ICD9CM|AB|863.40|Colon injury NOS-closed
C0160358|ICD9CM|PT|863.41|Injury to ascending [right] colon, without mention of open wound into cavity
C0160358|ICD9CM|AB|863.41|Ascending colon inj-clos
C0160359|ICD9CM|PT|863.42|Injury to transverse colon, without mention of open wound into cavity
C0160359|ICD9CM|AB|863.42|Transverse colon inj-cl
C0160360|ICD9CM|PT|863.43|Injury to descending [left] colon, without mention of open wound into cavity
C0160360|ICD9CM|AB|863.43|Descending colon inj-cl
C0160361|ICD9CM|PT|863.44|Injury to sigmoid colon, without mention of open wound into cavity
C0160361|ICD9CM|AB|863.44|Sigmoid colon inj-closed
C0160362|ICD9CM|PT|863.45|Injury to rectum, without mention of open wound into cavity
C0160362|ICD9CM|AB|863.45|Rectum injury-closed
C0160363|ICD9CM|PT|863.46|Injury to multiple sites in colon and rectum, without mention of open wound into cavity
C0160363|ICD9CM|AB|863.46|Colon inj mult site-clos
C0160365|ICD9CM|HT|863.5|Injury to colon or rectum with open wound into cavity
C0160366|ICD9CM|PT|863.50|Injury to colon, unspecified site, with open wound into cavity
C0160366|ICD9CM|AB|863.50|Colon injury NOS-open
C0160367|ICD9CM|PT|863.51|Injury to ascending [right] colon, with open wound into cavity
C0160367|ICD9CM|AB|863.51|Ascending colon inj-open
C0160368|ICD9CM|PT|863.52|Injury to transverse colon, with open wound into cavity
C0160368|ICD9CM|AB|863.52|Transverse colon inj-opn
C0160369|ICD9CM|PT|863.53|Injury to descending [left] colon, with open wound into cavity
C0160369|ICD9CM|AB|863.53|Descending colon inj-opn
C0160370|ICD9CM|PT|863.54|Injury to sigmoid colon, with open wound into cavity
C0160370|ICD9CM|AB|863.54|Sigmoid colon inj-open
C0160371|ICD9CM|PT|863.55|Injury to rectum, with open wound into cavity
C0160371|ICD9CM|AB|863.55|Rectum injury-open
C0160372|ICD9CM|PT|863.56|Injury to multiple sites in colon and rectum, with open wound into cavity
C0160372|ICD9CM|AB|863.56|Colon inj mult site-open
C0160374|ICD9CM|HT|863.8|Injury to other and unspecified gastrointestinal sites without mention of open wound into cavity
C0160375|ICD9CM|PT|863.80|Injury to gastrointestinal tract, unspecified site, without mention of open wound into cavity
C0160375|ICD9CM|AB|863.80|GI injury NOS-closed
C0160377|ICD9CM|PT|863.82|Injury to pancreas, body, without mention of open wound into cavity
C0160377|ICD9CM|AB|863.82|Pancreas, body inj-close
C0160378|ICD9CM|PT|863.83|Injury to pancreas, tail, without mention of open wound into cavity
C0160378|ICD9CM|AB|863.83|Pancreas, tail inj-close
C0160379|ICD9CM|PT|863.84|Injury to pancreas, multiple and unspecified sites, without mention of open wound into cavity
C0160379|ICD9CM|AB|863.84|Pancreas injury NOS-clos
C0160380|ICD9CM|PT|863.85|Injury to appendix, without mention of open wound into cavity
C0160380|ICD9CM|AB|863.85|Appendix injury-closed
C0160381|ICD9CM|PT|863.89|Injury to other gastrointestinal sites, without mention of open wound into cavity
C0160381|ICD9CM|AB|863.89|GI injury NEC-closed
C0160383|ICD9CM|PT|863.90|Injury to gastrointestinal tract, unspecified site, with open wound into cavity
C0160383|ICD9CM|AB|863.90|GI injury NOS-open
C0160384|ICD9CM|PT|863.91|Injury to pancreas, head, with open wound into cavity
C0160384|ICD9CM|AB|863.91|Pancreas, head inj-open
C0160385|ICD9CM|PT|863.92|Injury to pancreas, body, with open wound into cavity
C0160385|ICD9CM|AB|863.92|Pancreas, body inj-open
C0160386|ICD9CM|PT|863.93|Injury to pancreas, tail, with open wound into cavity
C0160386|ICD9CM|AB|863.93|Pancreas, tail inj-open
C0160387|ICD9CM|PT|863.94|Injury to pancreas, multiple and unspecified sites, with open wound into cavity
C0160387|ICD9CM|AB|863.94|Pancreas injury NOS-open
C0160388|ICD9CM|PT|863.95|Injury to appendix, with open wound into cavity
C0160388|ICD9CM|AB|863.95|Appendix injury-open
C0160389|ICD9CM|PT|863.99|Injury to other gastrointestinal sites, with open wound into cavity
C0160389|ICD9CM|HT|863.9|Injury to other and unspecified gastrointestinal sites, with open wound into cavity
C0160389|ICD9CM|AB|863.99|GI injury NEC-open
C0160390|ICD9CM|HT|864|Injury to liver
C0160392|ICD9CM|HT|864.0|Injury to liver without mention of open wound into cavity
C0160392|ICD9CM|AB|864.00|Liver injury NOS-closed
C0160392|ICD9CM|PT|864.00|Injury to liver without mention of open wound into cavity, unspecified injury
C0160393|ICD9CM|PT|864.01|Injury to liver without mention of open wound into cavity, hematoma and contusion
C0160393|ICD9CM|AB|864.01|Liver hematoma/contusion
C0160394|ICD9CM|PT|864.02|Injury to liver without mention of open wound into cavity, laceration, minor
C0160394|ICD9CM|AB|864.02|Liver laceration, minor
C0160396|ICD9CM|PT|864.04|Injury to liver without mention of open wound into cavity, laceration, major
C0160396|ICD9CM|AB|864.04|Liver laceration, major
C0160397|ICD9CM|PT|864.09|Other injury to liver without mention of open wound into cavity
C0160397|ICD9CM|AB|864.09|Liver injury NEC-closed
C0160399|ICD9CM|HT|864.1|Injury to liver with open wound into cavity
C0160399|ICD9CM|AB|864.10|Liver injury NOS-open
C0160399|ICD9CM|PT|864.10|Injury to liver with open wound into cavity, unspecified injury
C0160400|ICD9CM|PT|864.11|Injury to liver with open wound into cavity, hematoma and contusion
C0160400|ICD9CM|AB|864.11|Liver hematom/contus-opn
C0160401|ICD9CM|PT|864.12|Injury to liver with open wound into cavity, laceration, minor
C0160401|ICD9CM|AB|864.12|Liver lacerat, minor-opn
C0160402|ICD9CM|PT|864.13|Injury to liver with open wound into cavity, laceration, moderate
C0160402|ICD9CM|AB|864.13|Liver lacerat, mod-open
C0160404|ICD9CM|PT|864.19|Other injury to liver with open wound into cavity
C0160404|ICD9CM|AB|864.19|Liver injury NEC-open
C0160405|ICD9CM|HT|865|Injury to spleen
C0160407|ICD9CM|HT|865.0|Injury to spleen without mention of open wound into cavity
C0160407|ICD9CM|AB|865.00|Spleen injury NOS-closed
C0160407|ICD9CM|PT|865.00|Injury to spleen without mention of open wound into cavity, unspecified injury
C0160408|ICD9CM|PT|865.01|Injury to spleen without mention of open wound into cavity, hematoma without rupture of capsule
C0160408|ICD9CM|AB|865.01|Spleen hematoma-closed
C0160409|ICD9CM|PT|865.02|Injury to spleen without mention of open wound into cavity, capsular tears, without major disruption of parenchyma
C0160409|ICD9CM|AB|865.02|Spleen capsular tear
C0160410|ICD9CM|PT|865.03|Injury to spleen without mention of open wound into cavity, laceration extending into parenchyma
C0160410|ICD9CM|AB|865.03|Spleen parenchyma lacer
C0160411|ICD9CM|PT|865.04|Injury to spleen without mention of open wound into cavity, massive parenchymal disruption
C0160411|ICD9CM|AB|865.04|Spleen disruption-clos
C0160412|ICD9CM|PT|865.09|Other injury into spleen without mention of open wound into cavity
C0160412|ICD9CM|AB|865.09|Spleen injury NEC-closed
C0160414|ICD9CM|HT|865.1|Injury to spleen with open wound into cavity
C0160414|ICD9CM|AB|865.10|Spleen injury NOS-open
C0160414|ICD9CM|PT|865.10|Injury to spleen with open wound into cavity, unspecified injury
C0160415|ICD9CM|PT|865.11|Injury to spleen with open wound into cavity, hematoma without rupture of capsule
C0160415|ICD9CM|AB|865.11|Spleen hematoma-open
C0160416|ICD9CM|PT|865.12|Injury to spleen with open wound into cavity, capsular tears, without major disruption of parenchyma
C0160416|ICD9CM|AB|865.12|Spleen capsular tear-opn
C0160417|ICD9CM|PT|865.13|Injury to spleen with open wound into cavity, laceration extending into parenchyma
C0160417|ICD9CM|AB|865.13|Spleen parnchym lac-opn
C0160418|ICD9CM|PT|865.14|Injury to spleen with open wound into cavity, massive parenchyma disruption
C0160418|ICD9CM|AB|865.14|Spleen disruption-open
C0160419|ICD9CM|PT|865.19|Other injury to spleen with open wound into cavity
C0160419|ICD9CM|AB|865.19|Spleen injury NEC-open
C0160420|ICD9CM|HT|866|Injury to kidney
C0160422|ICD9CM|AB|866.00|Kidney injury NOS-closed
C0160422|ICD9CM|HT|866.0|Injury to kidney without mention of open wound into cavity
C0160422|ICD9CM|PT|866.00|Injury to kidney without mention of open wound into cavity, unspecified injury
C0160423|ICD9CM|PT|866.01|Injury to kidney without mention of open wound into cavity, hematoma without rupture of capsule
C0160423|ICD9CM|AB|866.01|Kidney hematoma-closed
C0160424|ICD9CM|AB|866.02|Kidney laceration-closed
C0160424|ICD9CM|PT|866.02|Injury to kidney without mention of open wound into cavity, laceration
C0160427|ICD9CM|HT|866.1|Injury to kidney with open wound into cavity
C0160427|ICD9CM|AB|866.10|Kidney injury NOS-open
C0160427|ICD9CM|PT|866.10|Injury to kidney with open wound into cavity, unspecified injury
C0160428|ICD9CM|AB|866.11|Kidney hematoma-open
C0160428|ICD9CM|PT|866.11|Injury to kidney with open wound into cavity, hematoma without rupture of capsule
C0160429|ICD9CM|AB|866.12|Kidney laceration-open
C0160429|ICD9CM|PT|866.12|Injury to kidney with open wound into cavity, laceration
C0160430|ICD9CM|PT|866.13|Injury to kidney with open wound into cavity, complete disruption of kidney parenchyma
C0160430|ICD9CM|AB|866.13|Kidney disruption-open
C0160432|ICD9CM|PT|867.0|Injury to bladder and urethra, without mention of open wound into cavity
C0160432|ICD9CM|AB|867.0|Bladder/urethra inj-clos
C0160433|ICD9CM|PT|867.1|Injury to bladder and urethra, with open wound into cavity
C0160433|ICD9CM|AB|867.1|Bladder/urethra inj-open
C0160434|ICD9CM|PT|867.2|Injury to ureter, without mention of open wound into cavity
C0160434|ICD9CM|AB|867.2|Ureter injury-closed
C0160435|ICD9CM|PT|867.3|Injury to ureter, with open wound into cavity
C0160435|ICD9CM|AB|867.3|Ureter injury-open
C0160436|ICD9CM|PT|867.4|Injury to uterus, without mention of open wound into cavity
C0160436|ICD9CM|AB|867.4|Uterus injury-closed
C0160437|ICD9CM|PT|867.5|Injury to uterus, with open wound into cavity
C0160437|ICD9CM|AB|867.5|Uterus injury-open
C0160438|ICD9CM|PT|867.6|Injury to other specified pelvic organs, without mention of open wound into cavity
C0160438|ICD9CM|AB|867.6|Pelvic organ inj NEC-cl
C0160439|ICD9CM|PT|867.7|Injury to other specified pelvic organs, with open wound into cavity
C0160439|ICD9CM|AB|867.7|Pelvic organ inj NEC-opn
C0160440|ICD9CM|PT|867.8|Injury to unspecified pelvic organ, without mention of open wound into cavity
C0160440|ICD9CM|AB|867.8|Pelvic organ inj NOS-cl
C0160441|ICD9CM|PT|867.9|Injury to unspecified pelvic organ, with open wound into cavity
C0160441|ICD9CM|AB|867.9|Pelvic organ inj NOS-opn
C0160443|ICD9CM|HT|868.0|Injury to other intra-abdominal organs without mention of open wound into cavity
C0160444|ICD9CM|PT|868.00|Injury to other intra-abdominal organs without mention of open wound into cavity, unspecified intra-abdominal organ
C0160444|ICD9CM|AB|868.00|Intra-abdom inj NOS-clos
C0160445|ICD9CM|PT|868.01|Injury to other intra-abdominal organs without mention of open wound into cavity, adrenal gland
C0160445|ICD9CM|AB|868.01|Adrenal gland injury-cl
C0160446|ICD9CM|PT|868.02|Injury to other intra-abdominal organs without mention of open wound into cavity, bile duct and gallbladder
C0160446|ICD9CM|AB|868.02|Biliary tract injury-cl
C0160447|ICD9CM|AB|868.03|Peritoneum injury-closed
C0160447|ICD9CM|PT|868.03|Injury to other intra-abdominal organs without mention of open wound into cavity, peritoneum
C0160448|ICD9CM|PT|868.04|Injury to other intra-abdominal organs without mention of open wound into cavity, retroperitoneum
C0160448|ICD9CM|AB|868.04|Retroperitoneum inj-cl
C0160449|ICD9CM|PT|868.09|Injury to other and multiple intra-abdominal organs without mention of open wound into cavity
C0160449|ICD9CM|AB|868.09|Intra-abdom inj NEC-clos
C0160450|ICD9CM|HT|868.1|Injury to other intra-abdominal organs with open wound into cavity
C0160451|ICD9CM|PT|868.10|Injury to other intra-abdominal organs with open wound into cavity, unspecified intra-abdominal organ
C0160451|ICD9CM|AB|868.10|Intra-abdom inj NOS-open
C0160452|ICD9CM|PT|868.11|Injury to other intra-abdominal organs with open wound into cavity, adrenal gland
C0160452|ICD9CM|AB|868.11|Adrenal gland injury-opn
C0160453|ICD9CM|PT|868.12|Injury to other intra-abdominal organs with open wound into cavity, bile duct and gallbladder
C0160453|ICD9CM|AB|868.12|Biliary tract injury-opn
C0160454|ICD9CM|AB|868.13|Peritoneum injury-open
C0160454|ICD9CM|PT|868.13|Injury to other intra-abdominal organs with open wound into cavity, peritoneum
C0160455|ICD9CM|PT|868.14|Injury to other intra-abdominal organs with open wound into cavity, retroperitoneum
C0160455|ICD9CM|AB|868.14|Retroperitoneum inj-open
C0160456|ICD9CM|PT|868.19|Injury to other and multiple intra-abdominal organs, with open wound into cavity
C0160456|ICD9CM|AB|868.19|Intra-abdom inj NEC-open
C0160457|ICD9CM|HT|869|Internal injury to unspecified or ill-defined organs
C0160458|ICD9CM|PT|869.1|Internal injury to unspecified or ill-defined organs with open wound into cavity
C0160458|ICD9CM|AB|869.1|Internal injury NOS-open
C0160459|ICD9CM|HT|870|Open wound of ocular adnexa
C0160460|ICD9CM|PT|870.0|Laceration of skin of eyelid and periocular area
C0160460|ICD9CM|AB|870.0|Lac eyelid skn/perioculr
C0160464|ICD9CM|PT|870.4|Penetrating wound of orbit with foreign body
C0160464|ICD9CM|AB|870.4|Penetrat wnd orbit w FB
C0160465|ICD9CM|PT|870.8|Other specified open wounds of ocular adnexa
C0160465|ICD9CM|AB|870.8|Opn wnd ocular adnex NEC
C0160466|ICD9CM|PT|870.9|Unspecified open wound of ocular adnexa
C0160466|ICD9CM|AB|870.9|Opn wnd ocular adnex NOS
C0160468|ICD9CM|PT|871.1|Ocular laceration with prolapse or exposure of intraocular tissue
C0160468|ICD9CM|AB|871.1|Ocular lacera w prolapse
C0160469|ICD9CM|PT|871.2|Rupture of eye with partial loss of intraocular tissue
C0160469|ICD9CM|AB|871.2|Rupture eye w tissu loss
C0160470|ICD9CM|AB|871.4|Laceration of eye NOS
C0160470|ICD9CM|PT|871.4|Unspecified laceration of eye
C0160471|ICD9CM|PT|871.5|Penetration of eyeball with magnetic foreign body
C0160471|ICD9CM|AB|871.5|Penetrat magnet FB eye
C0160472|ICD9CM|PT|871.6|Penetration of eyeball with (nonmagnetic) foreign body
C0160472|ICD9CM|AB|871.6|Penetrat FB NEC eye
C0160474|ICD9CM|HT|871|Open wound of eyeball
C0160474|ICD9CM|PT|871.9|Unspecified open wound of eyeball
C0160474|ICD9CM|AB|871.9|Opn wound of eyeball NOS
C0160475|ICD9CM|HT|872|Open wound of ear
C0160475|ICD9CM|AB|872.8|Open wound of ear NOS
C0160475|ICD9CM|PT|872.8|Open wound of ear, part unspecified, without mention of complication
C0160476|ICD9CM|HT|872.0|Open wound of external ear, without mention of complication
C0160481|ICD9CM|PT|872.10|Open wound of external ear, unspecified site, complicated
C0160481|ICD9CM|AB|872.10|Opn wnd ex ear NOS-compl
C0160482|ICD9CM|PT|872.11|Open wound of auricle, ear, complicated
C0160482|ICD9CM|AB|872.11|Open wound auricle-compl
C0160483|ICD9CM|PT|872.12|Open wound of auditory canal, complicated
C0160483|ICD9CM|AB|872.12|Open wnd aud canal-compl
C0160484|ICD9CM|HT|872.6|Open wound of other specified parts of ear, without mention of complication
C0160489|ICD9CM|HT|872.7|Open wound of other specified parts of ear, complicated
C0160490|ICD9CM|PT|872.71|Open wound of ear drum, complicated
C0160490|ICD9CM|AB|872.71|Open wnd ear drum-compl
C0160491|ICD9CM|PT|872.72|Open wound of ossicles, complicated
C0160491|ICD9CM|AB|872.72|Open wnd ossicles-compl
C0160492|ICD9CM|PT|872.73|Open wound of eustachian tube, complicated
C0160492|ICD9CM|AB|872.73|Opn wnd eustach tb-compl
C0160493|ICD9CM|PT|872.74|Open wound of cochlea, complicated
C0160493|ICD9CM|AB|872.74|Open wound cochlea-compl
C0160496|ICD9CM|HT|873|Other open wound of head
C0160498|ICD9CM|PT|873.1|Open wound of scalp, complicated
C0160498|ICD9CM|AB|873.1|Open wound scalp-compl
C0160502|ICD9CM|AB|873.22|Open wound nasal cavity
C0160502|ICD9CM|PT|873.22|Open wound of nasal cavity, without mention of complication
C0160503|ICD9CM|AB|873.23|Open wound nasal sinus
C0160503|ICD9CM|PT|873.23|Open wound of nasal sinus, without mention of complication
C0160505|ICD9CM|PT|873.30|Open wound of nose, unspecified site, complicated
C0160505|ICD9CM|HT|873.3|Open wound of nose, complicated
C0160505|ICD9CM|AB|873.30|Open wnd nose NOS-compl
C0160507|ICD9CM|PT|873.31|Open wound of nasal septum, complicated
C0160507|ICD9CM|AB|873.31|Opn wnd nas septum-compl
C0160508|ICD9CM|PT|873.32|Open wound of nasal cavity, complicated
C0160508|ICD9CM|AB|873.32|Open wnd nasal cav-compl
C0160509|ICD9CM|PT|873.33|Open wound of nasal sinus, complicated
C0160509|ICD9CM|AB|873.33|Open wnd nas sinus-compl
C0160511|ICD9CM|HT|873.4|Open wound of face, without mention of complication
C0160517|ICD9CM|PT|873.50|Open wound of face, unspecified site, complicated
C0160517|ICD9CM|HT|873.5|Open wound of face, complicated
C0160517|ICD9CM|AB|873.50|Open wnd face NOS-compl
C0160519|ICD9CM|PT|873.51|Open wound of cheek, complicated
C0160519|ICD9CM|AB|873.51|Open wound cheek-compl
C0160520|ICD9CM|PT|873.52|Open wound of forehead, complicated
C0160520|ICD9CM|AB|873.52|Open wnd forehead-compl
C0160521|ICD9CM|PT|873.53|Open wound of lip, complicated
C0160521|ICD9CM|AB|873.53|Open wound lip-complicat
C0160522|ICD9CM|PT|873.54|Open wound of jaw, complicated
C0160522|ICD9CM|AB|873.54|Open wound jaw-complicat
C0160523|ICD9CM|HT|873.6|Open wound of internal structures of mouth, without mention of complication
C0160529|ICD9CM|HT|873.7|Open wound of internal structure of mouth, complicated
C0160531|ICD9CM|PT|873.71|Open wound of buccal mucosa, complicated
C0160531|ICD9CM|AB|873.71|Opn wnd buc mucosa-compl
C0160533|ICD9CM|AB|873.73|Broken tooth-complicated
C0160533|ICD9CM|PT|873.73|Open wound of tooth (broken) (fractured) (due to trauma), complicated
C0160534|ICD9CM|PT|873.74|Open wound of tongue and floor of mouth, complicated
C0160534|ICD9CM|AB|873.74|Open wound tongue-compl
C0160535|ICD9CM|PT|873.75|Open wound of palate, complicated
C0160535|ICD9CM|AB|873.75|Open wound palate-compl
C0160536|ICD9CM|PT|873.8|Other and unspecified open wound of head without mention of complication
C0160536|ICD9CM|AB|873.8|Open wound of head NEC
C0160537|ICD9CM|PT|873.9|Other and unspecified open wound of head, complicated
C0160537|ICD9CM|AB|873.9|Open wnd head NEC-compl
C0160538|ICD9CM|HT|874|Open wound of neck
C0160539|ICD9CM|PT|874.00|Open wound of larynx with trachea, without mention of complication
C0160539|ICD9CM|HT|874.0|Open wound of larynx and trachea, without mention of complication
C0160539|ICD9CM|AB|874.00|Opn wnd larynx w trachea
C0160543|ICD9CM|PT|874.10|Open wound of larynx with trachea, complicated
C0160543|ICD9CM|HT|874.1|Open wound of larynx and trachea, complicated
C0160543|ICD9CM|AB|874.10|Opn wnd lary w trac-comp
C0160544|ICD9CM|PT|874.11|Open wound of larynx, complicated
C0160544|ICD9CM|AB|874.11|Open wound larynx-compl
C0160545|ICD9CM|PT|874.12|Open wound of trachea, complicated
C0160545|ICD9CM|AB|874.12|Open wound trachea-compl
C0160547|ICD9CM|PT|874.3|Open wound of thyroid gland, complicated
C0160547|ICD9CM|AB|874.3|Open wound thyroid-compl
C0160549|ICD9CM|PT|874.5|Open wound of pharynx, complicated
C0160549|ICD9CM|AB|874.5|Open wound pharynx-compl
C0160550|ICD9CM|PT|874.8|Open wound of other and unspecified parts of neck, without mention of complication
C0160550|ICD9CM|AB|874.8|Open wound of neck NEC
C0160551|ICD9CM|PT|874.9|Open wound of other and unspecified parts of neck, complicated
C0160551|ICD9CM|AB|874.9|Opn wound neck NEC-compl
C0160552|ICD9CM|HT|875|Open wound of chest (wall)
C0160555|ICD9CM|HT|876|Open wound of back
C0160557|ICD9CM|PT|876.1|Open wound of back, complicated
C0160557|ICD9CM|AB|876.1|Open wound back-compl
C0160558|ICD9CM|HT|877|Open wound of buttock
C0160560|ICD9CM|PT|877.1|Open wound of buttock, complicated
C0160560|ICD9CM|AB|877.1|Open wound buttock-compl
C0160561|ICD9CM|HT|878|Open wound of genital organs (external), including traumatic amputation
C0160562|ICD9CM|AB|878.0|Open wound of penis
C0160562|ICD9CM|PT|878.0|Open wound of penis, without mention of complication
C0160563|ICD9CM|PT|878.1|Open wound of penis, complicated
C0160563|ICD9CM|AB|878.1|Open wound penis-compl
C0160565|ICD9CM|PT|878.3|Open wound of scrotum and testes, complicated
C0160565|ICD9CM|AB|878.3|Opn wnd scrot/test-compl
C0160567|ICD9CM|PT|878.5|Open wound of vulva, complicated
C0160567|ICD9CM|AB|878.5|Open wound vulva-compl
C0160569|ICD9CM|PT|878.7|Open wound of vagina, complicated
C0160569|ICD9CM|AB|878.7|Open wound vagina-compl
C0160570|ICD9CM|PT|878.8|Open wound of other and unspecified parts of genital organs (external), without mention of complication
C0160570|ICD9CM|AB|878.8|Open wound genital NEC
C0160571|ICD9CM|PT|878.9|Open wound of other and unspecified parts of genital organs (external), complicated
C0160571|ICD9CM|AB|878.9|Opn wnd genital NEC-comp
C0160572|ICD9CM|HT|879|Open wound of other and unspecified sites, except limbs
C0160574|ICD9CM|PT|879.1|Open wound of breast, complicated
C0160574|ICD9CM|AB|879.1|Open wound breast-compl
C0160575|ICD9CM|PT|879.2|Open wound of abdominal wall, anterior, without mention of complication
C0160575|ICD9CM|AB|879.2|Opn wnd anterior abdomen
C0160576|ICD9CM|PT|879.3|Open wound of abdominal wall, anterior, complicated
C0160576|ICD9CM|AB|879.3|Opn wnd ant abdomen-comp
C0160577|ICD9CM|PT|879.4|Open wound of abdominal wall, lateral, without mention of complication
C0160577|ICD9CM|AB|879.4|Opn wnd lateral abdomen
C0160578|ICD9CM|PT|879.5|Open wound of abdominal wall, lateral, complicated
C0160578|ICD9CM|AB|879.5|Opn wnd lat abdomen-comp
C0160579|ICD9CM|PT|879.6|Open wound of other and unspecified parts of trunk, without mention of complication
C0160579|ICD9CM|AB|879.6|Open wound of trunk NEC
C0160580|ICD9CM|PT|879.7|Open wound of other and unspecified parts of trunk, complicated
C0160580|ICD9CM|AB|879.7|Open wnd trunk NEC-compl
C0160584|ICD9CM|HT|880.0|Open wound of shoulder and upper arm, without mention of complication
C0160586|ICD9CM|PT|880.01|Open wound of scapular region, without mention of complication
C0160586|ICD9CM|AB|880.01|Open wound of scapula
C0160587|ICD9CM|PT|880.02|Open wound of axillary region, without mention of complication
C0160587|ICD9CM|AB|880.02|Open wound of axilla
C0160588|ICD9CM|AB|880.03|Open wound of upper arm
C0160588|ICD9CM|PT|880.03|Open wound of upper arm, without mention of complication
C0160590|ICD9CM|HT|880.1|Open wound of shoulder and upper arm, complicated
C0160591|ICD9CM|PT|880.10|Open wound of shoulder region, complicated
C0160591|ICD9CM|AB|880.10|Open wnd shoulder-compl
C0160592|ICD9CM|PT|880.11|Open wound of scapular region, complicated
C0160592|ICD9CM|AB|880.11|Open wound scapula-compl
C0160593|ICD9CM|PT|880.12|Open wound of axillary region, complicated
C0160593|ICD9CM|AB|880.12|Open wound axilla-compl
C0160594|ICD9CM|PT|880.13|Open wound of upper arm, complicated
C0160594|ICD9CM|AB|880.13|Open wnd upper arm-compl
C0160595|ICD9CM|PT|880.19|Open wound of multiple sites of shoulder and upper arm, complicated
C0160595|ICD9CM|AB|880.19|Mult opn wnd should-comp
C0160596|ICD9CM|HT|880.2|Open wound of shoulder and upper arm, with tendon involvement
C0160597|ICD9CM|PT|880.20|Open wound of shoulder region, with tendon involvement
C0160597|ICD9CM|AB|880.20|Opn wnd shouldr w tendon
C0160598|ICD9CM|PT|880.21|Open wound of scapular region, with tendon involvement
C0160598|ICD9CM|AB|880.21|Opn wnd scapula w tendon
C0160599|ICD9CM|PT|880.22|Open wound of axillary region, with tendon involvement
C0160599|ICD9CM|AB|880.22|Open wnd axilla w tendon
C0160600|ICD9CM|PT|880.23|Open wound of upper arm, with tendon involvement
C0160600|ICD9CM|AB|880.23|Open wnd up arm w tendon
C0160601|ICD9CM|PT|880.29|Open wound of multiple sites of shoulder and upper arm, with tendon involvement
C0160601|ICD9CM|AB|880.29|Mlt opn wnd shldr w tend
C0160602|ICD9CM|HT|881|Open wound of elbow, forearm, and wrist
C0160603|ICD9CM|HT|881.0|Open wound of elbow, forearm, and wrist, without mention of complication
C0160604|ICD9CM|AB|881.00|Open wound of forearm
C0160604|ICD9CM|PT|881.00|Open wound of forearm, without mention of complication
C0160605|ICD9CM|AB|881.01|Open wound of elbow
C0160605|ICD9CM|PT|881.01|Open wound of elbow, without mention of complication
C0160606|ICD9CM|PT|881.02|Open wound of wrist, without mention of complication
C0160606|ICD9CM|AB|881.02|Open wound of wrist
C0160607|ICD9CM|HT|881.1|Open wound of elbow, forearm, and wrist, complicated
C0160608|ICD9CM|PT|881.10|Open wound of forearm, complicated
C0160608|ICD9CM|AB|881.10|Open wound forearm-compl
C0160609|ICD9CM|PT|881.11|Open wound of elbow, complicated
C0160609|ICD9CM|AB|881.11|Open wound elbow-complic
C0160610|ICD9CM|PT|881.12|Open wound of wrist, complicated
C0160610|ICD9CM|AB|881.12|Open wound wrist-complic
C0160611|ICD9CM|HT|881.2|Open wound of elbow, forearm, and wrist, with tendon involvement
C0160612|ICD9CM|PT|881.20|Open wound of forearm, with tendon involvement
C0160612|ICD9CM|AB|881.20|Open wnd forearm w tendn
C0160613|ICD9CM|PT|881.21|Open wound of elbow, with tendon involvement
C0160613|ICD9CM|AB|881.21|Opn wound elbow w tendon
C0160614|ICD9CM|PT|881.22|Open wound of wrist, with tendon involvement
C0160614|ICD9CM|AB|881.22|Opn wound wrist w tendon
C0160615|ICD9CM|HT|882|Open wound of hand except finger(s) alone
C0160616|ICD9CM|PT|882.0|Open wound of hand except finger(s) alone, without mention of complication
C0160616|ICD9CM|AB|882.0|Open wound of hand
C0160617|ICD9CM|PT|882.1|Open wound of hand except finger(s) alone, complicated
C0160617|ICD9CM|AB|882.1|Opn wound hand-complicat
C0160618|ICD9CM|PT|882.2|Open wound of hand except finger(s) alone, with tendon involvement
C0160618|ICD9CM|AB|882.2|Open wound hand w tendon
C0160621|ICD9CM|PT|883.1|Open wound of finger(s), complicated
C0160621|ICD9CM|AB|883.1|Open wound finger-compl
C0160622|ICD9CM|PT|883.2|Open wound of finger(s), with tendon involvement
C0160622|ICD9CM|AB|883.2|Open wnd finger w tendon
C0160623|ICD9CM|PT|884.0|Multiple and unspecified open wound of upper limb, without mention of complication
C0160623|ICD9CM|AB|884.0|Open wound arm mult/NOS
C0160625|ICD9CM|PT|884.1|Multiple and unspecified open wound of upper limb, complicated
C0160625|ICD9CM|AB|884.1|Open wound arm NOS-compl
C0160626|ICD9CM|PT|884.2|Multiple and unspecified open wound of upper limb, with tendon involvement
C0160626|ICD9CM|AB|884.2|Opn wnd arm NOS w tendon
C0160627|ICD9CM|HT|885|Traumatic amputation of thumb (complete) (partial)
C0160629|ICD9CM|PT|885.1|Traumatic amputation of thumb (complete)(partial), complicated
C0160629|ICD9CM|AB|885.1|Amputation thumb-compl
C0160630|ICD9CM|HT|886|Traumatic amputation of other finger(s) (complete) (partial)
C0160631|ICD9CM|PT|886.0|Traumatic amputation of other finger(s) (complete) (partial), without mention of complication
C0160631|ICD9CM|AB|886.0|Amputation finger
C0160632|ICD9CM|PT|886.1|Traumatic amputation of other finger(s) (complete) (partial), complicated
C0160632|ICD9CM|AB|886.1|Amputation finger-compl
C0160633|ICD9CM|HT|887|Traumatic amputation of arm and hand (complete) (partial)
C0160634|ICD9CM|PT|887.0|Traumatic amputation of arm and hand (complete) (partial), unilateral, below elbow, without mention of complication
C0160634|ICD9CM|AB|887.0|Amput below elb, unilat
C0160636|ICD9CM|PT|887.2|Traumatic amputation of arm and hand (complete) (partial), unilateral, at or above elbow, without mention of complication
C0160636|ICD9CM|AB|887.2|Amput abv elbow, unilat
C0160638|ICD9CM|PT|887.4|Traumatic amputation of arm and hand (complete) (partial), unilateral, level not specified, without mention of complication
C0160638|ICD9CM|AB|887.4|Amputat arm, unilat NOS
C0160639|ICD9CM|PT|887.5|Traumatic amputation of arm and hand (complete) (partial), unilateral, level not specified, complicated
C0160639|ICD9CM|AB|887.5|Amput arm, unil NOS-comp
C0160640|ICD9CM|PT|887.6|Traumatic amputation of arm and hand (complete) (partial), bilateral [any level], without mention of complication
C0160640|ICD9CM|AB|887.6|Amputation arm, bilat
C0160641|ICD9CM|PT|887.7|Traumatic amputation of arm and hand (complete) (partial), bilateral [any level], complicated
C0160641|ICD9CM|AB|887.7|Amputat arm, bilat-compl
C0160643|ICD9CM|HT|890|Open wound of hip and thigh
C0160644|ICD9CM|PT|890.1|Open wound of hip and thigh, complicated
C0160644|ICD9CM|AB|890.1|Open wnd hip/thigh-compl
C0160645|ICD9CM|PT|890.2|Open wound of hip and thigh, with tendon involvement
C0160645|ICD9CM|AB|890.2|Opn wnd hip/thigh w tend
C0160647|ICD9CM|PT|891.0|Open wound of knee, leg [except thigh], and ankle, without mention of complication
C0160647|ICD9CM|AB|891.0|Open wnd knee/leg/ankle
C0160648|ICD9CM|PT|891.1|Open wound of knee, leg [except thigh], and ankle, complicated
C0160648|ICD9CM|AB|891.1|Open wnd knee/leg-compl
C0160649|ICD9CM|PT|891.2|Open wound of knee, leg [except thigh], and ankle, with tendon involvement
C0160649|ICD9CM|AB|891.2|Opn wnd knee/leg w tendn
C0160650|ICD9CM|HT|892|Open wound of foot except toe(s) alone
C0160651|ICD9CM|PT|892.0|Open wound of foot except toe(s) alone, without mention of complication
C0160651|ICD9CM|AB|892.0|Open wound of foot
C0160652|ICD9CM|PT|892.1|Open wound of foot except toe(s) alone, complicated
C0160652|ICD9CM|AB|892.1|Open wound foot-compl
C0160653|ICD9CM|PT|892.2|Open wound of foot except toe(s) alone, with tendon involvement
C0160653|ICD9CM|AB|892.2|Open wound foot w tendon
C0160655|ICD9CM|PT|893.0|Open wound of toe(s), without mention of complication
C0160655|ICD9CM|AB|893.0|Open wound of toe
C0160658|ICD9CM|HT|894|Multiple and unspecified open wound of lower limb
C0160660|ICD9CM|PT|894.1|Multiple and unspecified open wound of lower limb, complicated
C0160660|ICD9CM|AB|894.1|Open wound leg NEC-compl
C0160661|ICD9CM|PT|894.2|Multiple and unspecified open wound of lower limb, with tendon involvement
C0160661|ICD9CM|AB|894.2|Opn wnd leg NEC w tendon
C0160662|ICD9CM|PT|895.0|Traumatic amputation of toe(s) (complete) (partial), without mention of complication
C0160662|ICD9CM|AB|895.0|Amputation toe
C0160665|ICD9CM|HT|896|Traumatic amputation of foot (complete) (partial)
C0160668|ICD9CM|PT|896.2|Traumatic amputation of foot (complete) (partial), bilateral, without mention of complication
C0160668|ICD9CM|AB|896.2|Amputation foot, bilat
C0160671|ICD9CM|PT|897.0|Traumatic amputation of leg(s) (complete) (partial), unilateral, below knee, without mention of complication
C0160671|ICD9CM|AB|897.0|Amput below knee, unilat
C0160672|ICD9CM|PT|897.1|Traumatic amputation of leg(s) (complete) (partial), unilateral, below knee, complicated
C0160672|ICD9CM|AB|897.1|Amputat bk, unilat-compl
C0160673|ICD9CM|PT|897.2|Traumatic amputation of leg(s) (complete) (partial), unilateral, at or above knee, without mention of complication
C0160673|ICD9CM|AB|897.2|Amput above knee, unilat
C0160674|ICD9CM|PT|897.3|Traumatic amputation of leg(s) (complete) (partial), unilateral, at or above knee, complicated
C0160674|ICD9CM|AB|897.3|Amput abv kn, unil-compl
C0160675|ICD9CM|HT|897|Traumatic amputation of leg(s) (complete) (partial)
C0160676|ICD9CM|PT|897.5|Traumatic amputation of leg(s) (complete) (partial), unilateral, level not specified, complicated
C0160676|ICD9CM|AB|897.5|Amput leg, unil NOS-comp
C0160677|ICD9CM|PT|897.6|Traumatic amputation of leg(s) (complete) (partial), bilateral [any level]), without mention of complication
C0160677|ICD9CM|AB|897.6|Amputation leg, bilat
C0160678|ICD9CM|PT|897.7|Traumatic amputation of leg(s) (complete) (partial), bilateral [any level], complicated
C0160678|ICD9CM|AB|897.7|Amputat leg, bilat-compl
C0160679|ICD9CM|HT|900|Injury to blood vessels of head and neck
C0160679|ICD9CM|PT|900.9|Injury to unspecified blood vessel of head and neck
C0160679|ICD9CM|AB|900.9|Inj head/neck vessel NOS
C0160680|ICD9CM|HT|900.0|Injury to carotid artery
C0160680|ICD9CM|PT|900.00|Injury to carotid artery, unspecified
C0160680|ICD9CM|AB|900.00|Injur carotid artery NOS
C0160681|ICD9CM|PT|900.01|Injury to common carotid artery
C0160681|ICD9CM|AB|900.01|Inj common carotid arter
C0160682|ICD9CM|PT|900.02|Injury to external carotid artery
C0160682|ICD9CM|AB|900.02|Inj external carotid art
C0160683|ICD9CM|PT|900.03|Injury to internal carotid artery
C0160683|ICD9CM|AB|900.03|Inj internal carotid art
C0160684|ICD9CM|PT|900.1|Injury to internal jugular vein
C0160684|ICD9CM|AB|900.1|Inj internl jugular vein
C0160685|ICD9CM|HT|900.8|Injury to other specified blood vessels of head and neck
C0160685|ICD9CM|PT|900.89|Injury to other specified blood vessels of head and neck
C0160685|ICD9CM|AB|900.89|Inj head/neck vessel NEC
C0160686|ICD9CM|PT|900.81|Injury to external jugular vein
C0160686|ICD9CM|AB|900.81|Inj extern jugular vein
C0160687|ICD9CM|PT|900.82|Injury to multiple blood vessels of head and neck
C0160687|ICD9CM|AB|900.82|Inj mlt head/neck vessel
C0160689|ICD9CM|HT|901|Injury to blood vessels of thorax
C0160689|ICD9CM|PT|901.9|Injury to unspecified blood vessel of thorax
C0160689|ICD9CM|AB|901.9|Inj thoracic vessel NOS
C0160690|ICD9CM|PT|901.0|Injury to thoracic aorta
C0160690|ICD9CM|AB|901.0|Injury thoracic aorta
C0160692|ICD9CM|PT|901.2|Injury to superior vena cava
C0160692|ICD9CM|AB|901.2|Inj superior vena cava
C0160693|ICD9CM|PT|901.3|Injury to innominate and subclavian veins
C0160693|ICD9CM|AB|901.3|Inj innomin/subclav vein
C0160696|ICD9CM|PT|901.41|Injury to pulmonary artery
C0160696|ICD9CM|AB|901.41|Injury pulmonary artery
C0160697|ICD9CM|PT|901.42|Injury to pulmonary vein
C0160697|ICD9CM|AB|901.42|Injury pulmonary vein
C0160698|ICD9CM|HT|901.8|Injury to other specified blood vessels of thorax
C0160698|ICD9CM|PT|901.89|Injury to other specified blood vessels of thorax
C0160698|ICD9CM|AB|901.89|Inj thoracic vessel NEC
C0160700|ICD9CM|PT|901.82|Injury to internal mammary artery or vein
C0160700|ICD9CM|AB|901.82|Inj int mammary art/vein
C0160701|ICD9CM|PT|901.83|Injury to multiple blood vessels of thorax
C0160701|ICD9CM|AB|901.83|Inj mult thoracic vessel
C0160703|ICD9CM|HT|902|Injury to blood vessels of abdomen and pelvis
C0160703|ICD9CM|PT|902.9|Injury to unspecified blood vessel of abdomen and pelvis
C0160703|ICD9CM|AB|902.9|Inj abdominal vessel NOS
C0160704|ICD9CM|PT|902.0|Injury to abdominal aorta
C0160704|ICD9CM|AB|902.0|Injury abdominal aorta
C0160705|ICD9CM|HT|902.1|Injury to inferior vena cava
C0160705|ICD9CM|PT|902.10|Injury to inferior vena cava, unspecified
C0160705|ICD9CM|AB|902.10|Inj infer vena cava NOS
C0160706|ICD9CM|PT|902.11|Injury to hepatic veins
C0160706|ICD9CM|AB|902.11|Injury hepatic veins
C0160707|ICD9CM|PT|902.19|Injury to inferior vena cava, other
C0160707|ICD9CM|AB|902.19|Inj infer vena cava NEC
C0160708|ICD9CM|HT|902.2|Injury to celiac and mesenteric arteries
C0160708|ICD9CM|PT|902.20|Injury to celiac and mesenteric arteries, unspecified
C0160708|ICD9CM|AB|902.20|Inj celiac/mesen art NOS
C0160709|ICD9CM|PT|902.21|Injury to gastric artery
C0160709|ICD9CM|AB|902.21|Injury gastric artery
C0160710|ICD9CM|PT|902.22|Injury to hepatic artery
C0160710|ICD9CM|AB|902.22|Injury hepatic artery
C0160711|ICD9CM|PT|902.23|Injury to splenic artery
C0160711|ICD9CM|AB|902.23|Injury splenic artery
C0160712|ICD9CM|PT|902.24|Injury to other specified branches of celiac axis
C0160712|ICD9CM|AB|902.24|Injury celiac axis NEC
C0160714|ICD9CM|PT|902.26|Injury to primary branches of superior mesenteric artery
C0160714|ICD9CM|AB|902.26|Inj brnch sup mesent art
C0160715|ICD9CM|PT|902.27|Injury to inferior mesenteric artery
C0160715|ICD9CM|AB|902.27|Inj infer mesenteric art
C0160716|ICD9CM|PT|902.29|Injury to celiac and mesenteric arteries, other
C0160716|ICD9CM|AB|902.29|Inj mesenteric vess NEC
C0160717|ICD9CM|HT|902.3|Injury to portal and splenic veins
C0160718|ICD9CM|PT|902.31|Injury to superior mesenteric vein and primary subdivisions
C0160718|ICD9CM|AB|902.31|Inj superior mesent vein
C0160719|ICD9CM|PT|902.32|Injury to inferior mesenteric vein
C0160719|ICD9CM|AB|902.32|Inj inferior mesent vein
C0160720|ICD9CM|PT|902.33|Injury to portal vein
C0160720|ICD9CM|AB|902.33|Injury portal vein
C0160721|ICD9CM|PT|902.34|Injury to splenic vein
C0160721|ICD9CM|AB|902.34|Injury splenic vein
C0160722|ICD9CM|PT|902.39|Injury to portal and splenic veins, other
C0160722|ICD9CM|AB|902.39|Inj port/splen vess NEC
C0160723|ICD9CM|HT|902.4|Injury to renal blood vessels
C0160723|ICD9CM|AB|902.40|Injury renal vessel NOS
C0160723|ICD9CM|PT|902.40|Injury to renal vessel(s), unspecified
C0160725|ICD9CM|PT|902.41|Injury to renal artery
C0160725|ICD9CM|AB|902.41|Injury renal artery
C0160726|ICD9CM|PT|902.42|Injury to renal vein
C0160726|ICD9CM|AB|902.42|Injury renal vein
C0160727|ICD9CM|PT|902.49|Injury to renal blood vessels, other
C0160727|ICD9CM|AB|902.49|Injury renal vessel NEC
C0160728|ICD9CM|HT|902.5|Injury to iliac blood vessels
C0160728|ICD9CM|AB|902.50|Injury iliac vessel NOS
C0160728|ICD9CM|PT|902.50|Injury to iliac vessel(s), unspecified
C0160730|ICD9CM|PT|902.51|Injury to hypogastric artery
C0160730|ICD9CM|AB|902.51|Inj hypogastric artery
C0160731|ICD9CM|AB|902.52|Injury hypogastric vein
C0160731|ICD9CM|PT|902.52|Injury to hypogastric vein
C0160732|ICD9CM|PT|902.53|Injury to iliac artery
C0160732|ICD9CM|AB|902.53|Injury iliac artery
C0160733|ICD9CM|PT|902.54|Injury to iliac vein
C0160733|ICD9CM|AB|902.54|Injury iliac vein
C0160734|ICD9CM|PT|902.55|Injury to uterine artery
C0160734|ICD9CM|AB|902.55|Injury uterine artery
C0160735|ICD9CM|PT|902.56|Injury to uterine vein
C0160735|ICD9CM|AB|902.56|Injury uterine vein
C0160736|ICD9CM|PT|902.59|Injury to iliac blood vessels, other
C0160736|ICD9CM|AB|902.59|Injury iliac vessel NEC
C0160737|ICD9CM|HT|902.8|Injury to other specified blood vessels of abdomen and pelvis
C0160737|ICD9CM|PT|902.89|Injury to other specified blood vessels of abdomen and pelvis
C0160737|ICD9CM|AB|902.89|Inj abdominal vessel NEC
C0160738|ICD9CM|PT|902.81|Injury to ovarian artery
C0160738|ICD9CM|AB|902.81|Injury ovarian artery
C0160739|ICD9CM|PT|902.82|Injury to ovarian vein
C0160739|ICD9CM|AB|902.82|Injury ovarian vein
C0160740|ICD9CM|PT|902.87|Injury to multiple blood vessels of abdomen and pelvis
C0160740|ICD9CM|AB|902.87|Inj mult abd/pelv vessel
C0160742|ICD9CM|HT|903|Injury to blood vessels of upper extremity
C0160742|ICD9CM|PT|903.9|Injury to unspecified blood vessel of upper extremity
C0160742|ICD9CM|AB|903.9|Injury arm vessel NOS
C0160745|ICD9CM|PT|903.01|Injury to axillary artery
C0160745|ICD9CM|AB|903.01|Injury axillary artery
C0160746|ICD9CM|PT|903.02|Injury to axillary vein
C0160746|ICD9CM|AB|903.02|Injury axillary vein
C0160748|ICD9CM|PT|903.2|Injury to radial blood vessels
C0160748|ICD9CM|AB|903.2|Injury radial vessels
C0160749|ICD9CM|PT|903.3|Injury to ulnar blood vessels
C0160749|ICD9CM|AB|903.3|Injury ulnar vessels
C0160750|ICD9CM|PT|903.4|Injury to palmar artery
C0160750|ICD9CM|AB|903.4|Injury palmar artery
C0160751|ICD9CM|PT|903.5|Injury to digital blood vessels
C0160751|ICD9CM|AB|903.5|Injury finger vessels
C0160752|ICD9CM|PT|903.8|Injury to other specified blood vessels of upper extremity
C0160752|ICD9CM|AB|903.8|Injury arm vessels NEC
C0160754|ICD9CM|HT|904|Injury to blood vessels of lower extremity and unspecified sites
C0160755|ICD9CM|PT|904.0|Injury to common femoral artery
C0160755|ICD9CM|AB|904.0|Inj common femoral arter
C0160756|ICD9CM|PT|904.1|Injury to superficial femoral artery
C0160756|ICD9CM|AB|904.1|Inj superfic femoral art
C0160757|ICD9CM|PT|904.2|Injury to femoral veins
C0160757|ICD9CM|AB|904.2|Injury femoral vein
C0160758|ICD9CM|PT|904.3|Injury to saphenous veins
C0160758|ICD9CM|AB|904.3|Injury saphenous vein
C0160761|ICD9CM|PT|904.41|Injury to popliteal artery
C0160761|ICD9CM|AB|904.41|Injury popliteal artery
C0160762|ICD9CM|PT|904.42|Injury to popliteal vein
C0160762|ICD9CM|AB|904.42|Injury popliteal vein
C0160763|ICD9CM|HT|904.5|Injury to tibial blood vessels
C0160763|ICD9CM|AB|904.50|Injury tibial vessel NOS
C0160763|ICD9CM|PT|904.50|Injury to tibial vessel(s), unspecified
C0160765|ICD9CM|PT|904.51|Injury to anterior tibial artery
C0160765|ICD9CM|AB|904.51|Inj anter tibial artery
C0160766|ICD9CM|PT|904.52|Injury to anterior tibial vein
C0160766|ICD9CM|AB|904.52|Inj anterior tibial vein
C0160767|ICD9CM|PT|904.53|Injury to posterior tibial artery
C0160767|ICD9CM|AB|904.53|Inj post tibial artery
C0160768|ICD9CM|PT|904.54|Injury to posterior tibial vein
C0160768|ICD9CM|AB|904.54|Inj post tibial vein
C0160769|ICD9CM|PT|904.6|Injury to deep plantar blood vessels
C0160769|ICD9CM|AB|904.6|Inj deep plantar vessel
C0160770|ICD9CM|PT|904.7|Injury to other specified blood vessels of lower extremity
C0160770|ICD9CM|AB|904.7|Injury leg vessels NEC
C0160773|ICD9CM|HT|905|Late effects of musculoskeletal and connective tissue injuries
C0160774|ICD9CM|PT|905.0|Late effect of fracture of skull and face bones
C0160774|ICD9CM|AB|905.0|Late effec skull/face fx
C0160777|ICD9CM|PT|905.3|Late effect of fracture of neck of femur
C0160777|ICD9CM|AB|905.3|Late eff femoral neck fx
C0160778|ICD9CM|PT|905.4|Late effect of fracture of lower extremities
C0160778|ICD9CM|AB|905.4|Late effect leg fx
C0160779|ICD9CM|PT|905.5|Late effect of fracture of multiple and unspecified bones
C0160779|ICD9CM|AB|905.5|Late effect fracture NEC
C0160780|ICD9CM|PT|905.6|Late effect of dislocation
C0160780|ICD9CM|AB|905.6|Late effect dislocation
C0160781|ICD9CM|PT|905.7|Late effect of sprain and strain without mention of tendon injury
C0160781|ICD9CM|AB|905.7|Late effec sprain/strain
C0160782|ICD9CM|PT|905.8|Late effect of tendon injury
C0160782|ICD9CM|AB|905.8|Late effec tendon injury
C0160783|ICD9CM|PT|905.9|Late effect of traumatic amputation
C0160783|ICD9CM|AB|905.9|Late eff traumat amputat
C0160784|ICD9CM|HT|906|Late effects of injuries to skin and subcutaneous tissues
C0160785|ICD9CM|PT|906.0|Late effect of open wound of head, neck, and trunk
C0160785|ICD9CM|AB|906.0|Lt eff opn wnd head/trnk
C0160786|ICD9CM|PT|906.1|Late effect of open wound of extremities without mention of tendon injury
C0160786|ICD9CM|AB|906.1|Late eff open wnd extrem
C0160787|ICD9CM|PT|906.2|Late effect of superficial injury
C0160787|ICD9CM|AB|906.2|Late eff superficial inj
C0160788|ICD9CM|AB|906.3|Late effect of contusion
C0160788|ICD9CM|PT|906.3|Late effect of contusion
C0160790|ICD9CM|PT|906.5|Late effect of burn of eye, face, head, and neck
C0160790|ICD9CM|AB|906.5|Late eff head/neck burn
C0160791|ICD9CM|PT|906.6|Late effect of burn of wrist and hand
C0160791|ICD9CM|AB|906.6|Late eff wrist/hand burn
C0160792|ICD9CM|PT|906.7|Late effect of burn of other extremities
C0160792|ICD9CM|AB|906.7|Late eff burn extrem NEC
C0160793|ICD9CM|PT|906.8|Late effect of burns of other specified sites
C0160793|ICD9CM|AB|906.8|Late effect of burns NEC
C0160794|ICD9CM|PT|906.9|Late effect of burn of unspecified site
C0160794|ICD9CM|AB|906.9|Late effect of burn NOS
C0160795|ICD9CM|HT|907|Late effects of injuries to the nervous system
C0160796|ICD9CM|PT|907.1|Late effect of injury to cranial nerve
C0160796|ICD9CM|AB|907.1|Late eff cran nerve inj
C0160797|ICD9CM|PT|907.2|Late effect of spinal cord injury
C0160797|ICD9CM|AB|907.2|Late eff spinal cord inj
C0160798|ICD9CM|PT|907.3|Late effect of injury to nerve root(s), spinal plexus(es), and other nerves of trunk
C0160798|ICD9CM|AB|907.3|Lt eff nerv inj trnk NEC
C0160799|ICD9CM|PT|907.4|Late effect of injury to peripheral nerve of shoulder girdle and upper limb
C0160799|ICD9CM|AB|907.4|Lt eff nerv inj shld/arm
C0160800|ICD9CM|PT|907.5|Late effect of injury to peripheral nerve of pelvic girdle and lower limb
C0160800|ICD9CM|AB|907.5|Lt eff nerv inj pelv/leg
C0160801|ICD9CM|PT|907.9|Late effect of injury to other and unspecified nerve
C0160801|ICD9CM|AB|907.9|Late eff nerve inj NEC
C0160802|ICD9CM|HT|908|Late effects of other and unspecified injuries
C0160803|ICD9CM|PT|908.0|Late effect of internal injury to chest
C0160803|ICD9CM|AB|908.0|Late eff int injur chest
C0160805|ICD9CM|PT|908.2|Late effect of internal injury to other internal organs
C0160805|ICD9CM|AB|908.2|Late eff int injury NEC
C0160806|ICD9CM|PT|908.3|Late effect of injury to blood vessel of head, neck, and extremities
C0160806|ICD9CM|AB|908.3|Late eff inj periph vess
C0160807|ICD9CM|PT|908.4|Late effect of injury to blood vessel of thorax, abdomen, and pelvis
C0160807|ICD9CM|AB|908.4|Lt eff inj thor/abd vess
C0160808|ICD9CM|PT|908.5|Late effect of foreign body in orifice
C0160808|ICD9CM|AB|908.5|Late eff FB in orifice
C0160809|ICD9CM|PT|908.6|Late effect of certain complications of trauma
C0160809|ICD9CM|AB|908.6|Late eff complic trauma
C0160814|ICD9CM|AB|909.2|Late effect of radiation
C0160814|ICD9CM|PT|909.2|Late effect of radiation
C0160816|ICD9CM|PT|909.4|Late effect of certain other external causes
C0160816|ICD9CM|AB|909.4|Late eff cert ext cause
C0160818|ICD9CM|HT|910|Superficial injury of face, neck, and scalp except eye
C0160819|ICD9CM|PT|910.0|Abrasion or friction burn of face, neck, and scalp except eye, without mention of infection
C0160819|ICD9CM|AB|910.0|Abrasion head
C0160820|ICD9CM|PT|910.1|Abrasion or friction burn of face, neck, and scalp except eye, infected
C0160820|ICD9CM|AB|910.1|Abrasion head-infected
C0160821|ICD9CM|PT|910.2|Blister of face, neck, and scalp except eye, without mention of infection
C0160821|ICD9CM|AB|910.2|Blister head
C0160822|ICD9CM|PT|910.3|Blister of face, neck, and scalp except eye, infected
C0160822|ICD9CM|AB|910.3|Blister head-infected
C0160823|ICD9CM|PT|910.4|Insect bite, nonvenomous of face, neck, and scalp except eye, without mention of infection
C0160823|ICD9CM|AB|910.4|Insect bite head
C0160824|ICD9CM|PT|910.5|Insect bite, nonvenomous of face, neck, and scalp except eye, infected
C0160824|ICD9CM|AB|910.5|Insect bite head-infect
C0160825|ICD9CM|PT|910.6|Superficial foreign body (splinter) of face, neck, and scalp except eye, without major open wound and without mention of infection
C0160825|ICD9CM|AB|910.6|Foreign body head
C0160826|ICD9CM|PT|910.7|Superficial foreign body (splinter) of face, neck, and scalp except eye, without major open wound, infected
C0160826|ICD9CM|AB|910.7|Foreign body head-infect
C0160827|ICD9CM|PT|910.8|Other and unspecified superficial injury of face, neck, and scalp, without mention of infection
C0160827|ICD9CM|AB|910.8|Superfic inj head NEC
C0160828|ICD9CM|PT|910.9|Other and unspecified superficial injury of face, neck, and scalp, infected
C0160828|ICD9CM|AB|910.9|Superf inj head NEC-inf
C0160829|ICD9CM|HT|911|Superficial injury of trunk
C0160830|ICD9CM|PT|911.0|Abrasion or friction burn of trunk, without mention of infection
C0160830|ICD9CM|AB|911.0|Abrasion trunk
C0160831|ICD9CM|PT|911.1|Abrasion or friction burn of trunk, infected
C0160831|ICD9CM|AB|911.1|Abrasion trunk-infected
C0160832|ICD9CM|PT|911.2|Blister of trunk, without mention of infection
C0160832|ICD9CM|AB|911.2|Blister trunk
C0160833|ICD9CM|PT|911.3|Blister of trunk, infected
C0160833|ICD9CM|AB|911.3|Blister trunk-infected
C0160836|ICD9CM|PT|911.6|Superficial foreign body (splinter) of trunk, without major open wound and without mention of infection
C0160836|ICD9CM|AB|911.6|Foreign body trunk
C0160837|ICD9CM|PT|911.7|Superficial foreign body (splinter) of trunk, without major open wound, infected
C0160837|ICD9CM|AB|911.7|Foreign body trunk-infec
C0160839|ICD9CM|PT|911.9|Other and unspecified superficial injury of trunk, infected
C0160839|ICD9CM|AB|911.9|Superf inj trnk NEC-inf
C0160840|ICD9CM|HT|912|Superficial injury of shoulder and upper arm
C0160841|ICD9CM|PT|912.0|Abrasion or friction burn of shoulder and upper arm, without mention of infection
C0160841|ICD9CM|AB|912.0|Abrasion shoulder/arm
C0160842|ICD9CM|PT|912.1|Abrasion or friction burn of shoulder and upper arm, infected
C0160842|ICD9CM|AB|912.1|Abrasion shldr/arm-infec
C0160843|ICD9CM|PT|912.2|Blister of shoulder and upper arm, without mention of infection
C0160843|ICD9CM|AB|912.2|Blister shoulder & arm
C0160844|ICD9CM|PT|912.3|Blister of shoulder and upper arm, infected
C0160844|ICD9CM|AB|912.3|Blister shoulder/arm-inf
C0160845|ICD9CM|PT|912.4|Insect bite, nonvenomous of shoulder and upper arm, without mention of infection
C0160845|ICD9CM|AB|912.4|Insect bite shoulder/arm
C0160846|ICD9CM|PT|912.5|Insect bite, nonvenomous of shoulder and upper arm, infected
C0160846|ICD9CM|AB|912.5|Insect bite shld/arm-inf
C0160847|ICD9CM|PT|912.6|Superficial foreign body (splinter) of shoulder and upper arm, without major open wound and without mention of infection
C0160847|ICD9CM|AB|912.6|Foreign body shouldr/arm
C0160848|ICD9CM|PT|912.7|Superficial foreign body (splinter) of shoulder and upper arm, without major open wound, infected
C0160848|ICD9CM|AB|912.7|FB shoulder/arm-infect
C0160850|ICD9CM|PT|912.9|Other and unspecified superficial injury of shoulder and upper arm, infected
C0160850|ICD9CM|AB|912.9|Superf inj shldr NEC-inf
C0160851|ICD9CM|HT|913|Superficial injury of elbow, forearm, and wrist
C0160852|ICD9CM|PT|913.0|Abrasion or friction burn of elbow, forearm, and wrist, without mention of infection
C0160852|ICD9CM|AB|913.0|Abrasion forearm
C0160853|ICD9CM|PT|913.1|Abrasion or friction burn of elbow, forearm, and wrist, infected
C0160853|ICD9CM|AB|913.1|Abrasion forearm-infect
C0160854|ICD9CM|PT|913.2|Blister of elbow, forearm, and wrist, without mention of infection
C0160854|ICD9CM|AB|913.2|Blister forearm
C0160855|ICD9CM|PT|913.3|Blister of elbow, forearm, and wrist, infected
C0160855|ICD9CM|AB|913.3|Blister forearm-infected
C0160856|ICD9CM|PT|913.4|Insect bite, nonvenomous of elbow, forearm, and wrist, without mention of infection
C0160856|ICD9CM|AB|913.4|Insect bite forearm
C0160857|ICD9CM|PT|913.5|Insect bite, nonvenomous, of elbow, forearm, and wrist, infected
C0160857|ICD9CM|AB|913.5|Insect bite forearm-inf
C0160858|ICD9CM|PT|913.6|Superficial foreign body (splinter) of elbow, forearm, and wrist, without major open wound and without mention of infection
C0160858|ICD9CM|AB|913.6|Foreign body forearm
C0160859|ICD9CM|PT|913.7|Superficial foreign body (splinter) of elbow, forearm, and wrist, without major open wound, infected
C0160859|ICD9CM|AB|913.7|Foreign body forearm-inf
C0160860|ICD9CM|PT|913.8|Other and unspecified superficial injury of elbow, forearm, and wrist, without mention of infection
C0160860|ICD9CM|AB|913.8|Superf inj forearm NEC
C0160861|ICD9CM|PT|913.9|Other and unspecified superficial injury of elbow, forearm, and wrist, infected
C0160861|ICD9CM|AB|913.9|Suprf inj forarm NEC-inf
C0160863|ICD9CM|PT|914.0|Abrasion or friction burn of hand(s) except finger(s) alone, without mention of infection
C0160863|ICD9CM|AB|914.0|Abrasion hand
C0160864|ICD9CM|PT|914.1|Abrasion or friction burn of hand(s) except finger(s) alone, infected
C0160864|ICD9CM|AB|914.1|Abrasion hand-infected
C0160865|ICD9CM|PT|914.2|Blister of hand(s) except finger(s) alone, without mention of infection
C0160865|ICD9CM|AB|914.2|Blister hand
C0160866|ICD9CM|PT|914.3|Blister of hand(s) except finger(s) alone, infected
C0160866|ICD9CM|AB|914.3|Blister hand-infected
C0160867|ICD9CM|PT|914.4|Insect bite, nonvenomous, of hand(s) except finger(s) alone, without mention of infection
C0160867|ICD9CM|AB|914.4|Insect bite hand
C0160868|ICD9CM|PT|914.5|Insect bite, nonvenomous, of hand(s) except finger(s) alone, infected
C0160868|ICD9CM|AB|914.5|Insect bite hand-infect
C0160869|ICD9CM|PT|914.6|Superficial foreign body (splinter) of hand(s) except finger(s) alone, without major open wound and without mention of infection
C0160869|ICD9CM|AB|914.6|Foreign body hand
C0160870|ICD9CM|PT|914.7|Superficial foreign body (splinter) of hand(s) except finger(s) alone, without major open wound, infected
C0160870|ICD9CM|AB|914.7|Foreign body hand-infect
C0160871|ICD9CM|PT|914.8|Other and unspecified superficial injury of hand(s) except finger(s) alone, without mention of infection
C0160871|ICD9CM|AB|914.8|Superficial inj hand NEC
C0160872|ICD9CM|PT|914.9|Other and unspecified superficial injury of hand(s) except finger(s) alone, infected
C0160872|ICD9CM|AB|914.9|Superf inj hand NEC-inf
C0160875|ICD9CM|PT|915.1|Abrasion or friction burn of finger(s), infected
C0160875|ICD9CM|AB|915.1|Abrasion finger-infected
C0160876|ICD9CM|PT|915.2|Blister of finger(s), without mention of infection
C0160876|ICD9CM|AB|915.2|Blister finger
C0160877|ICD9CM|AB|915.3|Blister finger-infected
C0160877|ICD9CM|PT|915.3|Blister of finger(s), infected
C0160879|ICD9CM|PT|915.5|Insect bite, nonvenomous of finger(s), infected
C0160879|ICD9CM|AB|915.5|Insect bite finger-infec
C0160880|ICD9CM|PT|915.6|Superficial foreign body (splinter) of finger(s), without major open wound and without mention of infection
C0160880|ICD9CM|AB|915.6|Foreign body finger
C0160881|ICD9CM|PT|915.7|Superficial foreign body (splinter) of finger(s), without major open wound, infected
C0160881|ICD9CM|AB|915.7|Foreign body finger-inf
C0160882|ICD9CM|PT|915.8|Other and unspecified superficial injury of fingers without mention of infection
C0160882|ICD9CM|AB|915.8|Superfic inj finger-NEC
C0160883|ICD9CM|PT|915.9|Other and unspecified superficial injury of fingers, infected
C0160883|ICD9CM|AB|915.9|Suprf inj finger NEC-inf
C0160884|ICD9CM|HT|916|Superficial injury of hip, thigh, leg, and ankle
C0160885|ICD9CM|PT|916.0|Abrasion or friction burn of hip, thigh, leg, and ankle, without mention of infection
C0160885|ICD9CM|AB|916.0|Abrasion hip & leg
C0160886|ICD9CM|PT|916.1|Abrasion or friction burn of hip, thigh, leg, and ankle, infected
C0160886|ICD9CM|AB|916.1|Abrasion hip/leg-infect
C0160887|ICD9CM|PT|916.2|Blister of hip, thigh, leg, and ankle, without mention of infection
C0160887|ICD9CM|AB|916.2|Blister hip & leg
C0160888|ICD9CM|PT|916.3|Blister of hip, thigh, leg, and ankle, infected
C0160888|ICD9CM|AB|916.3|Blister hip & leg-infect
C0160889|ICD9CM|PT|916.4|Insect bite, nonvenomous, of hip, thigh, leg, and ankle, without mention of infection
C0160889|ICD9CM|AB|916.4|Insect bite hip & leg
C0160890|ICD9CM|PT|916.5|Insect bite, nonvenomous of hip, thigh, leg, and ankle, infected
C0160890|ICD9CM|AB|916.5|Insect bite hip/leg-inf
C0160891|ICD9CM|PT|916.6|Superficial foreign body (splinter) of hip, thigh, leg, and ankle, without major open wound and without mention of infection
C0160891|ICD9CM|AB|916.6|Foreign body hip/leg
C0160892|ICD9CM|PT|916.7|Superficial foreign body (splinter) of hip, thigh, leg, and ankle, without major open wound, infected
C0160892|ICD9CM|AB|916.7|Foreign bdy hip/leg-inf
C0160893|ICD9CM|PT|916.8|Other and unspecified superficial injury of hip, thigh, leg, and ankle, without mention of infection
C0160893|ICD9CM|AB|916.8|Superfic inj hip/leg NEC
C0160894|ICD9CM|PT|916.9|Other and unspecified superficial injury of hip, thigh, leg, and ankle, infected
C0160894|ICD9CM|AB|916.9|Superf inj leg NEC-infec
C0160895|ICD9CM|HT|917|Superficial injury of foot and toe(s)
C0160902|ICD9CM|PT|917.6|Superficial foreign body (splinter) of foot and toe(s), without major open wound and without mention of infection
C0160902|ICD9CM|AB|917.6|Foreign body foot & toe
C0160903|ICD9CM|PT|917.7|Superficial foreign body (splinter) of foot and toe(s), without major open wound, infected
C0160903|ICD9CM|AB|917.7|Foreign bdy foot/toe-inf
C0160904|ICD9CM|PT|917.8|Other and unspecified superficial injury of foot and toes, without mention of infection
C0160904|ICD9CM|AB|917.8|Superf inj foot/toe NEC
C0160905|ICD9CM|PT|917.9|Other and unspecified superficial injury of foot and toes, infected
C0160905|ICD9CM|AB|917.9|Superf inj foot NEC-inf
C0160906|ICD9CM|HT|918|Superficial injury of eye and adnexa
C0160907|ICD9CM|PT|918.0|Superficial injury of eyelids and periocular area
C0160907|ICD9CM|AB|918.0|Superfic inj periocular
C0160908|ICD9CM|PT|918.2|Superficial injury of conjunctiva
C0160908|ICD9CM|AB|918.2|Superfic inj conjunctiva
C0160909|ICD9CM|PT|918.9|Other and unspecified superficial injuries of eye
C0160909|ICD9CM|AB|918.9|Superficial inj eye NEC
C0160910|ICD9CM|HT|919|Superficial injury of other, multiple, and unspecified sites
C0160911|ICD9CM|PT|919.1|Abrasion or friction burn of other, multiple, and unspecified sites, infected
C0160911|ICD9CM|AB|919.1|Abrasion NEC-infected
C0160912|ICD9CM|PT|919.3|Blister of other, multiple, and unspecified sites, infected
C0160912|ICD9CM|AB|919.3|Blister NEC-infected
C0160913|ICD9CM|PT|919.5|Insect bite, nonvenomous, of other, multiple, and unspecified sites, infected
C0160913|ICD9CM|AB|919.5|Insect bite NEC-infected
C0160914|ICD9CM|PT|919.6|Superficial foreign body (splinter) of other, multiple, and unspecified sites, without major open wound and without mention of infection
C0160914|ICD9CM|AB|919.6|Superfic foreign bdy NEC
C0160915|ICD9CM|PT|919.7|Superficial foreign body (splinter) of other, multiple, and unspecified sites, without major open wound, infected
C0160915|ICD9CM|AB|919.7|Superficial FB NEC-infec
C0160916|ICD9CM|PT|919.8|Other and unspecified superficial injury of other, multiple, and unspecified sites, without mention of infection
C0160916|ICD9CM|AB|919.8|Superficial injury NEC
C0160917|ICD9CM|PT|919.9|Other and unspecified superficial injury of other, multiple, and unspecified sites, infected
C0160917|ICD9CM|AB|919.9|Superfic inj NEC-infect
C0160918|ICD9CM|PT|920|Contusion of face, scalp, and neck except eye(s)
C0160918|ICD9CM|AB|920|Contusion face/scalp/nck
C0160919|ICD9CM|HT|921|Contusion of eye and adnexa
C0160920|ICD9CM|PT|921.1|Contusion of eyelids and periocular area
C0160920|ICD9CM|AB|921.1|Contusion periocular
C0160921|ICD9CM|PT|921.2|Contusion of orbital tissues
C0160921|ICD9CM|AB|921.2|Contusion orbital tissue
C0160923|ICD9CM|HT|922|Contusion of trunk
C0160923|ICD9CM|AB|922.9|Contusion trunk NOS
C0160923|ICD9CM|PT|922.9|Contusion of unspecified part of trunk
C0160924|ICD9CM|AB|922.0|Contusion of breast
C0160924|ICD9CM|PT|922.0|Contusion of breast
C0160925|ICD9CM|AB|922.1|Contusion of chest wall
C0160925|ICD9CM|PT|922.1|Contusion of chest wall
C0160926|ICD9CM|PT|922.2|Contusion of abdominal wall
C0160926|ICD9CM|AB|922.2|Contusion abdominal wall
C0160927|ICD9CM|HT|922.3|Contusion of back
C0160927|ICD9CM|PT|922.31|Contusion of back
C0160927|ICD9CM|AB|922.31|Back contusion
C0160928|ICD9CM|PT|922.4|Contusion of genital organs
C0160928|ICD9CM|AB|922.4|Contusion genital organs
C0160929|ICD9CM|PT|922.8|Contusion of multiple sites of trunk
C0160929|ICD9CM|AB|922.8|Multiple contusion trunk
C0160931|ICD9CM|HT|923|Contusion of upper limb
C0160931|ICD9CM|AB|923.9|Contusion upper limb NOS
C0160931|ICD9CM|PT|923.9|Contusion of unspecified part of upper limb
C0160932|ICD9CM|HT|923.0|Contusion of shoulder and upper arm
C0160933|ICD9CM|PT|923.00|Contusion of shoulder region
C0160933|ICD9CM|AB|923.00|Contusion shoulder reg
C0160934|ICD9CM|PT|923.01|Contusion of scapular region
C0160934|ICD9CM|AB|923.01|Contusion scapul region
C0160935|ICD9CM|PT|923.02|Contusion of axillary region
C0160935|ICD9CM|AB|923.02|Contusion axillary reg
C0160936|ICD9CM|AB|923.03|Contusion of upper arm
C0160936|ICD9CM|PT|923.03|Contusion of upper arm
C0160937|ICD9CM|PT|923.09|Contusion of multiple sites of shoulder and upper arm
C0160937|ICD9CM|AB|923.09|Contusion shoulder & arm
C0160938|ICD9CM|HT|923.1|Contusion of elbow and forearm
C0160941|ICD9CM|HT|923.2|Contusion of wrist and hand(s), except finger(s) alone
C0160943|ICD9CM|AB|923.21|Contusion of wrist
C0160943|ICD9CM|PT|923.21|Contusion of wrist
C0160945|ICD9CM|PT|923.8|Contusion of multiple sites of upper limb
C0160945|ICD9CM|AB|923.8|Multiple contusion arm
C0160947|ICD9CM|HT|924|Contusion of lower limb and of other and unspecified sites
C0160948|ICD9CM|HT|924.0|Contusion of hip and thigh
C0160949|ICD9CM|AB|924.00|Contusion of thigh
C0160949|ICD9CM|PT|924.00|Contusion of thigh
C0160950|ICD9CM|AB|924.01|Contusion of hip
C0160950|ICD9CM|PT|924.01|Contusion of hip
C0160951|ICD9CM|HT|924.1|Contusion of knee and lower leg
C0160952|ICD9CM|AB|924.10|Contusion of lower leg
C0160952|ICD9CM|PT|924.10|Contusion of lower leg
C0160953|ICD9CM|AB|924.11|Contusion of knee
C0160953|ICD9CM|PT|924.11|Contusion of knee
C0160955|ICD9CM|AB|924.20|Contusion of foot
C0160955|ICD9CM|PT|924.20|Contusion of foot
C0160956|ICD9CM|AB|924.21|Contusion of ankle
C0160956|ICD9CM|PT|924.21|Contusion of ankle
C0160957|ICD9CM|AB|924.3|Contusion of toe
C0160957|ICD9CM|PT|924.3|Contusion of toe
C0160958|ICD9CM|PT|924.4|Contusion of multiple sites of lower limb
C0160958|ICD9CM|AB|924.4|Multiple contusion leg
C0160960|MTH|PN|NOCODE|Contusion of multiple sites, NEC in ICD9CM_2014
C0160960|ICD9CM|PT|924.8|Contusion of multiple sites, not elsewhere classified
C0160960|ICD9CM|AB|924.8|Multiple contusions NEC
C0160961|ICD9CM|HT|925|Crushing injury of face, scalp, and neck
C0160962|ICD9CM|HT|926|Crushing injury of trunk
C0160962|ICD9CM|PT|926.9|Crushing injury of unspecified site of trunk
C0160962|ICD9CM|AB|926.9|Crushing inj trunk NOS
C0160963|ICD9CM|PT|926.0|Crushing injury of external genitalia
C0160963|ICD9CM|AB|926.0|Crush inj ext genitalia
C0160964|ICD9CM|HT|926.1|Crushing injury of other specified sites of trunk
C0160964|ICD9CM|PT|926.19|Crushing injury of other specified sites of trunk
C0160964|ICD9CM|AB|926.19|Crushing inj trunk NEC
C0160965|ICD9CM|PT|926.11|Crushing injury of back
C0160965|ICD9CM|AB|926.11|Crushing injury back
C0160966|ICD9CM|PT|926.12|Crushing injury of buttock
C0160966|ICD9CM|AB|926.12|Crushing injury buttock
C0160967|ICD9CM|PT|926.8|Crushing injury of multiple sites of trunk
C0160967|ICD9CM|AB|926.8|Mult crushing inj trunk
C0160969|ICD9CM|HT|927|Crushing injury of upper limb
C0160969|ICD9CM|PT|927.9|Crushing injury of unspecified site of upper limb
C0160969|ICD9CM|AB|927.9|Crushing injury arm NOS
C0160970|ICD9CM|HT|927.0|Crushing injury of shoulder and upper arm
C0160971|ICD9CM|PT|927.00|Crushing injury of shoulder region
C0160971|ICD9CM|AB|927.00|Crush inj shoulder reg
C0160972|ICD9CM|PT|927.01|Crushing injury of scapular region
C0160972|ICD9CM|AB|927.01|Crush inj scapul region
C0160973|ICD9CM|PT|927.02|Crushing injury of axillary region
C0160973|ICD9CM|AB|927.02|Crush inj axillary reg
C0160974|ICD9CM|PT|927.03|Crushing injury of upper arm
C0160974|ICD9CM|AB|927.03|Crushing inj upper arm
C0160975|ICD9CM|PT|927.09|Crushing injury of multiple sites of upper arm
C0160975|ICD9CM|AB|927.09|Crush inj shoulder & arm
C0160976|ICD9CM|HT|927.1|Crushing injury of elbow and forearm
C0160977|ICD9CM|PT|927.10|Crushing injury of forearm
C0160977|ICD9CM|AB|927.10|Crushing injury forearm
C0160978|ICD9CM|PT|927.11|Crushing injury of elbow
C0160978|ICD9CM|AB|927.11|Crushing injury elbow
C0160979|ICD9CM|HT|927.2|Crushing injury of wrist and hand(s), except finger(s) alone
C0160981|ICD9CM|AB|927.21|Crushing injury of wrist
C0160981|ICD9CM|PT|927.21|Crushing injury of wrist
C0160983|ICD9CM|PT|927.8|Crushing injury of multiple sites of upper limb
C0160983|ICD9CM|AB|927.8|Mult crushing injury arm
C0160985|ICD9CM|AB|928.9|Crushing injury leg NOS
C0160985|ICD9CM|HT|928|Crushing injury of lower limb
C0160985|ICD9CM|PT|928.9|Crushing injury of unspecified site of lower limb
C0160986|ICD9CM|HT|928.0|Crushing injury of hip and thigh
C0160987|ICD9CM|PT|928.00|Crushing injury of thigh
C0160987|ICD9CM|AB|928.00|Crushing injury thigh
C0160988|ICD9CM|PT|928.01|Crushing injury of hip
C0160988|ICD9CM|AB|928.01|Crushing injury hip
C0160989|ICD9CM|HT|928.1|Crushing injury of knee and lower leg
C0160990|ICD9CM|PT|928.10|Crushing injury of lower leg
C0160990|ICD9CM|AB|928.10|Crushing inj lower leg
C0160991|ICD9CM|PT|928.11|Crushing injury of knee
C0160991|ICD9CM|AB|928.11|Crushing injury knee
C0160992|ICD9CM|HT|928.2|Crushing injury of ankle and foot, excluding toe(s) alone
C0160993|ICD9CM|PT|928.20|Crushing injury of foot
C0160993|ICD9CM|AB|928.20|Crushing injury foot
C0160994|ICD9CM|PT|928.21|Crushing injury of ankle
C0160994|ICD9CM|AB|928.21|Crushing injury ankle
C0160996|ICD9CM|PT|928.8|Crushing injury of multiple sites of lower limb
C0160996|ICD9CM|AB|928.8|Mult crushing injury leg
C0161001|ICD9CM|HT|930|Foreign body on external eye
C0161001|ICD9CM|PT|930.9|Foreign body in unspecified site on external eye
C0161001|ICD9CM|AB|930.9|Foreign bdy ext eye NOS
C0161002|ICD9CM|AB|930.0|Corneal foreign body
C0161002|ICD9CM|PT|930.0|Corneal foreign body
C0161003|ICD9CM|PT|930.1|Foreign body in conjunctival sac
C0161003|ICD9CM|AB|930.1|FB in conjunctival sac
C0161004|ICD9CM|PT|930.2|Foreign body in lacrimal punctum
C0161004|ICD9CM|AB|930.2|FB in lacrimal punctum
C0161005|ICD9CM|PT|930.8|Foreign body in other and combined sites on external eye
C0161005|ICD9CM|AB|930.8|Foreign bdy ext eye NEC
C0161007|ICD9CM|AB|931|Foreign body in ear
C0161007|ICD9CM|PT|931|Foreign body in ear
C0161008|ICD9CM|AB|932|Foreign body in nose
C0161008|ICD9CM|PT|932|Foreign body in nose
C0161009|ICD9CM|HT|933|Foreign body in pharynx and larynx
C0161010|ICD9CM|AB|933.0|Foreign body in pharynx
C0161010|ICD9CM|PT|933.0|Foreign body in pharynx
C0161011|ICD9CM|AB|933.1|Foreign body in larynx
C0161011|ICD9CM|PT|933.1|Foreign body in larynx
C0161013|ICD9CM|AB|934.0|Foreign body in trachea
C0161013|ICD9CM|PT|934.0|Foreign body in trachea
C0161014|ICD9CM|PT|934.1|Foreign body in main bronchus
C0161014|ICD9CM|AB|934.1|Foreign body bronchus
C0161015|ICD9CM|PT|934.8|Foreign body in other specified parts bronchus and lung
C0161015|ICD9CM|AB|934.8|FB trach/bronch/lung NEC
C0161016|ICD9CM|PT|934.9|Foreign body in respiratory tree, unspecified
C0161016|ICD9CM|AB|934.9|FB respiratory tree NOS
C0161017|ICD9CM|HT|935|Foreign body in mouth, esophagus, and stomach
C0161018|ICD9CM|AB|935.0|Foreign body in mouth
C0161018|ICD9CM|PT|935.0|Foreign body in mouth
C0161019|ICD9CM|AB|935.2|Foreign body in stomach
C0161019|ICD9CM|PT|935.2|Foreign body in stomach
C0161020|ICD9CM|PT|936|Foreign body in intestine and colon
C0161020|ICD9CM|AB|936|FB in intestine & colon
C0161021|ICD9CM|PT|937|Foreign body in anus and rectum
C0161021|ICD9CM|AB|937|Foreign body anus/rectum
C0161022|ICD9CM|HT|939|Foreign body in genitourinary tract
C0161022|ICD9CM|PT|939.9|Foreign body in unspecified site in genitourinary tract
C0161022|ICD9CM|AB|939.9|Foreign bdy gu tract NOS
C0161023|ICD9CM|PT|939.0|Foreign body in bladder and urethra
C0161023|ICD9CM|AB|939.0|FB bladder & urethra
C0161025|ICD9CM|PT|939.2|Foreign body in vulva and vagina
C0161025|ICD9CM|AB|939.2|Foreign bdy vulva/vagina
C0161026|ICD9CM|PT|939.3|Foreign body in penis
C0161026|ICD9CM|AB|939.3|Foreign body penis
C0161029|ICD9CM|PT|940.1|Other burns of eyelids and periocular area
C0161029|ICD9CM|AB|940.1|Burn periocular area NEC
C0161030|ICD9CM|PT|940.2|Alkaline chemical burn of cornea and conjunctival sac
C0161030|ICD9CM|AB|940.2|Alkal burn cornea/conjun
C0161031|ICD9CM|PT|940.3|Acid chemical burn of cornea and conjunctival sac
C0161031|ICD9CM|AB|940.3|Acid burn cornea/conjunc
C0161033|ICD9CM|PT|940.5|Burn with resulting rupture and destruction of eyeball
C0161033|ICD9CM|AB|940.5|Burn w eyeball destruct
C0161036|ICD9CM|PT|941.01|Burn of unspecified degree of ear [any part]
C0161036|ICD9CM|AB|941.01|Burn NOS ear
C0161037|ICD9CM|PT|941.03|Burn of unspecified degree of lip(s)
C0161037|ICD9CM|AB|941.03|Burn NOS lip
C0161038|ICD9CM|PT|941.04|Burn of unspecified degree of chin
C0161038|ICD9CM|AB|941.04|Burn NOS chin
C0161041|ICD9CM|PT|941.07|Burn of unspecified degree of forehead and cheek
C0161041|ICD9CM|AB|941.07|Burn NOS face NEC
C0161043|ICD9CM|PT|941.09|Burn of unspecified degree of multiple sites [except with eye] of face, head, and neck
C0161043|ICD9CM|AB|941.09|Burn NOS head-mult
C0161044|ICD9CM|HT|941.1|Erythema due to burn [first degree] of face, head, and neck
C0161046|ICD9CM|PT|941.11|Erythema [first degree] of ear [any part]
C0161046|ICD9CM|AB|941.11|1st deg burn ear
C0161047|ICD9CM|PT|941.12|Erythema [first degree] of eye (with other parts face, head, and neck)
C0161047|ICD9CM|AB|941.12|1st deg burn eye
C0161048|ICD9CM|PT|941.13|Erythema [first degree] of lip(s)
C0161048|ICD9CM|AB|941.13|1st deg burn lip
C0161050|ICD9CM|PT|941.15|Erythema [first degree] of nose (septum)
C0161050|ICD9CM|AB|941.15|1st deg burn nose
C0161052|ICD9CM|PT|941.17|Erythema [first degree] of forehead and cheek
C0161052|ICD9CM|AB|941.17|1st deg burn face NEC
C0161053|ICD9CM|PT|941.18|Erythema [first degree] of neck
C0161053|ICD9CM|AB|941.18|1st deg burn neck
C0161054|ICD9CM|PT|941.19|Erythema [first degree] of multiple sites [except with eye] of face, head, and neck
C0161054|ICD9CM|AB|941.19|1st deg burn head-mult
C0161055|ICD9CM|HT|941.2|Blisters with epidermal loss due to burn [second degree] of face, head, and neck
C0161058|ICD9CM|PT|941.22|Blisters, epidermal loss [second degree] of eye (with other parts of face, head, and neck)
C0161058|ICD9CM|AB|941.22|2nd deg burn eye
C0161059|ICD9CM|PT|941.23|Blisters, epidermal loss [second degree] of lip(s)
C0161059|ICD9CM|AB|941.23|2nd deg burn lip
C0161060|ICD9CM|PT|941.24|Blisters, epidermal loss [second degree] of chin
C0161060|ICD9CM|AB|941.24|2nd deg burn chin
C0161061|ICD9CM|PT|941.25|Blisters, epidermal loss [second degree] of nose (septum)
C0161061|ICD9CM|AB|941.25|2nd deg burn nose
C0161062|ICD9CM|PT|941.26|Blisters, epidermal loss [second degree] of scalp [any part]
C0161062|ICD9CM|AB|941.26|2nd deg burn scalp
C0161063|ICD9CM|PT|941.27|Blisters, epidermal loss [second degree] of forehead and cheek
C0161063|ICD9CM|AB|941.27|2nd deg burn face NEC
C0161064|ICD9CM|PT|941.28|Blisters, epidermal loss [second degree] of neck
C0161064|ICD9CM|AB|941.28|2nd deg burn neck
C0161065|ICD9CM|PT|941.29|Blisters, epidermal loss [second degree] of multiple sites [except with eye] of face, head, and neck
C0161065|ICD9CM|AB|941.29|2nd deg burn head-mult
C0161066|ICD9CM|HT|941.3|Full-thickness skin loss due to burn [third degree NOS] of face, head, and neck
C0161067|ICD9CM|PT|941.30|Full-thickness skin loss [third degree, not otherwise specified] of face and head, unspecified site
C0161067|ICD9CM|AB|941.30|3rd deg burn head NOS
C0161068|ICD9CM|PT|941.31|Full-thickness skin loss [third degree, not otherwise specified] of ear [any part]
C0161068|ICD9CM|AB|941.31|3rd deg burn ear
C0161069|ICD9CM|PT|941.32|Full-thickness skin loss [third degree, not otherwise specified] of eye (with other parts of face, head, and neck)
C0161069|ICD9CM|AB|941.32|3rd deg burn eye
C0161070|ICD9CM|PT|941.33|Full-thickness skin loss [third degree, not otherwise specified] of lip(s)
C0161070|ICD9CM|AB|941.33|3rd deg burn lip
C0161071|ICD9CM|PT|941.34|Full-thickness skin loss [third degree, not otherwise specified] of chin
C0161071|ICD9CM|AB|941.34|3rd deg burn chin
C0161072|ICD9CM|PT|941.35|Full-thickness skin loss [third degree, not otherwise specified] of nose (septum)
C0161072|ICD9CM|AB|941.35|3rd deg burn nose
C0161073|ICD9CM|PT|941.36|Full-thickness skin loss [third degree, not otherwise specified] of scalp [any part]
C0161073|ICD9CM|AB|941.36|3rd deg burn scalp
C0161074|ICD9CM|PT|941.37|Full-thickness skin loss [third degree, not otherwise specified] of forehead and cheek
C0161074|ICD9CM|AB|941.37|3rd deg burn face NEC
C0161075|ICD9CM|PT|941.38|Full-thickness skin loss [third degree, not otherwise specified] of neck
C0161075|ICD9CM|AB|941.38|3rd deg burn neck
C0161076|ICD9CM|PT|941.39|Full-thickness skin loss [third degree, not otherwise specified] of multiple sites [except with eye] of face, head, and neck
C0161076|ICD9CM|AB|941.39|3rd deg burn head-mult
C0161077|ICD9CM|HT|941.4|Deep necrosis of underlying tissues due to burn [deep third degree] of face, head, and neck without mention of loss of a body part
C0161078|ICD9CM|PT|941.40|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, face and head, unspecified site
C0161078|ICD9CM|AB|941.40|Deep 3 deg burn head NOS
C0161079|ICD9CM|PT|941.41|Deep necrosis of underlying tissues [deep third degree]) without mention of loss of a body part, ear [any part]
C0161079|ICD9CM|AB|941.41|Deep 3rd deg burn ear
C0161080|ICD9CM|PT|941.42|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of eye (with other parts of face, head, and neck)
C0161080|ICD9CM|AB|941.42|Deep 3rd deg burn eye
C0161081|ICD9CM|PT|941.43|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of lip(s)
C0161081|ICD9CM|AB|941.43|Deep 3rd deg burn lip
C0161082|ICD9CM|PT|941.44|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of chin
C0161082|ICD9CM|AB|941.44|Deep 3rd deg burn chin
C0161083|ICD9CM|PT|941.45|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of nose (septum)
C0161083|ICD9CM|AB|941.45|Deep 3rd deg burn nose
C0161084|ICD9CM|PT|941.46|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part of scalp [any part]
C0161084|ICD9CM|AB|941.46|Deep 3rd deg burn scalp
C0161085|ICD9CM|PT|941.47|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of forehead and cheek
C0161085|ICD9CM|AB|941.47|Deep 3rd burn face NEC
C0161086|ICD9CM|PT|941.48|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of neck
C0161086|ICD9CM|AB|941.48|Deep 3rd deg burn neck
C0161087|ICD9CM|PT|941.49|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of multiple sites [except with eye] of face, head, and neck
C0161087|ICD9CM|AB|941.49|Deep 3 deg brn head-mult
C0161088|ICD9CM|HT|941.5|Deep necrosis of underlying tissues due to burn [deep third degree] of face, head, and neck with loss of a body part
C0161089|ICD9CM|PT|941.50|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of face and head, unspecified site
C0161089|ICD9CM|AB|941.50|3rd burn w loss-head NOS
C0161090|ICD9CM|PT|941.51|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of ear [any part]
C0161090|ICD9CM|AB|941.51|3rd deg burn w loss-ear
C0161091|ICD9CM|PT|941.52|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of eye (with other parts of face, head, and neck)
C0161091|ICD9CM|AB|941.52|3rd deg burn w loss-eye
C0161092|ICD9CM|PT|941.53|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of lip(s)
C0161092|ICD9CM|AB|941.53|3rd deg burn w loss-lip
C0161093|ICD9CM|PT|941.54|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of chin
C0161093|ICD9CM|AB|941.54|3rd deg burn w loss-chin
C0161094|ICD9CM|PT|941.55|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of nose (septum)
C0161094|ICD9CM|AB|941.55|3rd deg burn w loss-nose
C0161095|ICD9CM|PT|941.56|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of scalp [any part]
C0161095|ICD9CM|AB|941.56|3rd deg brn w loss-scalp
C0161096|ICD9CM|PT|941.57|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of forehead and cheek
C0161096|ICD9CM|AB|941.57|3rd burn w loss-face NEC
C0161097|ICD9CM|PT|941.58|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of neck
C0161097|ICD9CM|AB|941.58|3rd deg burn w loss-neck
C0161098|ICD9CM|PT|941.59|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of multiple sites [except with eye] of face, head, and neck
C0161098|ICD9CM|AB|941.59|3rd brn w loss-head mult
C0161099|ICD9CM|HT|942|Burn of trunk
C0161105|ICD9CM|PT|942.05|Burn of unspecified degree of genitalia
C0161105|ICD9CM|AB|942.05|Burn NOS genitalia
C0161106|ICD9CM|PT|942.09|Burn of unspecified degree of other and multiple sites of trunk
C0161106|ICD9CM|AB|942.09|Burn NOS trunk NEC
C0161107|ICD9CM|HT|942.1|Erythema due to burn [first degree] of trunk
C0161109|ICD9CM|PT|942.11|Erythema [first degree] of breast
C0161109|ICD9CM|AB|942.11|1st deg burn breast
C0161110|ICD9CM|PT|942.12|Erythema [first degree] of chest wall, excluding breast and nipple
C0161110|ICD9CM|AB|942.12|1st deg burn chest wall
C0161113|ICD9CM|PT|942.15|Erythema [first degree] of genitalia
C0161113|ICD9CM|AB|942.15|1st deg burn genitalia
C0161114|ICD9CM|PT|942.19|Erythema [first degree] of other and multiple sites of trunk
C0161114|ICD9CM|AB|942.19|1st deg burn trunk NEC
C0161118|ICD9CM|PT|942.22|Blisters, epidermal loss [second degree] of chest wall, excluding breast and nipple
C0161118|ICD9CM|AB|942.22|2nd deg burn chest wall
C0161121|ICD9CM|PT|942.25|Blisters, epidermal loss [second degree] of genitalia
C0161121|ICD9CM|AB|942.25|2nd deg burn genitalia
C0161122|ICD9CM|PT|942.29|Blisters, epidermal loss [second degree] of other and multiple sites of trunk
C0161122|ICD9CM|AB|942.29|2nd deg burn trunk NEC
C0161123|ICD9CM|HT|942.3|Full-thickness skin loss due to burn [third degree NOS] of trunk
C0161126|ICD9CM|PT|942.32|Full-thickness skin loss [third degree, not otherwise specified] of chest wall, excluding breast and nipple
C0161126|ICD9CM|AB|942.32|3rd deg burn chest wall
C0161129|ICD9CM|PT|942.35|Full-thickness skin loss [third degree, not otherwise specified] of genitalia
C0161129|ICD9CM|AB|942.35|3rd deg burn genitalia
C0161130|ICD9CM|PT|942.39|Full-thickness skin loss [third degree, not otherwise specified] of other and multiple sites of trunk
C0161130|ICD9CM|AB|942.39|3rd deg burn trunk NEC
C0161132|ICD9CM|PT|942.40|Deep necrosis of underlying tissues [deep third degree] ) without mention of loss of a body part, of trunk, unspecified site
C0161132|ICD9CM|HT|942.4|Deep necrosis of underlying tissues due to burn [deep third degree] of trunk without mention of loss of body part
C0161132|ICD9CM|AB|942.40|Deep 3rd burn trunk NOS
C0161133|ICD9CM|PT|942.41|Deep necrosis of underlying tissues [deep third degree]) without mention of loss of a body part, of breast
C0161133|ICD9CM|AB|942.41|Deep 3rd deg burn breast
C0161134|ICD9CM|PT|942.42|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of chest wall, excluding breast and nipple
C0161134|ICD9CM|AB|942.42|Deep 3rd burn chest wall
C0161138|ICD9CM|PT|942.49|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of other and multiple sites of trunk
C0161138|ICD9CM|AB|942.49|Deep 3rd burn trunk NEC
C0161139|ICD9CM|HT|942.5|Deep necrosis of underlying tissues due to burn [deep third degree] of trunk with loss of a body part
C0161140|ICD9CM|PT|942.50|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, trunk, unspecified site
C0161140|ICD9CM|AB|942.50|3rd brn w loss-trunk NOS
C0161141|ICD9CM|PT|942.51|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of breast
C0161141|ICD9CM|AB|942.51|3rd burn w loss-breast
C0161142|ICD9CM|PT|942.52|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of chest wall, excluding breast and nipple
C0161142|ICD9CM|AB|942.52|3rd brn w loss-chest wll
C0161146|ICD9CM|PT|942.59|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of other and multiple sites of trunk,
C0161146|ICD9CM|AB|942.59|3rd brn w loss-trunk NEC
C0161151|ICD9CM|PT|943.03|Burn of unspecified degree of upper arm
C0161151|ICD9CM|AB|943.03|Burn NOS upper arm
C0161155|ICD9CM|PT|943.09|Burn of unspecified degree of multiple sites of upper limb, except wrist and hand
C0161155|ICD9CM|AB|943.09|Burn NOS arm-multiple
C0161156|ICD9CM|HT|943.1|Erythema due to burn [first degree] of upper limb, except wrist and hand
C0161157|ICD9CM|PT|943.10|Erythema [first degree] of upper limb, unspecified site
C0161157|ICD9CM|AB|943.10|1st deg burn arm NOS
C0161158|ICD9CM|PT|943.11|Erythema [first degree] of forearm
C0161158|ICD9CM|AB|943.11|1st deg burn forearm
C0161159|ICD9CM|PT|943.12|Erythema [first degree] of elbow
C0161159|ICD9CM|AB|943.12|1st deg burn elbow
C0161160|ICD9CM|PT|943.13|Erythema [first degree] of upper arm
C0161160|ICD9CM|AB|943.13|1st deg burn upper arm
C0161161|ICD9CM|PT|943.14|Erythema [first degree] of axilla
C0161161|ICD9CM|AB|943.14|1st deg burn axilla
C0161162|ICD9CM|PT|943.15|Erythema [first degree] of shoulder
C0161162|ICD9CM|AB|943.15|1st deg burn shoulder
C0161163|ICD9CM|PT|943.16|Erythema [first degree] of scapular region
C0161163|ICD9CM|AB|943.16|1st deg burn scapula
C0161164|ICD9CM|PT|943.19|Erythema [first degree] of multiple sites of upper limb, except wrist and hand
C0161164|ICD9CM|AB|943.19|1st deg burn arm-mult
C0161165|ICD9CM|HT|943.2|Blisters with epidermal loss due to burn [second degree] of upper limb, except wrist and hand
C0161166|ICD9CM|PT|943.20|Blisters, epidermal loss [second degree] of upper limb, unspecified site
C0161166|ICD9CM|AB|943.20|2nd deg burn arm NOS
C0161167|ICD9CM|PT|943.21|Blisters, epidermal loss [second degree] of forearm
C0161167|ICD9CM|AB|943.21|2nd deg burn forearm
C0161168|ICD9CM|PT|943.22|Blisters, epidermal loss [second degree] of elbow
C0161168|ICD9CM|AB|943.22|2nd deg burn elbow
C0161169|ICD9CM|PT|943.23|Blisters, epidermal loss [second degree] of upper arm
C0161169|ICD9CM|AB|943.23|2nd deg burn upper arm
C0161170|ICD9CM|PT|943.24|Blisters, epidermal loss [second degree] of axilla
C0161170|ICD9CM|AB|943.24|2nd deg burn axilla
C0161171|ICD9CM|PT|943.25|Blisters, epidermal loss [second degree] of shoulder
C0161171|ICD9CM|AB|943.25|2nd deg burn shoulder
C0161172|ICD9CM|PT|943.26|Blisters, epidermal loss [second degree] of scapular region
C0161172|ICD9CM|AB|943.26|2nd deg burn scapula
C0161173|ICD9CM|PT|943.29|Blisters, epidermal loss [second degree] of multiple sites of upper limb, except wrist and hand
C0161173|ICD9CM|AB|943.29|2nd deg burn arm-mult
C0161174|ICD9CM|HT|943.3|Full-thickness skin loss due to burn [third degree NOS] of upper limb, except wrist and hand
C0161175|ICD9CM|PT|943.30|Full-thickness skin [third degree, not otherwise specified] of upper limb, unspecified site
C0161175|ICD9CM|AB|943.30|3rd deg burn arm NOS
C0161176|ICD9CM|PT|943.31|Full-thickness skin loss [third degree, not otherwise specified] of forearm
C0161176|ICD9CM|AB|943.31|3rd deg burn forearm
C0161177|ICD9CM|PT|943.32|Full-thickness skin loss [third degree, not otherwise specified] of elbow
C0161177|ICD9CM|AB|943.32|3rd deg burn elbow
C0161178|ICD9CM|PT|943.33|Full-thickness skin loss [third degree, not otherwise specified] of upper arm
C0161178|ICD9CM|AB|943.33|3rd deg burn upper arm
C0161180|ICD9CM|PT|943.35|Full-thickness skin loss [third degree, not otherwise specified] of shoulder
C0161180|ICD9CM|AB|943.35|3rd deg burn shoulder
C0161181|ICD9CM|PT|943.36|Full-thickness skin loss [third degree, not otherwise specified] of scapular region
C0161181|ICD9CM|AB|943.36|3rd deg burn scapula
C0161182|ICD9CM|PT|943.39|Full-thickness skin loss [third degree, not otherwise specified] of multiple sites of upper limb, except wrist and hand
C0161182|ICD9CM|AB|943.39|3rd deg burn arm-mult
C0161183|ICD9CM|HT|943.4|Deep necrosis of underlying tissues due to burn [deep third degree] of upper limb, except wrist and hand, without mention of loss of a body part
C0161184|ICD9CM|PT|943.40|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of upper limb,unspecified site
C0161184|ICD9CM|AB|943.40|Deep 3 deg burn arm NOS
C0161185|ICD9CM|PT|943.41|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of forearm
C0161185|ICD9CM|AB|943.41|Deep 3 deg burn forearm
C0161186|ICD9CM|PT|943.42|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of elbow
C0161186|ICD9CM|AB|943.42|Deep 3 deg burn elbow
C0161187|ICD9CM|PT|943.43|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of upper arm
C0161187|ICD9CM|AB|943.43|Deep 3 deg brn upper arm
C0161188|ICD9CM|PT|943.44|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of axilla
C0161188|ICD9CM|AB|943.44|Deep 3 deg burn axilla
C0161189|ICD9CM|PT|943.45|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of shoulder
C0161189|ICD9CM|AB|943.45|Deep 3 deg burn shoulder
C0161190|ICD9CM|PT|943.46|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of scapular region
C0161190|ICD9CM|AB|943.46|Deep 3 deg burn scapula
C0161191|ICD9CM|PT|943.49|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of multiple sites of upper limb, except wrist and hand
C0161191|ICD9CM|AB|943.49|Deep 3 deg burn arm-mult
C0161193|ICD9CM|PT|943.50|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of upper limb, unspecified site
C0161193|ICD9CM|AB|943.50|3rd burn w loss-arm NOS
C0161194|ICD9CM|PT|943.51|Deep necrosis of underlying tissues [deep third degree) with loss of a body part, of forearm
C0161194|ICD9CM|AB|943.51|3rd burn w loss-forearm
C0161195|ICD9CM|PT|943.52|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of elbow
C0161195|ICD9CM|AB|943.52|3rd burn w loss-elbow
C0161196|ICD9CM|PT|943.53|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of upper arm
C0161196|ICD9CM|AB|943.53|3rd brn w loss-upper arm
C0161197|ICD9CM|PT|943.54|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of axilla
C0161197|ICD9CM|AB|943.54|3rd burn w loss-axilla
C0161198|ICD9CM|PT|943.55|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of shoulder
C0161198|ICD9CM|AB|943.55|3rd burn w loss-shoulder
C0161199|ICD9CM|PT|943.56|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of scapular region
C0161199|ICD9CM|AB|943.56|3rd burn w loss-scapula
C0161200|ICD9CM|PT|943.59|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of multiple sites of upper limb, except wrist and hand
C0161200|ICD9CM|AB|943.59|3rd burn w loss arm-mult
C0161203|ICD9CM|PT|944.01|Burn of unspecified degree of single digit (finger (nail) other than thumb
C0161203|ICD9CM|AB|944.01|Burn NOS finger
C0161204|ICD9CM|PT|944.02|Burn of unspecified degree of thumb (nail)
C0161204|ICD9CM|AB|944.02|Burn NOS thumb
C0161205|ICD9CM|PT|944.03|Burn of unspecified degree of two or more digits of hand, not including thumb
C0161205|ICD9CM|AB|944.03|Burn NOS mult fingers
C0161206|ICD9CM|PT|944.04|Burn of unspecified degree of two or more digits of hand, including thumb
C0161206|ICD9CM|AB|944.04|Burn NOS finger w thumb
C0161207|ICD9CM|AB|944.05|Burn NOS palm
C0161207|ICD9CM|PT|944.05|Burn of unspecified degree of palm
C0161208|ICD9CM|PT|944.06|Burn of unspecified degree of back of hand
C0161208|ICD9CM|AB|944.06|Burn NOS back of hand
C0161210|ICD9CM|PT|944.08|Burn of unspecified degree of multiple sites of wrist(s) and hand(s)
C0161210|ICD9CM|AB|944.08|Burn NOS hand-multiple
C0161211|ICD9CM|HT|944.1|Erythema due to burn [first degree] of wrist(s) and hand(s)
C0161213|ICD9CM|PT|944.11|Erythema [first degree] of single digit (finger (nail)) other than thumb
C0161213|ICD9CM|AB|944.11|1st deg burn finger
C0161214|ICD9CM|PT|944.12|Erythema [first degree] of thumb (nail)
C0161214|ICD9CM|AB|944.12|1st deg burn thumb
C0161215|ICD9CM|PT|944.13|Erythema [first degree] of two or more digits of hand, not including thumb
C0161215|ICD9CM|AB|944.13|1st deg burn mult finger
C0161217|ICD9CM|PT|944.15|Erythema [first degree] of palm
C0161217|ICD9CM|AB|944.15|1st deg burn palm
C0161220|ICD9CM|PT|944.18|Erythema [first degree] of multiple sites of wrist(s) and hand(s)
C0161220|ICD9CM|AB|944.18|1st deg burn hand-mult
C0161221|ICD9CM|HT|944.2|Blisters with epidermal loss due to burn [second degree] of wrist(s) and hand(s)
C0161223|ICD9CM|PT|944.21|Blisters, epidermal loss [second degree] of single digit [finger (nail)] other than thumb
C0161223|ICD9CM|AB|944.21|2nd deg burn finger
C0161224|ICD9CM|PT|944.22|Blisters, epidermal loss [second degree] of thumb (nail)
C0161224|ICD9CM|AB|944.22|2nd deg burn thumb
C0161225|ICD9CM|PT|944.23|Blisters, epidermal loss [second degree] of two or more digits of hand, not including thumb
C0161225|ICD9CM|AB|944.23|2nd deg burn mult finger
C0161226|ICD9CM|PT|944.24|Blisters, epidermal loss [second degree] of two or more digits of hand including thumb
C0161226|ICD9CM|AB|944.24|2 deg burn fingr w thumb
C0161227|ICD9CM|PT|944.25|Blisters, epidermal loss [second degree] of palm
C0161227|ICD9CM|AB|944.25|2nd deg burn palm
C0161228|ICD9CM|PT|944.26|Blisters , epidermal loss [second degree] of back of hand
C0161228|ICD9CM|AB|944.26|2 deg burn back of hand
C0161230|ICD9CM|PT|944.28|Blisters, epidermal loss [second degree] of multiple sites of wrist(s) and hand(s)
C0161230|ICD9CM|AB|944.28|2nd deg burn hand-mult
C0161232|ICD9CM|PT|944.30|Full-thickness skin loss [third degree, not otherwise specified] of hand, unspecified site
C0161232|ICD9CM|AB|944.30|3rd deg burn hand NOS
C0161233|ICD9CM|PT|944.31|Full-thickness skin loss [third degree, not otherwise specified] of single digit [finger (nail)] other than thumb
C0161233|ICD9CM|AB|944.31|3rd deg burn finger
C0161234|ICD9CM|PT|944.32|Full-thickness skin loss [third degree, not otherwise specified] of thumb (nail)
C0161234|ICD9CM|AB|944.32|3rd deg burn thumb
C0161235|ICD9CM|PT|944.33|Full-thickness skin loss [third degree, not otherwise specified]of two or more digits of hand, not including thumb
C0161235|ICD9CM|AB|944.33|3rd deg burn mult finger
C0161236|ICD9CM|PT|944.34|Full-thickness skin loss [third degree, not otherwise specified] of two or more digits of hand including thumb
C0161236|ICD9CM|AB|944.34|3 deg burn fingr w thumb
C0161237|ICD9CM|PT|944.35|Full-thickness skin loss [third degree, not otherwise specified] of palm of hand
C0161237|ICD9CM|AB|944.35|3rd deg burn palm
C0161238|ICD9CM|PT|944.36|Full-thickness skin loss [third degree, not otherwise specified] of back of hand
C0161238|ICD9CM|AB|944.36|3 deg burn back of hand
C0161240|ICD9CM|PT|944.38|Full-thickness skin loss [third degree, not otherwise specified] of multiple sites of wrist(s) and hand(s)
C0161240|ICD9CM|AB|944.38|3rd deg burn hand-mult
C0161241|ICD9CM|HT|944.4|Deep necrosis of underlying tissues due to burn [deep third degree] of wrist(s) and hand(s), without mention of loss of a body part
C0161242|ICD9CM|PT|944.40|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, hand, unspecified site
C0161242|ICD9CM|AB|944.40|Deep 3 deg brn hand NOS
C0161243|ICD9CM|PT|944.41|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, single digit [finger (nail)] other than thumb
C0161243|ICD9CM|AB|944.41|Deep 3 deg burn finger
C0161244|ICD9CM|PT|944.42|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, thumb (nail)
C0161244|ICD9CM|AB|944.42|Deep 3 deg burn thumb
C0161245|ICD9CM|PT|944.43|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, two or more digits of hand, not including thumb
C0161245|ICD9CM|AB|944.43|Deep 3rd brn mult finger
C0161246|ICD9CM|PT|944.44|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, two or more digits of hand including thumb
C0161246|ICD9CM|AB|944.44|Deep 3rd brn fngr w thmb
C0161247|ICD9CM|PT|944.45|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of palm of hand
C0161247|ICD9CM|AB|944.45|Deep 3 deg burn palm
C0161248|ICD9CM|PT|944.46|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of back of hand
C0161248|ICD9CM|AB|944.46|Deep 3rd brn back of hnd
C0161249|ICD9CM|PT|944.47|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of wrist
C0161249|ICD9CM|AB|944.47|Deep 3 deg burn wrist
C0161250|ICD9CM|PT|944.48|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of multiple sites of wrist(s) and hand(s)
C0161250|ICD9CM|AB|944.48|Deep 3 deg brn hand-mult
C0161251|ICD9CM|HT|944.5|Deep necrosis of underlying tissues due to burn [deep third degree] of wrist(s) and hand(s), with loss of a body part
C0161252|ICD9CM|PT|944.50|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of hand, unspecified site
C0161252|ICD9CM|AB|944.50|3rd brn w loss-hand NOS
C0161253|ICD9CM|PT|944.51|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of single digit [finger (nail)] other than thumb
C0161253|ICD9CM|AB|944.51|3rd burn w loss-finger
C0161254|ICD9CM|PT|944.52|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of thumb (nail)
C0161254|ICD9CM|AB|944.52|3rd burn w loss-thumb
C0161255|ICD9CM|PT|944.53|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of two or more digits of hand, not including thumb
C0161255|ICD9CM|AB|944.53|3rd brn w loss-mult fngr
C0161256|ICD9CM|PT|944.54|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of two or more digits of hand including thumb
C0161256|ICD9CM|AB|944.54|3rd brn w loss-fngr/thmb
C0161257|ICD9CM|PT|944.55|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of palm of hand
C0161257|ICD9CM|AB|944.55|3rd burn w loss-palm
C0161258|ICD9CM|PT|944.56|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of back of hand
C0161258|ICD9CM|AB|944.56|3rd brn w loss-bk of hnd
C0161259|ICD9CM|PT|944.57|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of wrist
C0161259|ICD9CM|AB|944.57|3rd burn w loss-wrist
C0161260|ICD9CM|PT|944.58|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of multiple sites of wrist(s) and hand(s)
C0161260|ICD9CM|AB|944.58|3rd brn w loss hand-mult
C0161263|ICD9CM|PT|945.01|Burn of unspecified degree of toe(s) (nail)
C0161263|ICD9CM|AB|945.01|Burn NOS toe
C0161269|ICD9CM|PT|945.09|Burn of unspecified degree of multiple sites of lower limb(s)
C0161269|ICD9CM|AB|945.09|Burn NOS leg-multiple
C0161270|ICD9CM|HT|945.1|Erythema due to burn [first degree] of lower limb(s)
C0161271|ICD9CM|PT|945.10|Erythema [first degree] of lower limb [leg], unspecified site
C0161271|ICD9CM|AB|945.10|1st deg burn leg NOS
C0161272|ICD9CM|PT|945.11|Erythema [first degree] of toe(s) (nail)
C0161272|ICD9CM|AB|945.11|1st deg burn toe
C0161273|ICD9CM|PT|945.12|Erythema [first degree] of foot
C0161273|ICD9CM|AB|945.12|1st deg burn foot
C0161274|ICD9CM|PT|945.13|Erythema [first degree] of ankle
C0161274|ICD9CM|AB|945.13|1st deg burn ankle
C0161275|ICD9CM|PT|945.14|Erythema [first degree] of lower leg
C0161275|ICD9CM|AB|945.14|1st deg burn lower leg
C0161276|ICD9CM|PT|945.15|Erythema [first degree] of knee
C0161276|ICD9CM|AB|945.15|1st deg burn knee
C0161277|ICD9CM|PT|945.16|Erythema [first degree] of thigh [any part]
C0161277|ICD9CM|AB|945.16|1st deg burn thigh
C0161278|ICD9CM|PT|945.19|Erythema [first degree] of multiple sites of lower limb(s)
C0161278|ICD9CM|AB|945.19|1st deg burn leg-mult
C0161279|ICD9CM|HT|945.2|Blisters with epidermal loss due to burn [second degree] of lower limb(s)
C0161280|ICD9CM|PT|945.20|Blisters, epidermal loss [second degree] of lower limb [leg], unspecified site
C0161280|ICD9CM|AB|945.20|2nd deg burn leg NOS
C0161281|ICD9CM|PT|945.21|Blisters, epidermal loss [second degree] of toe(s) (nail)
C0161281|ICD9CM|AB|945.21|2nd deg burn toe
C0161282|ICD9CM|PT|945.22|Blisters, epidermal loss [second degree] of foot
C0161282|ICD9CM|AB|945.22|2nd deg burn foot
C0161283|ICD9CM|PT|945.23|Blisters, epidermal loss [second degree] of ankle
C0161283|ICD9CM|AB|945.23|2nd deg burn ankle
C0161284|ICD9CM|PT|945.24|Blisters, epidermal loss [second degree] of lower leg
C0161284|ICD9CM|AB|945.24|2nd deg burn lower leg
C0161285|ICD9CM|PT|945.25|Blisters, epidermal loss [second degree] of knee
C0161285|ICD9CM|AB|945.25|2nd deg burn knee
C0161286|ICD9CM|PT|945.26|Blisters, epidermal loss [second degree] of thigh [any part]
C0161286|ICD9CM|AB|945.26|2nd deg burn thigh
C0161287|ICD9CM|PT|945.29|Blisters, epidermal loss [second degree] of multiple sites of lower limb(s)
C0161287|ICD9CM|AB|945.29|2nd deg burn leg-mult
C0161288|ICD9CM|HT|945.3|Full-thickness skin loss due to burn [third degree NOS] of lower limb(s)
C0161289|ICD9CM|PT|945.30|Full-thickness skin loss [third degree NOS] of lower limb [leg] unspecified site
C0161289|ICD9CM|AB|945.30|3rd deg burn leg NOS
C0161290|ICD9CM|PT|945.31|Full-thickness skin loss [third degree NOS] of toe(s) (nail)
C0161290|ICD9CM|AB|945.31|3rd deg burn toe
C0161291|ICD9CM|PT|945.32|Full-thickness skin loss [third degree NOS] of foot
C0161291|ICD9CM|AB|945.32|3rd deg burn foot
C0161292|ICD9CM|PT|945.33|Full-thickness skin loss [third degree NOS] of ankle
C0161292|ICD9CM|AB|945.33|3rd deg burn ankle
C0161293|ICD9CM|PT|945.34|Full-thickness skin loss [third degree nos] of lower leg
C0161293|ICD9CM|AB|945.34|3rd deg burn low leg
C0161294|ICD9CM|PT|945.35|Full-thickness skin loss [third degree NOS] of knee
C0161294|ICD9CM|AB|945.35|3rd deg burn knee
C0161295|ICD9CM|PT|945.36|Full-thickness skin loss [third degree NOS] of thigh [any part]
C0161295|ICD9CM|AB|945.36|3rd deg burn thigh
C0161296|ICD9CM|PT|945.39|Full-thickness skin loss [third degree NOS] of multiple sites of lower limb(s)
C0161296|ICD9CM|AB|945.39|3rd deg burn leg-mult
C0161298|ICD9CM|HT|945.4|Deep necrosis of underlying tissues due to burn [deep third degree] of lower limb(s) without mention of loss of a body part
C0161298|ICD9CM|PT|945.40|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, lower limb [leg], unspecified site
C0161298|ICD9CM|AB|945.40|Deep 3rd deg brn leg NOS
C0161300|ICD9CM|PT|945.42|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of foot
C0161300|ICD9CM|AB|945.42|Deep 3rd deg burn foot
C0161301|ICD9CM|PT|945.43|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of ankle
C0161301|ICD9CM|AB|945.43|Deep 3rd deg burn ankle
C0161302|ICD9CM|PT|945.44|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of lower leg
C0161302|ICD9CM|AB|945.44|Deep 3rd deg brn low leg
C0161303|ICD9CM|PT|945.45|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of knee
C0161303|ICD9CM|AB|945.45|Deep 3rd deg burn knee
C0161304|ICD9CM|PT|945.46|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of thigh [any part]
C0161304|ICD9CM|AB|945.46|Deep 3rd deg burn thigh
C0161305|ICD9CM|PT|945.49|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of multiple sites of lower limb(s)
C0161305|ICD9CM|AB|945.49|Deep 3 deg burn leg-mult
C0161307|ICD9CM|HT|945.5|Deep necrosis of underlying tissues due to burn [deep third degree] of lower limb(s) with loss of a body part
C0161307|ICD9CM|PT|945.50|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of lower limb [leg], unspecified site
C0161307|ICD9CM|AB|945.50|3 deg brn w loss-leg NOS
C0161309|ICD9CM|PT|945.52|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of foot
C0161309|ICD9CM|AB|945.52|3 deg burn w loss-foot
C0161310|ICD9CM|PT|945.53|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of ankle
C0161310|ICD9CM|AB|945.53|3 deg burn w loss-ankle
C0161311|ICD9CM|PT|945.54|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of lower leg
C0161311|ICD9CM|AB|945.54|3 deg brn w loss-low leg
C0161312|ICD9CM|PT|945.55|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of knee
C0161312|ICD9CM|AB|945.55|3 deg burn w loss-knee
C0161313|ICD9CM|PT|945.56|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of thigh [any part]
C0161313|ICD9CM|AB|945.56|3 deg burn w loss-thigh
C0161314|ICD9CM|PT|945.59|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of multiple sites of lower limb(s)
C0161314|ICD9CM|AB|945.59|3 deg brn w loss leg-mlt
C0161316|ICD9CM|PT|946.1|Erythema [first degree] of multiple specified sites
C0161316|ICD9CM|AB|946.1|1st deg burn mult site
C0161317|ICD9CM|PT|946.2|Blisters, epidermal loss [second degree] of multiple specified sites
C0161317|ICD9CM|AB|946.2|2nd deg burn mult site
C0161318|ICD9CM|PT|946.3|Full-thickness skin loss [third degree NOS] of multiple specified sites
C0161318|ICD9CM|AB|946.3|3rd deg burn mult site
C0161319|ICD9CM|PT|946.4|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of multiple specified sites
C0161319|ICD9CM|AB|946.4|Deep 3 deg brn mult site
C0161320|ICD9CM|PT|946.5|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of multiple specified sites
C0161320|ICD9CM|AB|946.5|3rd brn w loss-mult site
C0161321|ICD9CM|PT|947.0|Burn of mouth and pharynx
C0161321|ICD9CM|AB|947.0|Burn of mouth & pharynx
C0161322|ICD9CM|PT|947.1|Burn of larynx, trachea, and lung
C0161322|ICD9CM|AB|947.1|Burn larynx/trachea/lung
C0161323|ICD9CM|PT|947.3|Burn of gastrointestinal tract
C0161323|ICD9CM|AB|947.3|Burn of GI tract
C0161325|ICD9CM|PT|947.8|Burn of other specified sites of internal organs
C0161325|ICD9CM|AB|947.8|Burn internal organ NEC
C0161327|ICD9CM|HT|948.0|Burn [any degree] involving less than 10 percent of body surface
C0161328|ICD9CM|PT|948.00|Burn [any degree] involving less than 10 percent of body surface with third degree burn, less than 10 percent or unspecified
C0161328|ICD9CM|AB|948.00|Bdy brn < 10%/3d deg NOS
C0161329|ICD9CM|HT|948.1|Burn [any degree] involving 10-19 percent of body surface
C0161330|ICD9CM|PT|948.10|Burn [any degree] involving 10-19 percent of body surface with third degree burn, less than 10 percent or unspecified
C0161330|ICD9CM|AB|948.10|10-19% bdy brn/3 deg NOS
C0161331|ICD9CM|PT|948.11|Burn [any degree] involving 10-19 percent of body surface with third degree burn, 10-19%
C0161331|ICD9CM|AB|948.11|10-19% bdy brn/10-19% 3d
C0161332|ICD9CM|HT|948.2|Burn [any degree] involving 20-29 percent of body surface
C0161333|ICD9CM|PT|948.20|Burn [any degree] involving 20-29 percent of body surface with third degree burn, less than 10 percent or unspecified
C0161333|ICD9CM|AB|948.20|20-29% bdy brn/3 deg NOS
C0161334|ICD9CM|PT|948.21|Burn [any degree] involving 20-29 percent of body surface with third degree burn, 10-19%
C0161334|ICD9CM|AB|948.21|20-29% bdy brn/10-19% 3d
C0161335|ICD9CM|PT|948.22|Burn [any degree] involving 20-29 percent of body surface with third degree burn, 20-29%
C0161335|ICD9CM|AB|948.22|20-29% bdy brn/20-29% 3d
C0161336|ICD9CM|HT|948.3|Burn [any degree] involving 30-39 percent of body surface
C0161337|ICD9CM|PT|948.30|Burn [any degree] involving 30-39 percent of body surface with third degree burn, less than 10 percent or unspecified
C0161337|ICD9CM|AB|948.30|30-39% bdy brn/3 deg NOS
C0161338|ICD9CM|PT|948.31|Burn [any degree] involving 30-39 percent of body surface with third degree burn, 10-19%
C0161338|ICD9CM|AB|948.31|30-39% bdy brn/10-19% 3d
C0161339|ICD9CM|PT|948.32|Burn [any degree] involving 30-39 percent of body surface with third degree burn, 20-29%
C0161339|ICD9CM|AB|948.32|30-39% bdy brn/20-29% 3d
C0161340|ICD9CM|PT|948.33|Burn [any degree] involving 30-39 percent of body surface with third degree burn, 30-39%
C0161340|ICD9CM|AB|948.33|30-39% bdy brn/30-39% 3d
C0161341|ICD9CM|HT|948.4|Burn [any degree] involving 40-49 percent of body surface
C0161342|ICD9CM|PT|948.40|Burn [any degree] involving 40-49 percent of body surface with third degree burn, less than 10 percent or unspecified
C0161342|ICD9CM|AB|948.40|40-49% bdy brn/3 deg NOS
C0161343|ICD9CM|PT|948.41|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 10-19%
C0161343|ICD9CM|AB|948.41|40-49% bdy brn/10-19% 3d
C0161344|ICD9CM|PT|948.42|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 20-29%
C0161344|ICD9CM|AB|948.42|40-49% bdy brn/20-29% 3d
C0161345|ICD9CM|PT|948.43|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 30-39%
C0161345|ICD9CM|AB|948.43|40-49% bdy brn/30-39% 3d
C0161346|ICD9CM|PT|948.44|Burn [any degree] involving 40-49 percent of body surface with third degree burn, 40-49%
C0161346|ICD9CM|AB|948.44|40-49% bdy brn/40-49% 3d
C0161347|ICD9CM|HT|948.5|Burn [any degree] involving 50-59 percent of body surface
C0161348|ICD9CM|PT|948.50|Burn [any degree] involving 50-59 percent of body surface with third degree burn, less than 10 percent or unspecified
C0161348|ICD9CM|AB|948.50|50-59% bdy brn/3 deg NOS
C0161349|ICD9CM|PT|948.51|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 10-19%
C0161349|ICD9CM|AB|948.51|50-59% bdy brn/10-19% 3d
C0161350|ICD9CM|PT|948.52|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 20-29%
C0161350|ICD9CM|AB|948.52|50-59% bdy brn/20-29% 3d
C0161351|ICD9CM|PT|948.53|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 30-39%
C0161351|ICD9CM|AB|948.53|50-59% bdy brn/30-39% 3d
C0161352|ICD9CM|PT|948.54|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 40-49%
C0161352|ICD9CM|AB|948.54|50-59% bdy brn/40-49% 3d
C0161353|ICD9CM|PT|948.55|Burn [any degree] involving 50-59 percent of body surface with third degree burn, 50-59%
C0161353|ICD9CM|AB|948.55|50-59% bdy brn/50-59% 3d
C0161354|ICD9CM|HT|948.6|Burn [any degree] involving 60-69 percent of body surface
C0161355|ICD9CM|PT|948.60|Burn [any degree] involving 60-69 percent of body surface with third degree burn, less than 10 percent or unspecified
C0161355|ICD9CM|AB|948.60|60-69% bdy brn/3 deg NOS
C0161356|ICD9CM|PT|948.61|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 10-19%
C0161356|ICD9CM|AB|948.61|60-69% bdy brn/10-19% 3d
C0161357|ICD9CM|PT|948.62|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 20-29%
C0161357|ICD9CM|AB|948.62|60-69% bdy brn/20-29% 3d
C0161358|ICD9CM|PT|948.63|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 30-39%
C0161358|ICD9CM|AB|948.63|60-69% bdy brn/30-39% 3d
C0161359|ICD9CM|PT|948.64|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 40-49%
C0161359|ICD9CM|AB|948.64|60-69% bdy brn/40-49% 3d
C0161360|ICD9CM|PT|948.65|Burn (any degree) involving 60-69 percent of body surface with third degree burn, 50-59%
C0161360|ICD9CM|AB|948.65|60-69% bdy brn/50-59% 3d
C0161361|ICD9CM|PT|948.66|Burn [any degree] involving 60-69 percent of body surface with third degree burn, 60-69%
C0161361|ICD9CM|AB|948.66|60-69% bdy brn/60-69% 3d
C0161362|ICD9CM|HT|948.7|Burn [any degree] involving 70-79 percent of body surface
C0161363|ICD9CM|PT|948.70|Burn [any degree] involving 70-79 percent of body surface with third degree burn, less than 10 percent or unspecified
C0161363|ICD9CM|AB|948.70|70-79% bdy brn/3 deg NOS
C0161364|ICD9CM|PT|948.71|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 10-19%
C0161364|ICD9CM|AB|948.71|70-79% bdy brn/10-19% 3d
C0161365|ICD9CM|PT|948.72|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 20-29%
C0161365|ICD9CM|AB|948.72|70-79% bdy brn/20-29% 3d
C0161366|ICD9CM|PT|948.73|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 30-39%
C0161366|ICD9CM|AB|948.73|70-79% bdy brn/30-39% 3d
C0161367|ICD9CM|PT|948.74|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 40-49%
C0161367|ICD9CM|AB|948.74|70-79% bdy brn/40-49% 3d
C0161368|ICD9CM|PT|948.75|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 50-59%
C0161368|ICD9CM|AB|948.75|70-79% bdy brn/50-59% 3d
C0161369|ICD9CM|PT|948.76|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 60-69%
C0161369|ICD9CM|AB|948.76|70-79% bdy brn/60-69% 3d
C0161370|ICD9CM|PT|948.77|Burn [any degree] involving 70-79 percent of body surface with third degree burn, 70-79%
C0161370|ICD9CM|AB|948.77|70-79% bdy brn/70-79% 3d
C0161371|ICD9CM|HT|948.8|Burn [any degree] involving 80-89 percent of body surface
C0161372|ICD9CM|PT|948.80|Burn [any degree] involving 80-89 percent of body surface with third degree burn, less than 10 percent or unspecified
C0161372|ICD9CM|AB|948.80|80-89% bdy brn/3 deg NOS
C0161373|ICD9CM|PT|948.81|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 10-19%
C0161373|ICD9CM|AB|948.81|80-89% bdy brn/10-19% 3d
C0161374|ICD9CM|PT|948.82|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 20-29%
C0161374|ICD9CM|AB|948.82|80-89% bdy brn/20-29% 3d
C0161375|ICD9CM|PT|948.83|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 30-39%
C0161375|ICD9CM|AB|948.83|80-89% bdy brn/30-39% 3d
C0161376|ICD9CM|PT|948.84|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 40-49%
C0161376|ICD9CM|AB|948.84|80-89% bdy brn/40-49% 3d
C0161377|ICD9CM|PT|948.85|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 50-59%
C0161377|ICD9CM|AB|948.85|80-89% bdy brn/50-59% 3d
C0161378|ICD9CM|PT|948.86|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 60-69%
C0161378|ICD9CM|AB|948.86|80-89% bdy brn/60-69% 3d
C0161379|ICD9CM|PT|948.87|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 70-79%
C0161379|ICD9CM|AB|948.87|80-89% bdy brn/70-79% 3d
C0161380|ICD9CM|PT|948.88|Burn [any degree] involving 80-89 percent of body surface with third degree burn, 80-89%
C0161380|ICD9CM|AB|948.88|80-89% bdy brn/80-89% 3d
C0161381|ICD9CM|HT|948.9|Burn [any degree] involving 90 percent or more of body surface
C0161382|ICD9CM|PT|948.90|Burn [any degree] involving 90 percent or more of body surface with third degree burn, less than 10 percent or unspecified
C0161382|ICD9CM|AB|948.90|90% + bdy brn/3d deg NOS
C0161383|ICD9CM|PT|948.91|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 10-19%
C0161383|ICD9CM|AB|948.91|90% + bdy brn/10-19% 3rd
C0161384|ICD9CM|PT|948.92|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 20-29%
C0161384|ICD9CM|AB|948.92|90% + bdy brn/20-29% 3rd
C0161385|ICD9CM|PT|948.93|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 30-39%
C0161385|ICD9CM|AB|948.93|90% + bdy brn/30-39% 3rd
C0161386|ICD9CM|PT|948.94|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 40-49%
C0161386|ICD9CM|AB|948.94|90% + bdy brn/40-49% 3rd
C0161387|ICD9CM|PT|948.95|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 50-59%
C0161387|ICD9CM|AB|948.95|90% + bdy brn/50-59% 3rd
C0161388|ICD9CM|PT|948.96|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 60-69%
C0161388|ICD9CM|AB|948.96|90% + bdy brn/60-69% 3rd
C0161389|ICD9CM|PT|948.97|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 70-79%
C0161389|ICD9CM|AB|948.97|90% + bdy brn/70-79% 3rd
C0161390|ICD9CM|PT|948.98|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 80-89%
C0161390|ICD9CM|AB|948.98|90% + bdy brn/80-89% 3rd
C0161391|ICD9CM|PT|948.99|Burn [any degree] involving 90 percent or more of body surface with third degree burn, 90% or more of body surface
C0161391|ICD9CM|AB|948.99|90% + bdy brn/90% + 3rd
C0161395|ICD9CM|PT|949.4|Deep necrosis of underlying tissue [deep third degree] without mention of loss of a body part, unspecified
C0161395|ICD9CM|AB|949.4|Deep 3rd deg burn NOS
C0161396|ICD9CM|PT|949.5|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, unspecified
C0161396|ICD9CM|AB|949.5|3rd burn w loss-site NOS
C0161397|ICD9CM|HT|950|Injury to optic nerve and pathways
C0161397|ICD9CM|PT|950.9|Injury to unspecified optic nerve and pathways
C0161397|ICD9CM|AB|950.9|Inj optic nerv/path NOS
C0161398|ICD9CM|AB|950.0|Optic nerve injury
C0161398|ICD9CM|PT|950.0|Optic nerve injury
C0161399|ICD9CM|AB|950.1|Injury to optic chiasm
C0161399|ICD9CM|PT|950.1|Injury to optic chiasm
C0161400|ICD9CM|AB|950.2|Injury to optic pathways
C0161400|ICD9CM|PT|950.2|Injury to optic pathways
C0161401|ICD9CM|AB|950.3|Injury to visual cortex
C0161401|ICD9CM|PT|950.3|Injury to visual cortex
C0161405|ICD9CM|PT|951.1|Injury to trochlear nerve
C0161405|ICD9CM|AB|951.1|Injury trochlear nerve
C0161406|ICD9CM|PT|951.2|Injury to trigeminal nerve
C0161406|ICD9CM|AB|951.2|Injury trigeminal nerve
C0161407|ICD9CM|AB|951.3|Injury abducens nerve
C0161407|ICD9CM|PT|951.3|Injury to abducens nerve
C0161408|ICD9CM|AB|951.4|Injury to facial nerve
C0161408|ICD9CM|PT|951.4|Injury to facial nerve
C0161409|ICD9CM|AB|951.5|Injury to acoustic nerve
C0161409|ICD9CM|PT|951.5|Injury to acoustic nerve
C0161410|ICD9CM|PT|951.6|Injury to accessory nerve
C0161410|ICD9CM|AB|951.6|Injury accessory nerve
C0161411|ICD9CM|PT|951.7|Injury to hypoglossal nerve
C0161411|ICD9CM|AB|951.7|Injury hypoglossal nerve
C0161412|ICD9CM|PT|951.8|Injury to other specified cranial nerves
C0161412|ICD9CM|AB|951.8|Injury cranial nerve NEC
C0161414|ICD9CM|HT|952|Spinal cord injury without evidence of spinal bone injury
C0161416|ICD9CM|PT|952.00|C1-C4 level with unspecified spinal cord injury
C0161416|ICD9CM|AB|952.00|C1-c4 spin cord inj NOS
C0161417|ICD9CM|PT|952.01|C1-C4 level with complete lesion of spinal cord
C0161417|ICD9CM|AB|952.01|Complete les cord/c1-c4
C0161418|ICD9CM|PT|952.02|C1-C4 level with anterior cord syndrome
C0161418|ICD9CM|AB|952.02|Anterior cord synd/c1-c4
C0161419|ICD9CM|PT|952.03|C1-C4 level with central cord syndrome
C0161419|ICD9CM|AB|952.03|Central cord synd/c1-c4
C0161420|ICD9CM|PT|952.04|C1-C4 level with other specified spinal cord injury
C0161420|ICD9CM|AB|952.04|C1-c4 spin cord inj NEC
C0161421|ICD9CM|PT|952.05|C5-C7 level with unspecified spinal cord injury
C0161421|ICD9CM|AB|952.05|C5-c7 spin cord inj NOS
C0161422|ICD9CM|PT|952.06|C5-C7 level with complete lesion of spinal cord
C0161422|ICD9CM|AB|952.06|Complete les cord/c5-c7
C0161423|ICD9CM|PT|952.07|C5-C7 level with anterior cord syndrome
C0161423|ICD9CM|AB|952.07|Anterior cord synd/c5-c7
C0161424|ICD9CM|PT|952.08|C5-C7 level with central cord syndrome
C0161424|ICD9CM|AB|952.08|Central cord synd/c5-c7
C0161425|ICD9CM|PT|952.09|C5-C7 level with other specified spinal cord injury
C0161425|ICD9CM|AB|952.09|C5-c7 spin cord inj NEC
C0161426|ICD9CM|HT|952.1|Dorsal [thoracic] spinal cord injury without evidence of spinal bone injury
C0161427|ICD9CM|PT|952.10|T1-T6 level with unspecified spinal cord injury
C0161427|ICD9CM|AB|952.10|T1-t6 spin cord inj NOS
C0161432|ICD9CM|PT|952.15|T7-T12 level with unspecified spinal cord injury
C0161432|ICD9CM|AB|952.15|T7-t12 spin cord inj NOS
C0161436|ICD9CM|PT|952.19|T7-T12 level with other specified spinal cord injury
C0161436|ICD9CM|AB|952.19|T7-t12 spin cord inj NEC
C0161439|ICD9CM|AB|952.4|Cauda equina injury
C0161439|ICD9CM|PT|952.4|Cauda equina spinal cord injury without evidence of spinal bone injury
C0161440|ICD9CM|PT|952.8|Multiple sites of spinal cord injury without evidence of spinal bone injury
C0161440|ICD9CM|AB|952.8|Spin cord inj-mult site
C0161441|ICD9CM|PT|953.9|Injury to unspecified site of nerve roots and spinal plexus
C0161441|ICD9CM|HT|953|Injury to nerve roots and spinal plexus
C0161441|ICD9CM|AB|953.9|Inj nerve root/plex NOS
C0161442|ICD9CM|PT|953.0|Injury to cervical nerve root
C0161442|ICD9CM|AB|953.0|Cervical root injury
C0161444|ICD9CM|PT|953.2|Injury to lumbar nerve root
C0161444|ICD9CM|AB|953.2|Lumbar root injury
C0161445|ICD9CM|PT|953.3|Injury to sacral nerve root
C0161445|ICD9CM|AB|953.3|Sacral root injury
C0161446|ICD9CM|PT|953.4|Injury to brachial plexus
C0161446|ICD9CM|AB|953.4|Brachial plexus injury
C0161447|ICD9CM|PT|953.5|Injury to lumbosacral plexus
C0161447|ICD9CM|AB|953.5|Lumbosacral plex injury
C0161448|ICD9CM|PT|953.8|Injury to multiple sites of nerve roots and spinal plexus
C0161448|ICD9CM|AB|953.8|Mult nerve root/plex inj
C0161451|ICD9CM|PT|954.0|Injury to cervical sympathetic nerve, excluding shoulder and pelvic girdles
C0161451|ICD9CM|AB|954.0|Inj cerv sympath nerve
C0161452|ICD9CM|PT|954.1|Injury to other sympathetic nerve, excluding shoulder and pelvic girdles
C0161452|ICD9CM|AB|954.1|Inj sympath nerve NEC
C0161453|ICD9CM|PT|954.8|Injury to other specified nerve(s) of trunk, excluding shoulder and pelvic girdles
C0161453|ICD9CM|AB|954.8|Injury trunk nerve NEC
C0161454|ICD9CM|PT|954.9|Injury to unspecified nerve of trunk, excluding shoulder and pelvic girdles
C0161454|ICD9CM|AB|954.9|Injury trunk nerve NOS
C0161456|ICD9CM|PT|955.0|Injury to axillary nerve
C0161456|ICD9CM|AB|955.0|Injury axillary nerve
C0161457|ICD9CM|PT|955.1|Injury to median nerve
C0161457|ICD9CM|AB|955.1|Injury median nerve
C0161458|ICD9CM|PT|955.2|Injury to ulnar nerve
C0161458|ICD9CM|AB|955.2|Injury ulnar nerve
C0161459|ICD9CM|PT|955.3|Injury to radial nerve
C0161459|ICD9CM|AB|955.3|Injury radial nerve
C0161460|ICD9CM|PT|955.4|Injury to musculocutaneous nerve
C0161460|ICD9CM|AB|955.4|Inj musculocutan nerve
C0161461|ICD9CM|PT|955.5|Injury to cutaneous sensory nerve, upper limb
C0161461|ICD9CM|AB|955.5|Inj cutan senso nerv/arm
C0161462|ICD9CM|PT|955.6|Injury to digital nerve, upper limb
C0161462|ICD9CM|AB|955.6|Injury digital nerve
C0161463|ICD9CM|PT|955.7|Injury to other specified nerve(s) of shoulder girdle and upper limb
C0161463|ICD9CM|AB|955.7|Inj nerve shldr/arm NEC
C0161467|ICD9CM|PT|956.0|Injury to sciatic nerve
C0161467|ICD9CM|AB|956.0|Injury sciatic nerve
C0161468|ICD9CM|PT|956.1|Injury to femoral nerve
C0161468|ICD9CM|AB|956.1|Injury femoral nerve
C0161471|ICD9CM|PT|956.4|Injury to cutaneous sensory nerve, lower limb
C0161471|ICD9CM|AB|956.4|Inj cutan senso nerv/leg
C0161473|ICD9CM|PT|956.8|Injury to multiple nerves of pelvic girdle and lower limb
C0161473|ICD9CM|AB|956.8|Inj mult nerve pelv/leg
C0161475|ICD9CM|HT|957|Injury to other and unspecified nerves
C0161476|ICD9CM|PT|957.0|Injury to superficial nerves of head and neck
C0161476|ICD9CM|AB|957.0|Inj superf nerv head/nck
C0161478|ICD9CM|PT|957.8|Injury to multiple nerves in several parts
C0161478|ICD9CM|AB|957.8|Injury to mult nerves
C0161479|ICD9CM|AB|957.9|Injury to nerve NOS
C0161479|ICD9CM|PT|957.9|Injury to nerves, unspecified site
C0161480|ICD9CM|HT|958|Certain early complications of trauma
C0161483|ICD9CM|PT|959.2|Shoulder and upper arm injury
C0161483|ICD9CM|AB|959.2|Shldr/upper arm inj NOS
C0161484|ICD9CM|PT|959.6|Hip and thigh injury
C0161484|ICD9CM|AB|959.6|Hip & thigh injury NOS
C0161485|ICD9CM|HT|960|Poisoning by antibiotics
C0161485|ICD9CM|AB|960.9|Poisoning-antibiotic NOS
C0161485|ICD9CM|PT|960.9|Poisoning by unspecified antibiotic
C0161486|ICD9CM|PT|960.0|Poisoning by penicillins
C0161486|ICD9CM|AB|960.0|Poisoning-penicillins
C0161487|ICD9CM|PT|960.1|Poisoning by antifungal antibiotics
C0161487|ICD9CM|AB|960.1|Pois-antifungal antibiot
C0161488|ICD9CM|PT|960.2|Poisoning by chloramphenicol group
C0161488|ICD9CM|AB|960.2|Poison-chloramphenicol
C0161489|ICD9CM|PT|960.3|Poisoning by erythromycin and other macrolides
C0161489|ICD9CM|AB|960.3|Pois-erythromyc/macrolid
C0161493|ICD9CM|PT|960.7|Poisoning by antineoplastic antibiotics
C0161493|ICD9CM|AB|960.7|Pois-antineop antibiotic
C0161494|ICD9CM|PT|960.8|Poisoning by other specified antibiotics
C0161494|ICD9CM|AB|960.8|Poisoning-antibiotic NEC
C0161496|ICD9CM|HT|961|Poisoning by other anti-infectives
C0161497|ICD9CM|PT|961.0|Poisoning by sulfonamides
C0161497|ICD9CM|AB|961.0|Poisoning-sulfonamides
C0161498|ICD9CM|PT|961.1|Poisoning by arsenical anti-infectives
C0161498|ICD9CM|AB|961.1|Pois-arsenic anti-infec
C0161499|ICD9CM|PT|961.2|Poisoning by heavy metal anti-infectives
C0161499|ICD9CM|AB|961.2|Pois-heav met anti-infec
C0161501|ICD9CM|PT|961.4|Poisoning by antimalarials and drugs acting on other blood protozoa
C0161501|ICD9CM|AB|961.4|Poisoning-antimalarials
C0161502|ICD9CM|PT|961.5|Poisoning by other antiprotozoal drugs
C0161502|ICD9CM|AB|961.5|Pois-antiprotoz drug NEC
C0161504|ICD9CM|PT|961.7|Poisoning by antiviral drugs
C0161504|ICD9CM|AB|961.7|Poisoning-antiviral drug
C0161505|ICD9CM|PT|961.8|Poisoning by other antimycobacterial drugs
C0161505|ICD9CM|AB|961.8|Pois-antimycobac drg NEC
C0161506|ICD9CM|PT|961.9|Poisoning by other and unspecified anti-infectives
C0161506|ICD9CM|AB|961.9|Pois-anti-infect NEC/NOS
C0161508|ICD9CM|PT|962.0|Poisoning by adrenal cortical steroids
C0161508|ICD9CM|AB|962.0|Pois-corticosteroids
C0161509|ICD9CM|PT|962.1|Poisoning by androgens and anabolic congeners
C0161509|ICD9CM|AB|962.1|Poisoning-androgens
C0161512|ICD9CM|PT|962.4|Poisoning by anterior pituitary hormones
C0161512|ICD9CM|AB|962.4|Pois-ant pituitary horm
C0161513|ICD9CM|PT|962.5|Poisoning by posterior pituitary hormones
C0161513|ICD9CM|AB|962.5|Pois-post pituitary horm
C0161514|ICD9CM|PT|962.6|Poisoning by parathyroid and parathyroid derivatives
C0161514|ICD9CM|AB|962.6|Poisoning-parathyroids
C0161515|ICD9CM|PT|962.7|Poisoning by thyroid and thyroid derivatives
C0161515|ICD9CM|AB|962.7|Poisoning-thyroid/deriv
C0161516|ICD9CM|PT|962.8|Poisoning by antithyroid agents
C0161516|ICD9CM|AB|962.8|Poison-antithyroid agent
C0161517|ICD9CM|PT|962.9|Poisoning by other and unspecified hormones and synthetic substitutes
C0161517|ICD9CM|AB|962.9|Poisoning hormon NEC/NOS
C0161518|ICD9CM|PT|963.9|Poisoning by unspecified systemic agent
C0161518|ICD9CM|HT|963|Poisoning by primarily systemic agents
C0161518|ICD9CM|AB|963.9|Poisoning-system agt NOS
C0161519|ICD9CM|PT|963.0|Poisoning by antiallergic and antiemetic drugs
C0161519|ICD9CM|AB|963.0|Pois-antiallrg/antiemet
C0161521|ICD9CM|PT|963.2|Poisoning by acidifying agents
C0161521|ICD9CM|AB|963.2|Poisoning-acidifying agt
C0161522|ICD9CM|PT|963.3|Poisoning by alkalizing agents
C0161522|ICD9CM|AB|963.3|Poisoning-alkalizing agt
C0161525|ICD9CM|PT|963.8|Poisoning by other specified systemic agents
C0161525|ICD9CM|AB|963.8|Poisoning-system agt NEC
C0161527|ICD9CM|HT|964|Poisoning by agents primarily affecting blood constituents
C0161529|ICD9CM|PT|964.1|Poisoning by liver preparations and other antianemic agents
C0161529|ICD9CM|AB|964.1|Poison-liver/antianemics
C0161530|ICD9CM|PT|964.2|Poisoning by anticoagulants
C0161530|ICD9CM|AB|964.2|Poisoning-anticoagulants
C0161533|ICD9CM|PT|964.5|Poisoning by anticoagulant antagonists and other coagulants
C0161533|ICD9CM|AB|964.5|Poisoning-coagulants
C0161534|ICD9CM|PT|964.6|Poisoning by gamma globulin
C0161534|ICD9CM|AB|964.6|Poisoning-gamma globulin
C0161536|ICD9CM|PT|964.8|Poisoning by other specified agents affecting blood constituents
C0161536|ICD9CM|AB|964.8|Poisoning-blood agt NEC
C0161537|ICD9CM|PT|964.9|Poisoning by unspecified agent affecting blood constituents
C0161537|ICD9CM|AB|964.9|Poisoning-blood agt NOS
C0161538|ICD9CM|HT|965|Poisoning by analgesics, antipyretics, and antirheumatics
C0161540|ICD9CM|PT|965.00|Poisoning by opium (alkaloids), unspecified
C0161540|ICD9CM|AB|965.00|Poisoning-opium NOS
C0161541|ICD9CM|PT|965.01|Poisoning by heroin
C0161541|ICD9CM|AB|965.01|Poisoning-heroin
C0161542|ICD9CM|PT|965.02|Poisoning by methadone
C0161542|ICD9CM|AB|965.02|Poisoning-methadone
C0161543|ICD9CM|PT|965.09|Poisoning by other opiates and related narcotics
C0161543|ICD9CM|AB|965.09|Poisoning-opiates NEC
C0161544|ICD9CM|PT|965.1|Poisoning by salicylates
C0161544|ICD9CM|AB|965.1|Poisoning-salicylates
C0161546|ICD9CM|PT|965.5|Poisoning by pyrazole derivatives
C0161546|ICD9CM|AB|965.5|Poisoning-pyrazole deriv
C0161548|ICD9CM|PT|965.7|Poisoning by other non-narcotic analgesics
C0161548|ICD9CM|AB|965.7|Pois-no-narc analges NEC
C0161549|ICD9CM|PT|965.8|Poisoning by other specified analgesics and antipyretics
C0161549|ICD9CM|AB|965.8|Pois-analges/antipyr NEC
C0161552|ICD9CM|PT|966.0|Poisoning by oxazolidine derivatives
C0161552|ICD9CM|AB|966.0|Poison-oxazolidine deriv
C0161553|ICD9CM|PT|966.1|Poisoning by hydantoin derivatives
C0161553|ICD9CM|AB|966.1|Poison-hydantoin derivat
C0161554|ICD9CM|PT|966.2|Poisoning by succinimides
C0161554|ICD9CM|AB|966.2|Poisoning-succinimides
C0161555|ICD9CM|PT|966.3|Poisoning by other and unspecified anticonvulsants
C0161555|ICD9CM|AB|966.3|Pois-anticonvul NEC/NOS
C0161556|ICD9CM|PT|966.4|Poisoning by anti-Parkinsonism drugs
C0161556|ICD9CM|AB|966.4|Pois-anti-parkinson drug
C0161558|ICD9CM|PT|967.0|Poisoning by barbiturates
C0161558|ICD9CM|AB|967.0|Poisoning-barbiturates
C0161560|ICD9CM|PT|967.2|Poisoning by paraldehyde
C0161560|ICD9CM|AB|967.2|Poisoning-paraldehyde
C0161562|ICD9CM|PT|967.4|Poisoning by methaqualone compounds
C0161562|ICD9CM|AB|967.4|Poisoning-methaqualone
C0161563|ICD9CM|PT|967.5|Poisoning by glutethimide group
C0161563|ICD9CM|AB|967.5|Poisoning-glutethimide
C0161565|ICD9CM|PT|967.8|Poisoning by other sedatives and hypnotics
C0161565|ICD9CM|AB|967.8|Pois-sedative/hypnot NEC
C0161567|ICD9CM|HT|968|Poisoning by other central nervous system depressants and anesthetics
C0161568|ICD9CM|PT|968.0|Poisoning by central nervous system muscle-tone depressants
C0161568|ICD9CM|AB|968.0|Pois-cns muscle depress
C0161569|ICD9CM|PT|968.1|Poisoning by halothane
C0161569|ICD9CM|AB|968.1|Poisoning-halothane
C0161571|ICD9CM|PT|968.3|Poisoning by intravenous anesthetics
C0161571|ICD9CM|AB|968.3|Poison-intraven anesthet
C0161572|ICD9CM|PT|968.4|Poisoning by other and unspecified general anesthetics
C0161572|ICD9CM|AB|968.4|Pois-gen anesth NEC/NOS
C0161573|ICD9CM|PT|968.5|Surface (topical) and infiltration anesthetics
C0161573|ICD9CM|AB|968.5|Surfce-topic/infilt anes
C0161574|ICD9CM|PT|968.6|Poisoning by peripheral nerve- and plexus-blocking anesthetics
C0161574|ICD9CM|AB|968.6|Pois-nerve/plex-blk anes
C0161575|ICD9CM|PT|968.7|Poisoning by spinal anesthetics
C0161575|ICD9CM|AB|968.7|Poison-spinal anesthetic
C0161576|ICD9CM|PT|968.9|Poisoning by other and unspecified local anesthetics
C0161576|ICD9CM|AB|968.9|Pois-local anest NEC/NOS
C0161577|ICD9CM|HT|969|Poisoning by psychotropic agents
C0161577|ICD9CM|PT|969.9|Poisoning by unspecified psychotropic agent
C0161577|ICD9CM|AB|969.9|Poison-psychotropic NOS
C0161578|ICD9CM|HT|969.0|Poisoning by antidepressants
C0161581|ICD9CM|PT|969.3|Poisoning by other antipsychotics, neuroleptics, and major tranquilizers
C0161581|ICD9CM|AB|969.3|Poison-antipsychotic NEC
C0161583|ICD9CM|PT|969.5|Poisoning by other tranquilizers
C0161583|ICD9CM|AB|969.5|Poison-tranquilizer NEC
C0161584|ICD9CM|PT|969.6|Poisoning by psychodysleptics (hallucinogens)
C0161584|ICD9CM|AB|969.6|Poisoning-hallucinogens
C0161585|ICD9CM|HT|969.7|Poisoning by psychostimulants
C0161586|ICD9CM|PT|969.8|Poisoning by other specified psychotropic agents
C0161586|ICD9CM|AB|969.8|Poison-psychotropic NEC
C0161588|ICD9CM|HT|970|Poisoning by central nervous system stimulants
C0161588|ICD9CM|PT|970.9|Poisoning by unspecified central nervous system stimulant
C0161588|ICD9CM|AB|970.9|Pois-cns stimulant NOS
C0161589|ICD9CM|PT|970.0|Poisoning by analeptics
C0161589|ICD9CM|AB|970.0|Poisoning-analeptics
C0161590|ICD9CM|PT|970.1|Poisoning by opiate antagonists
C0161590|ICD9CM|AB|970.1|Poison-opiate antagonist
C0161591|ICD9CM|HT|970.8|Poisoning by other specified central nervous system stimulants
C0161593|ICD9CM|HT|971|Poisoning by drugs primarily affecting the autonomic nervous system
C0161598|ICD9CM|PT|971.9|Poisoning by unspecified drug primarily affecting autonomic nervous system
C0161598|ICD9CM|AB|971.9|Pois-autonomic agent NOS
C0161599|ICD9CM|HT|972|Poisoning by agents primarily affecting the cardiovascular system
C0161601|ICD9CM|PT|972.1|Poisoning by cardiotonic glycosides and drugs of similar action
C0161601|ICD9CM|AB|972.1|Poisoning-cardiotonics
C0161602|ICD9CM|PT|972.2|Poisoning by antilipemic and antiarteriosclerotic drugs
C0161602|ICD9CM|AB|972.2|Poisoning-antilipemics
C0161603|ICD9CM|PT|972.3|Poisoning by ganglion-blocking agents
C0161603|ICD9CM|AB|972.3|Pois-ganglion block agt
C0161604|ICD9CM|PT|972.4|Poisoning by coronary vasodilators
C0161604|ICD9CM|AB|972.4|Pois-coronary vasodilat
C0161605|ICD9CM|PT|972.5|Poisoning by other vasodilators
C0161605|ICD9CM|AB|972.5|Poison-vasodilator NEC
C0161606|ICD9CM|PT|972.6|Poisoning by other antihypertensive agents
C0161606|ICD9CM|AB|972.6|Pois-antihyperten agent
C0161607|ICD9CM|PT|972.7|Poisoning by antivaricose drugs, including sclerosing agents
C0161607|ICD9CM|AB|972.7|Poison-antivaricose drug
C0161608|ICD9CM|PT|972.8|Poisoning by capillary-active drugs
C0161608|ICD9CM|AB|972.8|Poison-capillary act agt
C0161609|ICD9CM|PT|972.9|Poisoning by other and unspecified agents primarily affecting the cardiovascular system
C0161609|ICD9CM|AB|972.9|Pois-cardiovasc agt NEC
C0161610|ICD9CM|HT|973|Poisoning by agents primarily affecting the gastrointestinal system
C0161611|ICD9CM|PT|973.0|Poisoning by antacids and antigastric secretion drugs
C0161611|ICD9CM|AB|973.0|Pois-antacid/antigastric
C0161612|ICD9CM|PT|973.1|Poisoning by irritant cathartics
C0161612|ICD9CM|AB|973.1|Pois-irritant cathartics
C0161613|ICD9CM|PT|973.2|Poisoning by emollient cathartics
C0161613|ICD9CM|AB|973.2|Pois-emollient cathartic
C0161615|ICD9CM|PT|973.4|Poisoning by digestants
C0161615|ICD9CM|AB|973.4|Poisoning-digestants
C0161616|ICD9CM|PT|973.5|Poisoning by antidiarrheal drugs
C0161616|ICD9CM|AB|973.5|Poisoning-antidiarrh agt
C0161617|ICD9CM|PT|973.6|Poisoning by emetics
C0161617|ICD9CM|AB|973.6|Poisoning-emetics
C0161618|ICD9CM|PT|973.8|Poisoning by other specified agents primarily affecting the gastrointestinal system
C0161618|ICD9CM|AB|973.8|Poisoning-gi agents NEC
C0161619|ICD9CM|PT|973.9|Poisoning by unspecified agent primarily affecting the gastrointestinal system
C0161619|ICD9CM|AB|973.9|Poisoning-gi agent NOS
C0161621|ICD9CM|PT|974.0|Poisoning by mercurial diuretics
C0161621|ICD9CM|AB|974.0|Pois-mercurial diuretics
C0161622|ICD9CM|PT|974.1|Poisoning by purine derivative diuretics
C0161622|ICD9CM|AB|974.1|Pois-purine diuretics
C0161623|ICD9CM|PT|974.2|Poisoning by carbonic acid anhydrase inhibitors
C0161623|ICD9CM|AB|974.2|Pois-h2co3 anhydra inhib
C0161624|ICD9CM|PT|974.3|Poisoning by saluretics
C0161624|ICD9CM|AB|974.3|Poisoning-saluretics
C0161625|ICD9CM|PT|974.4|Poisoning by other diuretics
C0161625|ICD9CM|AB|974.4|Poisoning-diuretics NEC
C0161626|ICD9CM|PT|974.5|Poisoning by electrolytic, caloric, and water-balance agents
C0161626|ICD9CM|AB|974.5|Pois-electro/cal/wat agt
C0161628|ICD9CM|PT|974.7|Poisoning by uric acid metabolism drugs
C0161628|ICD9CM|AB|974.7|Pois-uric acid metabol
C0161629|ICD9CM|HT|975|Poisoning by agents primarily acting on the smooth and skeletal muscles and respiratory system
C0161630|ICD9CM|PT|975.0|Poisoning by oxytocic agents
C0161630|ICD9CM|AB|975.0|Poisoning-oxytocic agent
C0161631|ICD9CM|PT|975.1|Poisoning by smooth muscle relaxants
C0161631|ICD9CM|AB|975.1|Pois-smooth muscle relax
C0161632|ICD9CM|PT|975.2|Poisoning by skeletal muscle relaxants
C0161632|ICD9CM|AB|975.2|Pois-skelet muscle relax
C0161633|ICD9CM|PT|975.3|Poisoning by other and unspecified drugs acting on muscles
C0161633|ICD9CM|AB|975.3|Poison-muscle agent NEC
C0161634|ICD9CM|PT|975.4|Poisoning by antitussives
C0161634|ICD9CM|AB|975.4|Poisoning-antitussives
C0161635|ICD9CM|PT|975.5|Poisoning by expectorants
C0161635|ICD9CM|AB|975.5|Poisoning-expectorants
C0161636|ICD9CM|PT|975.6|Poisoning by anti-common cold drugs
C0161636|ICD9CM|AB|975.6|Pois-anti-cold drugs
C0161637|ICD9CM|PT|975.7|Poisoning by antiasthmatics
C0161637|ICD9CM|AB|975.7|Poisoning-antiasthmatics
C0161639|ICD9CM|HT|976|Poisoning by agents primarily affecting skin and mucous membrane, ophthalmological, otorhinolaryngological, and dental drugs
C0161640|ICD9CM|PT|976.0|Poisoning by local anti-infectives and anti-inflammatory drugs
C0161640|ICD9CM|AB|976.0|Pois-local anti-infect
C0161641|ICD9CM|PT|976.1|Poisoning by antipruritics
C0161641|ICD9CM|AB|976.1|Poisoning-antipruritics
C0161642|ICD9CM|PT|976.2|Poisoning by local astringents and local detergents
C0161642|ICD9CM|AB|976.2|Pois-loc astring/deterg
C0161643|ICD9CM|PT|976.3|Poisoning by emollients, demulcents, and protectants
C0161643|ICD9CM|AB|976.3|Pois-emol/demul/protect
C0161644|ICD9CM|PT|976.4|Poisoning by keratolytics, keratoplastics, other hair treatment drugs and preparations
C0161644|ICD9CM|AB|976.4|Poison-hair/scalp prep
C0161645|ICD9CM|PT|976.5|Poisoning by eye anti-infectives and other eye drugs
C0161645|ICD9CM|AB|976.5|Pois-eye anti-infec/drug
C0161646|ICD9CM|PT|976.6|Poisoning by anti-infectives and other drugs and preparations for ear, nose, and throat
C0161646|ICD9CM|AB|976.6|Poison-ent preparation
C0161647|ICD9CM|PT|976.7|Poisoning by dental drugs topically applied
C0161647|ICD9CM|AB|976.7|Pois-topical dental drug
C0161648|ICD9CM|PT|976.8|Poisoning by other agents primarily affecting skin and mucous membrane
C0161648|ICD9CM|AB|976.8|Pois-skin/membr agnt NEC
C0161649|ICD9CM|PT|976.9|Poisoning by unspecified agent primarily affecting skin and mucous membrane
C0161649|ICD9CM|AB|976.9|Pois-skin/membr agnt NOS
C0161651|ICD9CM|PT|977.0|Poisoning by dietetics
C0161651|ICD9CM|AB|977.0|Poisoning-dietetics
C0161652|ICD9CM|PT|977.1|Poisoning by lipotropic drugs
C0161652|ICD9CM|AB|977.1|Poison-lipotropic drugs
C0161654|ICD9CM|PT|977.3|Poisoning by alcohol deterrents
C0161654|ICD9CM|AB|977.3|Poison-alcohol deterrent
C0161655|ICD9CM|PT|977.4|Poisoning by pharmaceutical excipients
C0161655|ICD9CM|AB|977.4|Pois-pharmaceut excipien
C0161656|ICD9CM|PT|977.8|Poisoning by other specified drugs and medicinal substances
C0161656|ICD9CM|AB|977.8|Poison-medicinal agt NEC
C0161658|ICD9CM|HT|978|Poisoning by bacterial vaccines
C0161659|ICD9CM|PT|978.0|Poisoning by BCG vaccine
C0161659|ICD9CM|AB|978.0|Poisoning-bcg vaccine
C0161661|ICD9CM|PT|978.2|Poisoning by cholera vaccine
C0161661|ICD9CM|AB|978.2|Poisoning-cholera vaccin
C0161662|ICD9CM|PT|978.3|Poisoning by plague vaccine
C0161662|ICD9CM|AB|978.3|Poisoning-plague vaccine
C0161663|ICD9CM|PT|978.4|Poisoning by tetanus vaccine
C0161663|ICD9CM|AB|978.4|Poisoning-tetanus vaccin
C0161664|ICD9CM|PT|978.5|Poisoning by diphtheria vaccine
C0161664|ICD9CM|AB|978.5|Pois-diphtheria vaccine
C0161666|ICD9CM|PT|978.8|Poisoning by other and unspecified bacterial vaccines
C0161666|ICD9CM|AB|978.8|Pois-bact vaccin NEC/NOS
C0161669|ICD9CM|PT|979.0|Poisoning by smallpox vaccine
C0161669|ICD9CM|AB|979.0|Poison-smallpox vaccine
C0161670|ICD9CM|PT|979.1|Poisoning by rabies vaccine
C0161670|ICD9CM|AB|979.1|Poison-rabies vaccine
C0161671|ICD9CM|PT|979.2|Poisoning by typhus vaccine
C0161671|ICD9CM|AB|979.2|Poison-typhus vaccine
C0161672|ICD9CM|PT|979.3|Poisoning by yellow fever vaccine
C0161672|ICD9CM|AB|979.3|Pois-yellow fever vaccin
C0161673|ICD9CM|PT|979.4|Poisoning by measles vaccine
C0161673|ICD9CM|AB|979.4|Poisoning-measles vaccin
C0161674|ICD9CM|PT|979.5|Poisoning by poliomyelitis vaccine
C0161674|ICD9CM|AB|979.5|Pois-poliomyelit vaccine
C0161675|ICD9CM|PT|979.6|Poisoning by other and unspecified viral and rickettsial vaccines
C0161675|ICD9CM|AB|979.6|Pois-viral/rick vacc NEC
C0161676|ICD9CM|PT|979.7|Poisoning by mixed viral-rickettsial and bacterial vaccines, except combinations with a pertussis component
C0161676|ICD9CM|AB|979.7|Poisoning-mixed vaccine
C0161677|ICD9CM|PT|979.9|Poisoning by other and unspecified vaccines and biological substances
C0161677|ICD9CM|HT|979|Poisoning by other vaccines and biological substances
C0161677|ICD9CM|AB|979.9|Pois-vaccine/biolog NEC
C0161678|ICD9CM|HT|980|Toxic effect of alcohol
C0161678|ICD9CM|AB|980.9|Toxic effect alcohol NOS
C0161678|ICD9CM|PT|980.9|Toxic effect of unspecified alcohol
C0161679|ICD9CM|PT|980.0|Toxic effect of ethyl alcohol
C0161679|ICD9CM|AB|980.0|Toxic eff ethyl alcohol
C0161680|ICD9CM|PT|980.1|Toxic effect of methyl alcohol
C0161680|ICD9CM|AB|980.1|Toxic eff methyl alcohol
C0161681|ICD9CM|PT|980.2|Toxic effect of isopropyl alcohol
C0161681|ICD9CM|AB|980.2|Toxic eff isopropyl alc
C0161682|ICD9CM|PT|980.3|Toxic effect of fusel oil
C0161682|ICD9CM|AB|980.3|Toxic effect fusel oil
C0161683|ICD9CM|PT|980.8|Toxic effect of other specified alcohols
C0161683|ICD9CM|AB|980.8|Toxic effect alcohol NEC
C0161685|ICD9CM|PT|981|Toxic effect of petroleum products
C0161685|ICD9CM|AB|981|Toxic eff petroleum prod
C0161687|ICD9CM|PT|982.0|Toxic effect of benzene and homologues
C0161687|ICD9CM|AB|982.0|Toxic effect benzene
C0161689|ICD9CM|PT|982.2|Toxic effect of carbon disulfide
C0161689|ICD9CM|AB|982.2|Toxic eff carbon disulfi
C0161691|ICD9CM|PT|982.4|Toxic effect of nitroglycol
C0161691|ICD9CM|AB|982.4|Toxic effect nitroglycol
C0161692|ICD9CM|PT|982.8|Toxic effect of other nonpetroleum-based solvents
C0161692|ICD9CM|AB|982.8|Toxic eff nonpetrol solv
C0161693|ICD9CM|HT|983|Toxic effect of corrosive aromatics, acids, and caustic alkalis
C0161694|ICD9CM|PT|983.0|Toxic effect of corrosive aromatics
C0161694|ICD9CM|AB|983.0|Tox eff corrosive aromat
C0161695|ICD9CM|PT|983.1|Toxic effect of acids
C0161695|ICD9CM|AB|983.1|Toxic effect acids
C0161696|ICD9CM|PT|983.2|Toxic effect of caustic alkalis
C0161696|ICD9CM|AB|983.2|Toxic eff caustic alkali
C0161699|ICD9CM|PT|984.0|Toxic effect of inorganic lead compounds
C0161699|ICD9CM|AB|984.0|Tx eff inorg lead compnd
C0161700|ICD9CM|PT|984.1|Toxic effect of organic lead compounds
C0161700|ICD9CM|AB|984.1|Tox eff org lead compnd
C0161701|ICD9CM|PT|984.8|Toxic effect of other lead compounds
C0161701|ICD9CM|AB|984.8|Tox eff lead compnd NEC
C0161708|ICD9CM|PT|985.6|Toxic effect of chromium
C0161708|ICD9CM|AB|985.6|Toxic effect chromium
C0161709|ICD9CM|PT|985.9|Toxic effect of unspecified metal
C0161709|ICD9CM|AB|985.9|Toxic effect metal NOS
C0161713|ICD9CM|PT|987.2|Toxic effect of nitrogen oxides
C0161713|ICD9CM|AB|987.2|Toxic eff nitrogen oxide
C0161714|ICD9CM|PT|987.3|Toxic effect of sulfur dioxide
C0161714|ICD9CM|AB|987.3|Toxic eff sulfur dioxide
C0161715|ICD9CM|PT|987.4|Toxic effect of freon
C0161715|ICD9CM|AB|987.4|Toxic effect freon
C0161716|ICD9CM|PT|987.5|Toxic effect of lacrimogenic gas
C0161716|ICD9CM|AB|987.5|Tox eff lacrimogenic gas
C0161717|ICD9CM|PT|987.6|Toxic effect of chlorine gas
C0161717|ICD9CM|AB|987.6|Toxic eff chlorine gas
C0161718|ICD9CM|PT|987.7|Toxic effect of hydrocyanic acid gas
C0161718|ICD9CM|AB|987.7|Tox eff hydrocyan acd gs
C0161719|ICD9CM|PT|987.8|Toxic effect of other specified gases, fumes, or vapors
C0161719|ICD9CM|AB|987.8|Toxic eff gas/vapor NEC
C0161721|ICD9CM|HT|988|Toxic effect of noxious substances eaten as food
C0161721|ICD9CM|PT|988.9|Toxic effect of unspecified noxious substance eaten as food
C0161721|ICD9CM|AB|988.9|Tox eff noxious food NOS
C0161722|ICD9CM|PT|988.0|Toxic effect of fish and shellfish eaten as food
C0161722|ICD9CM|AB|988.0|Toxic eff fish/shellfish
C0161723|ICD9CM|PT|988.8|Toxic effect of other specified noxious substances eaten as food
C0161723|ICD9CM|AB|988.8|Tox eff noxious food NEC
C0161725|ICD9CM|HT|989|Toxic effect of other substances, chiefly nonmedicinal as to source
C0161725|ICD9CM|HT|989.8|Toxic effect of other substances, chiefly nonmedicinal as to source
C0161725|ICD9CM|PT|989.89|Toxic effect of other substance, chiefly nonmedicinal as to source, not elsewhere classified
C0161725|ICD9CM|AB|989.89|Tox eff nonmed subst NEC
C0161726|ICD9CM|PT|989.0|Toxic effect of hydrocyanic acid and cyanides
C0161726|ICD9CM|AB|989.0|Toxic effect cyanides
C0161727|ICD9CM|PT|989.1|Toxic effect of strychnine and salts
C0161727|ICD9CM|AB|989.1|Toxic effect strychnine
C0161732|ICD9CM|PT|989.7|Toxic effect of aflatoxin and other mycotoxin (food contaminants)
C0161732|ICD9CM|AB|989.7|Tox eff aflatox/mycotox
C0161734|ICD9CM|PT|991.9|Unspecified effect of reduced temperature
C0161734|ICD9CM|HT|991|Effects of reduced temperature
C0161734|ICD9CM|PT|E901.9|Accident due to excessive cold of unspecified origin
C0161734|ICD9CM|AB|E901.9|Excessive cold NOS
C0161734|ICD9CM|AB|991.9|Effect reduced temp NOS
C0161735|ICD9CM|AB|991.0|Frostbite of face
C0161735|ICD9CM|PT|991.0|Frostbite of face
C0161736|ICD9CM|AB|991.1|Frostbite of hand
C0161736|ICD9CM|PT|991.1|Frostbite of hand
C0161737|ICD9CM|AB|991.2|Frostbite of foot
C0161737|ICD9CM|PT|991.2|Frostbite of foot
C0161738|ICD9CM|PT|991.8|Other specified effects of reduced temperature
C0161738|ICD9CM|AB|991.8|Effect reduced temp NEC
C0161741|ICD9CM|AB|992.7|Heat edema
C0161741|ICD9CM|PT|992.7|Heat edema
C0161742|ICD9CM|PT|992.8|Other specified heat effects
C0161742|ICD9CM|AB|992.8|Heat effect NEC
C0161744|ICD9CM|AB|993.0|Barotrauma, otitic
C0161744|ICD9CM|PT|993.0|Barotrauma, otitic
C0161745|ICD9CM|AB|993.1|Barotrauma, sinus
C0161745|ICD9CM|PT|993.1|Barotrauma, sinus
C0161747|ICD9CM|PT|993.8|Other specified effects of air pressure
C0161747|ICD9CM|AB|993.8|Effect air pressure NEC
C0161748|ICD9CM|PT|993.9|Unspecified effect of air pressure
C0161748|ICD9CM|AB|993.9|Effect air pressure NOS
C0161749|ICD9CM|PT|994.4|Exhaustion due to exposure
C0161749|ICD9CM|AB|994.4|Exhaustion-exposure
C0161750|ICD9CM|PT|994.5|Exhaustion due to excessive exertion
C0161750|ICD9CM|AB|994.5|Exhaustion-excess exert
C0161751|ICD9CM|PT|994.7|Asphyxiation and strangulation
C0161751|ICD9CM|AB|994.7|Asphyxiation/strangulat
C0161752|ICD9CM|PT|994.8|Electrocution and nonfatal effects of electric current
C0161752|ICD9CM|AB|994.8|Effects electric current
C0161759|ICD9CM|PT|996.01|Mechanical complication due to cardiac pacemaker (electrode)
C0161759|ICD9CM|AB|996.01|Malfunc cardiac pacemake
C0161760|ICD9CM|PT|996.02|Mechanical complication due to heart valve prosthesis
C0161760|ICD9CM|AB|996.02|Malfunc prosth hrt valve
C0161761|ICD9CM|PT|996.03|Mechanical complication due to coronary bypass graft
C0161761|ICD9CM|AB|996.03|Malfunc coron bypass grf
C0161762|ICD9CM|PT|996.09|Other mechanical complication of cardiac device, implant, and graft
C0161762|ICD9CM|AB|996.09|Malfunc card dev/grf NEC
C0161763|ICD9CM|PT|996.1|Mechanical complication of other vascular device, implant, and graft
C0161763|ICD9CM|AB|996.1|Malfunc vasc device/graf
C0161767|ICD9CM|PT|996.31|Mechanical complication due to urethral (indwelling) catheter
C0161767|ICD9CM|AB|996.31|Malfunc urethral cath
C0161768|ICD9CM|PT|996.32|Mechanical complication due to intrauterine contraceptive device
C0161768|ICD9CM|AB|996.32|Malfunction iud
C0161769|ICD9CM|PT|996.39|Other mechanical complication of genitourinary device, implant, and graft
C0161769|ICD9CM|AB|996.39|Malfunc gu dev/graft NEC
C0161770|ICD9CM|HT|996.4|Mechanical complication of internal orthopedic device, implant, and graft
C0161771|ICD9CM|HT|996.5|Mechanical complication of other specified prosthetic device, implant, and graft
C0161777|ICD9CM|HT|996.6|Infection and inflammatory reaction due to internal prosthetic device, implant, and graft
C0161778|ICD9CM|PT|996.60|Infection and inflammatory reaction due to unspecified device, implant, and graft
C0161778|ICD9CM|AB|996.60|Reaction-unsp devic/grft
C0161779|ICD9CM|PT|996.61|Infection and inflammatory reaction due to cardiac device, implant, and graft
C0161779|ICD9CM|AB|996.61|React-cardiac dev/graft
C0161780|ICD9CM|PT|996.62|Infection and inflammatory reaction due to other vascular device, implant, and graft
C0161780|ICD9CM|AB|996.62|React-oth vasc dev/graft
C0161781|ICD9CM|PT|996.63|Infection and inflammatory reaction due to nervous system device, implant, and graft
C0161781|ICD9CM|AB|996.63|React-nerv sys dev/graft
C0161782|ICD9CM|PT|996.64|Infection and inflammatory reaction due to indwelling urinary catheter
C0161782|ICD9CM|AB|996.64|React-indwell urin cath
C0161783|ICD9CM|PT|996.65|Infection and inflammatory reaction due to other genitourinary device, implant, and graft
C0161783|ICD9CM|AB|996.65|React-oth genitourin dev
C0161784|ICD9CM|PT|996.66|Infection and inflammatory reaction due to internal joint prosthesis
C0161784|ICD9CM|AB|996.66|React-inter joint prost
C0161785|ICD9CM|PT|996.67|Infection and inflammatory reaction due to other internal orthopedic device, implant, and graft
C0161785|ICD9CM|AB|996.67|React-oth int ortho dev
C0161786|ICD9CM|PT|996.69|Infection and inflammatory reaction due to other internal prosthetic device, implant, and graft
C0161786|ICD9CM|AB|996.69|React-int pros devic NEC
C0161787|ICD9CM|HT|996.7|Other complications of internal (biological) (synthetic) prosthetic device, implant, and graft
C0161788|ICD9CM|PT|996.70|Other complications due to unspecified device, implant, and graft
C0161788|ICD9CM|AB|996.70|Comp-unsp device/graft
C0161789|ICD9CM|PT|996.71|Other complications due to heart valve prosthesis
C0161789|ICD9CM|AB|996.71|Comp-heart valve prosth
C0161790|ICD9CM|PT|996.72|Other complications due to other cardiac device, implant, and graft
C0161790|ICD9CM|AB|996.72|Comp-oth cardiac device
C0161791|ICD9CM|PT|996.73|Other complications due to renal dialysis device, implant, and graft
C0161791|ICD9CM|AB|996.73|Comp-ren dialys dev/grft
C0161792|ICD9CM|PT|996.74|Other complications due to other vascular device, implant, and graft
C0161792|ICD9CM|AB|996.74|Comp-oth vasc dev/graft
C0161794|ICD9CM|PT|996.76|Other complications due to genitourinary device, implant, and graft
C0161794|ICD9CM|AB|996.76|Comp-genitourin dev/grft
C0161795|ICD9CM|PT|996.77|Other complications due to internal joint prosthesis
C0161795|ICD9CM|AB|996.77|Comp-internal joint pros
C0161796|ICD9CM|PT|996.78|Other complications due to other internal orthopedic device, implant, and graft
C0161796|ICD9CM|AB|996.78|Comp-oth int ortho devic
C0161797|ICD9CM|PT|996.79|Other complications due to other internal prosthetic device, implant, and graft
C0161797|ICD9CM|AB|996.79|Comp-int prost devic NEC
C0161801|ICD9CM|PT|996.84|Complications of transplanted lung
C0161801|ICD9CM|AB|996.84|Compl lung transplant
C0161802|ICD9CM|PT|996.85|Complications of transplanted bone marrow
C0161802|ICD9CM|AB|996.85|Compl marrow transplant
C0161803|ICD9CM|PT|996.86|Complications of transplanted pancreas
C0161803|ICD9CM|AB|996.86|Compl pancreas transplnt
C0161804|ICD9CM|PT|996.89|Complications of other specified transplanted organ
C0161804|ICD9CM|AB|996.89|Comp oth organ transplnt
C0161805|ICD9CM|HT|996.9|Complications of reattached extremity or body part
C0161807|ICD9CM|PT|996.91|Complications of reattached forearm
C0161807|ICD9CM|AB|996.91|Compl reattached forearm
C0161808|ICD9CM|PT|996.92|Complications of reattached hand
C0161808|ICD9CM|AB|996.92|Compl reattached hand
C0161813|ICD9CM|PT|996.99|Complication of other specified reattached body part
C0161813|ICD9CM|AB|996.99|Compl reattach part NEC
C0161815|ICD9CM|PT|997.01|Central nervous system complication
C0161815|ICD9CM|AB|997.01|Surg complication - cns
C0161819|ICD9CM|HT|997.4|Digestive system complications
C0161821|ICD9CM|AB|997.60|Amputat stump compl NOS
C0161821|ICD9CM|PT|997.60|Unspecified complication of amputation stump
C0161824|ICD9CM|PT|997.62|Infection (chronic) of amputation stump
C0161824|ICD9CM|AB|997.62|Infection amputat stump
C0161829|ICD9CM|PT|998.2|Accidental puncture or laceration during a procedure, not elsewhere classified
C0161829|ICD9CM|AB|998.2|Accidental op laceration
C0161831|ICD9CM|PT|998.4|Foreign body accidentally left during a procedure
C0161831|ICD9CM|AB|998.4|FB left during procedure
C0161832|ICD9CM|PT|998.6|Persistent postoperative fistula
C0161832|ICD9CM|AB|998.6|Persist postop fistula
C0161833|ICD9CM|PT|998.7|Acute reaction to foreign substance accidentally left during a procedure
C0161833|ICD9CM|AB|998.7|Postop forgn subst react
C0161834|ICD9CM|PT|998.89|Other specified complications of procedures not elsewhere classified
C0161834|ICD9CM|AB|998.89|Oth spcf cmplc procd NEC
C0161841|ICD9CM|PT|E876.0|Mismatched blood in transfusion
C0161841|ICD9CM|AB|E876.0|Mismatch blood-transfusn
C0161848|ICD9CM|HT|01|Incision and excision of skull, brain, and cerebral meninges
C0161849|ICD9CM|PT|02.92|Repair of brain
C0161849|ICD9CM|AB|02.92|Brain repair
C0161850|ICD9CM|HT|02|Other operations on skull, brain, and cerebral meninges
C0161850|ICD9CM|HT|02.9|Other operations on skull, brain, and cerebral meninges
C0161850|ICD9CM|PT|02.99|Other operations on skull, brain, and cerebral meninges
C0161850|ICD9CM|AB|02.99|Skull & brain op NEC
C0161851|ICD9CM|HT|03|Operations on spinal cord and spinal canal structures
C0161852|ICD9CM|HT|04|Operations on cranial and peripheral nerves
C0161853|ICD9CM|HT|05|Operations on sympathetic nerves or ganglia
C0161855|ICD9CM|HT|07|Operations on other endocrine glands
C0161856|ICD9CM|HT|07.2|Partial adrenalectomy
C0161861|ICD9CM|HT|11.5|Repair of cornea
C0161862|ICD9CM|HT|12|Operations on iris, ciliary body, sclera, and anterior chamber
C0161864|ICD9CM|HT|14|Operations on retina, choroid, vitreous, and posterior chamber
C0161868|ICD9CM|HT|19|Reconstructive operations on middle ear
C0161869|ICD9CM|HT|19.2|Revision of stapedectomy
C0161870|ICD9CM|HT|20|Other operations on middle and inner ear
C0161870|ICD9CM|PT|20.99|Other operations on middle and inner ear
C0161870|ICD9CM|HT|20.9|Other operations on inner and middle ear
C0161870|ICD9CM|AB|20.99|Mid-inner ear ops NEC
C0161872|ICD9CM|HT|21.6|Turbinectomy
C0161874|ICD9CM|HT|23|Removal and restoration of teeth
C0161875|ICD9CM|HT|24|Other operations on teeth, gums, and alveoli
C0161878|ICD9CM|AB|27.24|Mouth biopsy NOS
C0161878|ICD9CM|PT|27.24|Biopsy of mouth, unspecified structure
C0161879|ICD9CM|HT|27.9|Other operations on mouth and face
C0161879|ICD9CM|HT|27|Other operations on mouth and face
C0161880|ICD9CM|AB|27.92|Mouth incision NOS
C0161880|ICD9CM|PT|27.92|Incision of mouth, unspecified structure
C0161884|ICD9CM|HT|31.2|Permanent tracheostomy
C0161885|ICD9CM|HT|31.9|Other operations on larynx and trachea
C0161885|ICD9CM|HT|31|Other operations on larynx and trachea
C0161887|ICD9CM|HT|33.9|Other operations on lung and bronchus
C0161887|ICD9CM|HT|33|Other operations on lung and bronchus
C0161888|ICD9CM|HT|34|Operations on chest wall, pleura, mediastinum, and diaphragm
C0161889|ICD9CM|AB|34.93|Repair of pleura
C0161889|ICD9CM|PT|34.93|Repair of pleura
C0161890|ICD9CM|HT|35|Operations on valves and septa of heart
C0161892|ICD9CM|HT|37|Other operations on heart and pericardium
C0161892|ICD9CM|HT|37.9|Other operations on heart and pericardium
C0161892|ICD9CM|PT|37.99|Other operations on heart and pericardium
C0161892|ICD9CM|AB|37.99|Other heart/pericard ops
C0161893|ICD9CM|HT|38|Incision, excision, and occlusion of vessels
C0161894|ICD9CM|HT|39|Other operations on vessels
C0161894|ICD9CM|HT|39.9|Other operations on vessels
C0161894|ICD9CM|PT|39.99|Other operations on vessels
C0161894|ICD9CM|AB|39.99|Vessel operation NEC
C0161896|ICD9CM|HT|41|Operations on bone marrow and spleen
C0161898|ICD9CM|HT|43|Incision and excision of stomach
C0161899|ICD9CM|HT|43.9|Total gastrectomy
C0161900|ICD9CM|HT|44|Other operations on stomach
C0161900|ICD9CM|HT|44.9|Other operations on stomach
C0161900|ICD9CM|PT|44.99|Other operations on stomach
C0161900|ICD9CM|AB|44.99|Gastric operation NEC
C0161901|ICD9CM|HT|45|Incision, excision, and anastomosis of intestine
C0161905|ICD9CM|HT|48|Operations on rectum, rectosigmoid and perirectal tissue
C0161906|ICD9CM|HT|48.7|Repair of rectum
C0161912|ICD9CM|HT|52.5|Partial pancreatectomy
C0161915|ICD9CM|HT|54.9|Other operations of abdominal region
C0161915|ICD9CM|PT|54.99|Other operations of abdominal region
C0161915|ICD9CM|HT|54|Other operations on abdominal region
C0161915|ICD9CM|AB|54.99|Abdomen region ops NEC
C0161918|ICD9CM|PT|56.73|Nephrocystanastomosis, not otherwise specified
C0161918|ICD9CM|AB|56.73|Nephrocystanastomosi NOS
C0161920|ICD9CM|HT|57|Operations on urinary bladder
C0161922|ICD9CM|HT|58.4|Repair of urethra
C0161924|ICD9CM|PT|59.00|Retroperitoneal dissection, not otherwise specified
C0161924|ICD9CM|AB|59.00|Retroperit dissect NOS
C0161925|ICD9CM|HT|60|Operations on prostate and seminal vesicles
C0161926|ICD9CM|HT|61|Operations on scrotum and tunica vaginalis
C0161928|ICD9CM|HT|63|Operations on spermatic cord, epididymis, and vas deferens
C0161930|ICD9CM|HT|65|Operations on ovary
C0161933|ICD9CM|HT|68|Other incision and excision of uterus
C0161934|ICD9CM|HT|69|Other operations on uterus and supporting structures
C0161935|ICD9CM|HT|70|Operations on vagina and cul-de-sac
C0161936|ICD9CM|HT|71|Operations on vulva and perineum
C0161937|ICD9CM|HT|72|Forceps, vacuum, and breech delivery
C0161939|ICD9CM|HT|73|Other procedures inducing or assisting delivery
C0161942|ICD9CM|HT|75|Other obstetric operations
C0161942|ICD9CM|HT|75.9|Other obstetric operations
C0161942|ICD9CM|PT|75.99|Other obstetric operations
C0161942|ICD9CM|AB|75.99|Obstetric operation NEC
C0161943|ICD9CM|HT|76|Operations on facial bones and joints
C0161944|ICD9CM|HT|77|Incision, excision, and division of other bones
C0161945|ICD9CM|HT|78|Other operations on bones, except facial bones
C0161946|ICD9CM|HT|79|Reduction of fracture and dislocation
C0161947|ICD9CM|HT|80|Incision and excision of joint structures
C0161948|ICD9CM|HT|81|Repair and plastic operations on joint structures
C0161950|ICD9CM|HT|83|Operations on muscle, tendon, fascia, and bursa, except hand
C0161954|ICD9CM|HT|86|Operations on skin and subcutaneous tissue
C0161955|ICD9CM|PT|86.60|Free skin graft, not otherwise specified
C0161955|ICD9CM|HT|86.6|Free skin graft
C0161955|ICD9CM|AB|86.60|Free skin graft NOS
C0161958|ICD9CM|HT|89|Interview, evaluation, consultation, and examination
C0161959|ICD9CM|HT|89.6|Circulatory monitoring
C0161960|ICD9CM|HT|90|Microscopic examination-I
C0161961|ICD9CM|HT|91|Microscopic examination-II
C0161962|ICD9CM|HT|93|Physical therapy, respiratory therapy, rehabilitation, and related procedures
C0161965|ICD9CM|HT|95|Ophthalmologic and otologic diagnosis and treatment
C0161966|ICD9CM|HT|96|Nonoperative intubation and irrigation
C0161967|ICD9CM|HT|97|Replacement and removal of therapeutic appliances
C0161968|ICD9CM|HT|98|Nonoperative removal of foreign body or calculus
C0161969|ICD9CM|HT|99|Other nonoperative procedures
C0161970|ICD9CM|PT|99.16|Injection of antidote
C0161970|ICD9CM|AB|99.16|Inject antidote
C0161972|ICD9CM|HT|670-677.99|COMPLICATIONS OF THE PUERPERIUM
C0161972|ICD9CM|HT|674.9|Unspecified complications of the puerperium
C0161972|ICD9CM|PT|674.90|Unspecified complications of puerperium, unspecified as to episode of care or not applicable
C0161972|ICD9CM|PT|674.94|Unspecified complications of puerperium, postpartum condition or complication
C0161972|ICD9CM|AB|674.94|Puerp compl NOS-postpart
C0161972|ICD9CM|AB|674.90|Puerp compl NOS-unspec
C0162019|ICD9CM|HT|376.4|Deformity of orbit
C0162019|ICD9CM|AB|376.40|Deformity of orbit NOS
C0162019|ICD9CM|PT|376.40|Deformity of orbit, unspecified
C0162164|ICD9CM|PT|746.02|Stenosis of pulmonary valve, congenital
C0162164|ICD9CM|AB|746.02|Cong pulmon valve stenos
C0162203|ICD9CM|PT|38.93|Venous catheterization, not elsewhere classified
C0162203|ICD9CM|AB|38.93|Venous cath NEC
C0162209|ICD9CM|PT|72.9|Unspecified instrumental delivery
C0162209|ICD9CM|AB|72.9|Instrument delivery NOS
C0162218|ICD9CM|PT|93.19|Exercise, not elsewhere classified
C0162218|ICD9CM|AB|93.19|Pt exercise NEC
C0162245|ICD9CM|PT|52.59|Other partial pancreatectomy
C0162245|ICD9CM|AB|52.59|Partial pancreatect NEC
C0162275|ICD9CM|AB|791.6|Acetonuria
C0162275|ICD9CM|PT|791.6|Acetonuria
C0162279|ICD9CM|HT|363.7|Choroidal detachment
C0162279|ICD9CM|AB|363.70|Choroidal detachment NOS
C0162279|ICD9CM|PT|363.70|Choroidal detachment, unspecified
C0162280|ICD9CM|AB|372.56|Conjunctival deposits
C0162280|ICD9CM|PT|372.56|Conjunctival deposits
C0162281|ICD9CM|AB|371.10|Corneal deposit NOS
C0162281|ICD9CM|PT|371.10|Corneal deposit, unspecified
C0162283|ICD9CM|PT|588.1|Nephrogenic diabetes insipidus
C0162283|ICD9CM|AB|588.1|Nephrogen diabetes insip
C0162285|ICD9CM|AB|374.82|Edema of eyelid
C0162285|ICD9CM|PT|374.82|Edema of eyelid
C0162286|ICD9CM|AB|947.2|Burn of esophagus
C0162286|ICD9CM|PT|947.2|Burn of esophagus
C0162287|ICD9CM|AB|787.7|Abnormal feces
C0162287|ICD9CM|PT|787.7|Abnormal feces
C0162291|ICD9CM|AB|362.84|Retinal ischemia
C0162291|ICD9CM|PT|362.84|Retinal ischemia
C0162292|ICD9CM|AB|378.55|External ophthalmoplegia
C0162292|ICD9CM|PT|378.55|External ophthalmoplegia
C0162296|ICD9CM|PT|719.49|Pain in joint, multiple sites
C0162296|ICD9CM|AB|719.49|Joint pain-mult jts
C0162297|ICD9CM|AB|799.1|Respiratory arrest
C0162297|ICD9CM|PT|799.1|Respiratory arrest
C0162299|ICD9CM|AB|246.2|Cyst of thyroid
C0162299|ICD9CM|PT|246.2|Cyst of thyroid
C0162301|ICD9CM|PT|594.2|Calculus in urethra
C0162301|ICD9CM|AB|594.2|Urethral calculus
C0162316|ICD9CM|HT|280|Iron deficiency anemias
C0162316|ICD9CM|PT|280.9|Iron deficiency anemia, unspecified
C0162316|ICD9CM|AB|280.9|Iron defic anemia NOS
C0162323|ICD9CM|PT|714.9|Unspecified inflammatory polyarthropathy
C0162323|ICD9CM|AB|714.9|Inflamm polyarthrop NOS
C0162352|ICD9CM|PT|99.12|Immunization for allergy
C0162352|ICD9CM|AB|99.12|Allergy immunization
C0162375|ICD9CM|PT|526.3|Central giant cell (reparative) granuloma
C0162375|ICD9CM|AB|526.3|Cent giant cell granulom
C0162423|ICD9CM|AB|705.1|Prickly heat
C0162423|ICD9CM|PT|705.1|Prickly heat
C0162482|ICD9CM|HT|665.2|Obstetrical inversion of uterus
C0162522|ICD9CM|PT|51.23|Laparoscopic cholecystectomy
C0162522|ICD9CM|AB|51.23|Laparoscopic cholecystec
C0162576|ICD9CM|AB|127.1|Anisakiasis
C0162576|ICD9CM|PT|127.1|Anisakiasis
C0162644|ICD9CM|PT|521.08|Dental caries of root surface
C0162644|ICD9CM|AB|521.08|Dental caries-root surf
C0162649|ICD9CM|PT|03.95|Spinal blood patch
C0162649|ICD9CM|AB|03.95|Spinal patch
C0162661|ICD9CM|HT|16.5|Exenteration of orbital contents
C0162662|ICD9CM|HT|16.3|Evisceration of eyeball
C0162674|ICD9CM|PT|378.72|Progressive external ophthalmoplegia
C0162674|ICD9CM|AB|378.72|Prog ext ophthalmoplegia
C0162678|ICD9CM|HT|237.7|Neurofibromatosis
C0162678|ICD9CM|AB|237.70|Neurofibromatosis NOS
C0162678|ICD9CM|PT|237.70|Neurofibromatosis, unspecified
C0162701|ICD9CM|AB|89.17|Polysomnogram
C0162701|ICD9CM|PT|89.17|Polysomnogram
C0162780|ICD9CM|AB|11.76|Epikeratophakia
C0162780|ICD9CM|PT|11.76|Epikeratophakia
C0162819|ICD9CM|PT|709.1|Vascular disorders of skin
C0162819|ICD9CM|AB|709.1|Vascular disord of skin
C0162849|ICD9CM|AB|697.1|Lichen nitidus
C0162849|ICD9CM|PT|697.1|Lichen nitidus
C0162870|ICD9CM|PT|442.2|Aneurysm of iliac artery
C0162870|ICD9CM|AB|442.2|Iliac artery aneurysm
C0175568|ICD9CM|HT|10.9|Other operations on conjunctiva
C0175568|ICD9CM|PT|10.99|Other operations on conjunctiva
C0175568|ICD9CM|AB|10.99|Conjunctival op NEC
C0175570|ICD9CM|HT|11.9|Other operations on cornea
C0175570|ICD9CM|PT|11.99|Other operations on cornea
C0175570|ICD9CM|AB|11.99|Corneal operation NEC
C0175572|ICD9CM|HT|13.5|Other extracapsular extraction of lens
C0175572|ICD9CM|PT|13.59|Other extracapsular extraction of lens
C0175572|ICD9CM|AB|13.59|Extracap lens extrac NEC
C0175574|ICD9CM|HT|24.9|Other dental operations
C0175574|ICD9CM|PT|24.99|Other dental operations
C0175574|ICD9CM|AB|24.99|Dental operation NEC
C0175578|ICD9CM|HT|29.5|Other repair of pharynx
C0175578|ICD9CM|PT|29.59|Other repair of pharynx
C0175578|ICD9CM|AB|29.59|Pharyngeal repair NEC
C0175580|ICD9CM|HT|29.9|Other operations on pharynx
C0175580|ICD9CM|PT|29.99|Other operations on pharynx
C0175580|ICD9CM|AB|29.99|Pharyngeal operation NEC
C0175582|ICD9CM|HT|30.2|Other partial laryngectomy
C0175582|ICD9CM|PT|30.29|Other partial laryngectomy
C0175582|ICD9CM|AB|30.29|Other part laryngectomy
C0175584|ICD9CM|HT|34.9|Other operations on thorax
C0175584|ICD9CM|PT|34.99|Other operations on thorax
C0175584|ICD9CM|AB|34.99|Thoracic operation NEC
C0175586|ICD9CM|HT|55.8|Other repair of kidney
C0175586|ICD9CM|PT|55.89|Other repair of kidney
C0175586|ICD9CM|AB|55.89|Renal repair NEC
C0175588|ICD9CM|HT|55.9|Other operations on kidney
C0175590|ICD9CM|HT|56.7|Other anastomosis or bypass of ureter
C0175590|ICD9CM|PT|56.79|Other anastomosis or bypass of ureter
C0175590|ICD9CM|AB|56.79|Ureteral anastomosis NEC
C0175594|ICD9CM|HT|57.9|Other operations on bladder
C0175594|ICD9CM|PT|57.99|Other operations on bladder
C0175594|ICD9CM|AB|57.99|Bladder operation NEC
C0175596|ICD9CM|HT|58.9|Other operations on urethra and periurethral tissue
C0175596|ICD9CM|PT|58.99|Other operations on urethra and periurethral tissue
C0175596|ICD9CM|AB|58.99|Ureth/periureth op NEC
C0175598|ICD9CM|HT|59|Other operations on urinary tract
C0175598|ICD9CM|HT|59.9|Other operations on urinary system
C0175598|ICD9CM|PT|59.99|Other operations on urinary system
C0175598|ICD9CM|AB|59.99|Urinary system op NEC
C0175600|ICD9CM|HT|60.9|Other operations on prostate
C0175600|ICD9CM|PT|60.99|Other operations on prostate
C0175600|ICD9CM|AB|60.99|Prostatic operation NEC
C0175608|ICD9CM|HT|65.9|Other operations on ovary
C0175608|ICD9CM|PT|65.99|Other operations on ovary
C0175608|ICD9CM|AB|65.99|Ovarian operation NEC
C0175610|ICD9CM|HT|66.9|Other operations on fallopian tubes
C0175610|ICD9CM|PT|66.99|Other operations on fallopian tubes
C0175610|ICD9CM|AB|66.99|Fallopian tube op NEC
C0175612|ICD9CM|HT|67.6|Other repair of cervix
C0175612|ICD9CM|PT|67.69|Other repair of cervix
C0175612|ICD9CM|AB|67.69|Cervical repair NEC
C0175614|ICD9CM|HT|70.7|Other repair of vagina
C0175614|ICD9CM|PT|70.79|Other repair of vagina
C0175614|ICD9CM|AB|70.79|Vaginal repair NEC
C0175616|ICD9CM|HT|75.6|Repair of other current obstetric laceration
C0175616|ICD9CM|PT|75.69|Repair of other current obstetric laceration
C0175616|ICD9CM|AB|75.69|Repair ob laceration NEC
C0175618|ICD9CM|HT|76.9|Other operations on facial bones and joints
C0175618|ICD9CM|PT|76.99|Other operations on facial bones and joints
C0175618|ICD9CM|AB|76.99|Facial bone/jnt op NEC
C0175620|ICD9CM|HT|81.9|Other operations on joint structures
C0175620|ICD9CM|PT|81.99|Other operations on joint structures
C0175620|ICD9CM|AB|81.99|Joint structure op NEC
C0175622|ICD9CM|HT|82.3|Other excision of soft tissue of hand
C0175622|ICD9CM|PT|82.39|Other excision of soft tissue of hand
C0175622|ICD9CM|AB|82.39|Hand soft tissue exc NEC
C0175624|ICD9CM|HT|17|Other miscellaneous procedures
C0175624|ICD9CM|PT|99.99|Other miscellaneous procedures
C0175624|ICD9CM|HT|99.9|Other miscellaneous procedures
C0175624|ICD9CM|AB|99.99|Miscellaneous proc NEC
C0175708|ICD9CM|HT|393-398.99|CHRONIC RHEUMATIC HEART DISEASE
C0175757|ICD9CM|AB|56.1|Ureteral meatotomy
C0175757|ICD9CM|PT|56.1|Ureteral meatotomy
C0175759|ICD9CM|AB|34.02|Exploratory thoracotomy
C0175759|ICD9CM|PT|34.02|Exploratory thoracotomy
C0175760|ICD9CM|PT|77.25|Wedge osteotomy, femur
C0175760|ICD9CM|AB|77.25|Femoral wedge osteotomy
C0175761|ICD9CM|AB|35.34|Infundibulectomy
C0175761|ICD9CM|PT|35.34|Infundibulectomy
C0175763|ICD9CM|AB|01.52|Hemispherectomy
C0175763|ICD9CM|PT|01.52|Hemispherectomy
C0175999|ICD9CM|PT|515|Postinflammatory pulmonary fibrosis
C0175999|ICD9CM|AB|515|Postinflam pulm fibrosis
C0176004|ICD9CM|HT|E829|Other road vehicle accidents
C0176004|ICD9CM|HT|E826-E829.9|OTHER ROAD VEHICLE ACCIDENTS
C0176005|ICD9CM|HT|E929|Late effects of accidental injury
C0176005|ICD9CM|HT|E929-E929.9|LATE EFFECTS OF ACCIDENTAL INJURY
C0176006|ICD9CM|PT|01.02|Ventriculopuncture through previously implanted catheter
C0176006|ICD9CM|AB|01.02|Ventricl shunt tube punc
C0176007|ICD9CM|PT|01.09|Other cranial puncture
C0176007|ICD9CM|AB|01.09|Cranial puncture NEC
C0176008|ICD9CM|HT|01.1|Diagnostic procedures on skull, brain, and cerebral meninges
C0176010|ICD9CM|PT|01.12|Open biopsy of cerebral meninges
C0176010|ICD9CM|AB|01.12|Open cereb meninges bx
C0176013|ICD9CM|PT|01.18|Other diagnostic procedures on brain and cerebral meninges
C0176013|ICD9CM|AB|01.18|Other brain dx procedure
C0176014|ICD9CM|PT|01.19|Other diagnostic procedures on skull
C0176014|ICD9CM|AB|01.19|Other skull dx procedure
C0176015|ICD9CM|HT|01.2|Craniotomy and craniectomy
C0176016|ICD9CM|AB|01.25|Other craniectomy
C0176016|ICD9CM|PT|01.25|Other craniectomy
C0176017|ICD9CM|HT|01.3|Incision of brain and cerebral meninges
C0176018|ICD9CM|PT|01.39|Other incision of brain
C0176018|ICD9CM|AB|01.39|Other brain incision
C0176019|ICD9CM|HT|01.4|Operations on thalamus and globus pallidus
C0176020|ICD9CM|PT|01.41|Operations on thalamus
C0176020|ICD9CM|AB|01.41|Thalamus operations
C0176022|ICD9CM|HT|01.5|Other excision or destruction of brain and meninges
C0176023|ICD9CM|PT|01.51|Excision of lesion or tissue of cerebral meninges
C0176023|ICD9CM|AB|01.51|Ex cereb meningeal les
C0176024|ICD9CM|PT|01.59|Other excision or destruction of lesion or tissue of brain
C0176024|ICD9CM|AB|01.59|Other brain excision
C0176025|ICD9CM|PT|02.03|Formation of cranial bone flap
C0176025|ICD9CM|AB|02.03|Skull flap formation
C0176026|ICD9CM|PT|02.06|Other cranial osteoplasty
C0176026|ICD9CM|AB|02.06|Cranial osteoplasty NEC
C0176027|ICD9CM|PT|02.12|Other repair of cerebral meninges
C0176027|ICD9CM|AB|02.12|Brain meninge repair NEC
C0176028|ICD9CM|PT|02.13|Ligation of meningeal vessel
C0176028|ICD9CM|AB|02.13|Meninge vessel ligation
C0176030|ICD9CM|PT|02.31|Ventricular shunt to structure in head and neck
C0176030|ICD9CM|AB|02.31|Ventricl shunt-head/neck
C0176031|ICD9CM|PT|02.33|Ventricular shunt to thoracic cavity
C0176031|ICD9CM|AB|02.33|Ventricl shunt-thorax
C0176032|ICD9CM|PT|02.34|Ventricular shunt to abdominal cavity and organs
C0176032|ICD9CM|AB|02.34|Ventricl shunt-abdomen
C0176034|ICD9CM|HT|02.4|Revision, removal, and irrigation of ventricular shunt
C0176036|ICD9CM|PT|02.91|Lysis of cortical adhesions
C0176036|ICD9CM|AB|02.91|Lysis cortical adhesion
C0176038|ICD9CM|PT|02.94|Insertion or replacement of skull tongs or halo traction device
C0176038|ICD9CM|AB|02.94|Insert/replac skull tong
C0176039|ICD9CM|PT|02.95|Removal of skull tongs or halo traction device
C0176039|ICD9CM|AB|02.95|Remove skull tongs
C0176040|ICD9CM|HT|03.0|Exploration and decompression of spinal canal structures
C0176044|ICD9CM|HT|03.3|Diagnostic procedures on spinal cord and spinal canal structures
C0176045|ICD9CM|PT|03.32|Biopsy of spinal cord or spinal meninges
C0176045|ICD9CM|AB|03.32|Spinal cord/meninges bx
C0176046|ICD9CM|PT|03.39|Other diagnostic procedures on spinal cord and spinal canal structures
C0176046|ICD9CM|AB|03.39|Other spinal dx proc
C0176047|ICD9CM|PT|03.4|Excision or destruction of lesion of spinal cord or spinal meninges
C0176047|ICD9CM|AB|03.4|Excis spinal cord lesion
C0176048|ICD9CM|HT|03.5|Plastic operations on spinal cord structures
C0176049|ICD9CM|PT|03.59|Other repair and plastic operations on spinal cord structures
C0176049|ICD9CM|AB|03.59|Spinal struct repair NEC
C0176050|ICD9CM|HT|03.7|Shunt of spinal theca
C0176051|ICD9CM|PT|03.79|Other shunt of spinal theca
C0176051|ICD9CM|AB|03.79|Oth spinal thecal shunt
C0176053|ICD9CM|PT|03.90|Insertion of catheter into spinal canal for infusion of therapeutic or palliative substances
C0176053|ICD9CM|AB|03.90|Insert spinal canal cath
C0176054|ICD9CM|PT|03.91|Injection of anesthetic into spinal canal for analgesia
C0176054|ICD9CM|AB|03.91|Anesth inject-spin canal
C0176056|ICD9CM|HT|04.0|Incision, division, and excision of cranial and peripheral nerves
C0176057|ICD9CM|PT|04.04|Other incision of cranial and peripheral nerves
C0176057|ICD9CM|AB|04.04|Periph nerve incis NEC
C0176058|ICD9CM|PT|04.06|Other cranial or peripheral ganglionectomy
C0176058|ICD9CM|AB|04.06|Periph ganglionect NEC
C0176059|ICD9CM|PT|04.07|Other excision or avulsion of cranial and peripheral nerves
C0176059|ICD9CM|AB|04.07|Periph nerv excision NEC
C0176060|ICD9CM|HT|04.1|Diagnostic procedures on peripheral nervous system
C0176061|ICD9CM|PT|04.11|Closed [percutaneous] [needle] biopsy of cranial or peripheral nerve or ganglion
C0176061|ICD9CM|AB|04.11|Clos periph nerve biopsy
C0176062|ICD9CM|PT|04.12|Open biopsy of cranial or peripheral nerve or ganglion
C0176062|ICD9CM|AB|04.12|Open periph nerve biopsy
C0176063|ICD9CM|PT|04.19|Other diagnostic procedures on cranial and peripheral nerves and ganglia
C0176063|ICD9CM|AB|04.19|Periph nerve dx proc NEC
C0176064|ICD9CM|PT|04.2|Destruction of cranial and peripheral nerves
C0176064|ICD9CM|AB|04.2|Periph nerve destruction
C0176065|ICD9CM|PT|04.3|Suture of cranial and peripheral nerves
C0176065|ICD9CM|AB|04.3|Peripheral nerve suture
C0176066|ICD9CM|HT|04.4|Lysis of adhesions and decompression of cranial and peripheral nerves
C0176067|ICD9CM|PT|04.42|Other cranial nerve decompression
C0176067|ICD9CM|AB|04.42|Cran nerv root decom NEC
C0176069|ICD9CM|PT|04.49|Other peripheral nerve or ganglion decompression or lysis of adhesions
C0176069|ICD9CM|AB|04.49|Per nerve adhesiolys NEC
C0176070|ICD9CM|PT|04.5|Cranial or peripheral nerve graft
C0176070|ICD9CM|AB|04.5|Peripheral nerve graft
C0176071|ICD9CM|HT|04.7|Other cranial or peripheral neuroplasty
C0176075|ICD9CM|PT|04.74|Other anastomosis of cranial or peripheral nerve
C0176075|ICD9CM|AB|04.74|Periph nerv anastom NEC
C0176076|ICD9CM|PT|04.75|Revision of previous repair of cranial and peripheral nerves
C0176076|ICD9CM|AB|04.75|Postop revis per nerv op
C0176077|ICD9CM|PT|04.76|Repair of old traumatic injury of cranial and peripheral nerves
C0176077|ICD9CM|AB|04.76|Late repair per nerv inj
C0176078|ICD9CM|AB|04.79|Other neuroplasty
C0176078|ICD9CM|PT|04.79|Other neuroplasty
C0176079|ICD9CM|HT|04.8|Injection into peripheral nerve
C0176081|ICD9CM|PT|04.89|Injection of other agent, except neurolytic
C0176081|ICD9CM|AB|04.89|Periph nerve inject NEC
C0176082|ICD9CM|HT|04.9|Other operations on cranial and peripheral nerves
C0176082|ICD9CM|PT|04.99|Other operations on cranial and peripheral nerves
C0176082|ICD9CM|AB|04.99|Peripheral nerve ops NEC
C0176085|ICD9CM|PT|05.0|Division of sympathetic nerve or ganglion
C0176085|ICD9CM|AB|05.0|Sympath nerve division
C0176086|ICD9CM|HT|05.1|Diagnostic procedures on sympathetic nerves or ganglia
C0176087|ICD9CM|PT|05.11|Biopsy of sympathetic nerve or ganglion
C0176087|ICD9CM|AB|05.11|Sympathetic nerve biopsy
C0176088|ICD9CM|PT|05.19|Other diagnostic procedures on sympathetic nerves or ganglia
C0176088|ICD9CM|AB|05.19|Sympath nrv dx proc NEC
C0176089|ICD9CM|HT|05.3|Injection into sympathetic nerve or ganglion
C0176091|ICD9CM|PT|05.39|Other injection into sympathetic nerve or ganglion
C0176091|ICD9CM|AB|05.39|Sympath nerve inject NEC
C0176092|ICD9CM|HT|05.8|Other operations on sympathetic nerves or ganglia
C0176092|ICD9CM|PT|05.89|Other operations on sympathetic nerves or ganglia
C0176092|ICD9CM|AB|05.89|Sympathetic nerve op NEC
C0176093|ICD9CM|PT|05.81|Repair of sympathetic nerve or ganglion
C0176093|ICD9CM|AB|05.81|Sympathetic nerve repair
C0176094|ICD9CM|PT|05.9|Other operations on nervous system
C0176094|ICD9CM|AB|05.9|Other nervous system ops
C0176095|ICD9CM|HT|06.0|Incision of thyroid field
C0176098|ICD9CM|PT|06.09|Other incision of thyroid field
C0176098|ICD9CM|AB|06.09|Incis thyroid field NEC
C0176099|ICD9CM|HT|06.1|Diagnostic procedures on thyroid and parathyroid glands
C0176100|ICD9CM|PT|06.11|Closed [percutaneous] [needle] biopsy of thyroid gland
C0176100|ICD9CM|AB|06.11|Closed thyroid gland bx
C0176101|ICD9CM|PT|06.12|Open biopsy of thyroid gland
C0176101|ICD9CM|AB|06.12|Open thyroid gland bx
C0176102|ICD9CM|PT|06.19|Other diagnostic procedures on thyroid and parathyroid glands
C0176102|ICD9CM|AB|06.19|Thyr/parathy dx proc NEC
C0176103|ICD9CM|PT|06.7|Excision of thyroglossal duct or tract
C0176103|ICD9CM|AB|06.7|Thyrogloss duct excision
C0176104|ICD9CM|HT|06.9|Other operations on thyroid (region) and parathyroid
C0176106|ICD9CM|PT|06.92|Ligation of thyroid vessels
C0176106|ICD9CM|AB|06.92|Thyroid vessel ligation
C0176108|ICD9CM|PT|06.95|Parathyroid tissue reimplantation
C0176108|ICD9CM|AB|06.95|Parathyroid reimplant
C0176109|ICD9CM|PT|06.98|Other operations on thyroid glands
C0176109|ICD9CM|AB|06.98|Other thyroid operations
C0176110|ICD9CM|PT|06.99|Other operations on parathyroid glands
C0176110|ICD9CM|AB|06.99|Other parathyroid ops
C0176112|ICD9CM|PT|07.01|Unilateral exploration of adrenal field
C0176112|ICD9CM|AB|07.01|Unilat adrenal explorat
C0176114|ICD9CM|HT|07.1|Diagnostic procedures on adrenal glands, pituitary gland, pineal gland, and thymus
C0176117|ICD9CM|PT|07.13|Biopsy of pituitary gland, transfrontal approach
C0176117|ICD9CM|AB|07.13|Transfront pituitary bx
C0176118|ICD9CM|PT|07.14|Biopsy of pituitary gland, transsphenoidal approach
C0176118|ICD9CM|AB|07.14|Transphen pituitary bx
C0176120|ICD9CM|PT|07.17|Biopsy of pineal gland
C0176120|ICD9CM|AB|07.17|Pineal biopsy
C0176121|ICD9CM|PT|07.19|Other diagnostic procedures on adrenal glands, pituitary gland, pineal gland, and thymus
C0176121|ICD9CM|AB|07.19|Endocrine dx proc NEC
C0176122|ICD9CM|PT|07.29|Other partial adrenalectomy
C0176122|ICD9CM|AB|07.29|Part adrenalectomy NEC
C0176123|ICD9CM|HT|07.4|Other operations on adrenal glands, nerves, and vessels
C0176123|ICD9CM|PT|07.49|Other operations on adrenal glands, nerves, and vessels
C0176123|ICD9CM|AB|07.49|Adrenal operation NEC
C0176124|ICD9CM|PT|07.43|Ligation of adrenal vessels
C0176124|ICD9CM|AB|07.43|Adrenal vessel ligation
C0176127|ICD9CM|PT|07.51|Exploration of pineal field
C0176127|ICD9CM|AB|07.51|Pineal field exploration
C0176128|ICD9CM|PT|07.59|Other operations on pineal gland
C0176128|ICD9CM|AB|07.59|Pineal operation NEC
C0176134|ICD9CM|PT|07.68|Total excision of pituitary gland, other specified approach
C0176134|ICD9CM|AB|07.68|Total exc pituitary NEC
C0176135|ICD9CM|HT|07.7|Other operations on hypophysis
C0176135|ICD9CM|PT|07.79|Other operations on hypophysis
C0176135|ICD9CM|AB|07.79|Pituitary operation NEC
C0176136|ICD9CM|PT|07.71|Exploration of pituitary fossa
C0176136|ICD9CM|AB|07.71|Pituitary fossa explorat
C0176137|ICD9CM|HT|07.9|Other operations on thymus
C0176138|ICD9CM|PT|07.91|Exploration of thymus field
C0176138|ICD9CM|AB|07.91|Thymus field exploration
C0176140|ICD9CM|PT|08.09|Other incision of eyelid
C0176140|ICD9CM|AB|08.09|Other eyelid incision
C0176142|ICD9CM|PT|08.19|Other diagnostic procedures on eyelid
C0176142|ICD9CM|AB|08.19|Eyelid dx procedure NEC
C0176144|ICD9CM|PT|08.21|Excision of chalazion
C0176144|ICD9CM|AB|08.21|Chalazion excision
C0176145|ICD9CM|PT|08.22|Excision of other minor lesion of eyelid
C0176145|ICD9CM|AB|08.22|Excise minor les lid NEC
C0176146|ICD9CM|HT|08.3|Repair of blepharoptosis and lid retraction
C0176149|ICD9CM|HT|08.4|Repair of entropion or ectropion
C0176150|ICD9CM|PT|08.41|Repair of entropion or ectropion by thermocauterization
C0176150|ICD9CM|AB|08.41|Thermocaut/entropion rep
C0176153|ICD9CM|PT|08.44|Repair of entropion or ectropion with lid reconstruction
C0176153|ICD9CM|AB|08.44|Lid recons entropion rep
C0176154|ICD9CM|PT|08.49|Other repair of entropion or ectropion
C0176154|ICD9CM|AB|08.49|Entropion/ectrop rep NEC
C0176155|ICD9CM|HT|08.5|Other adjustment of lid position
C0176155|ICD9CM|PT|08.59|Other adjustment of lid position
C0176155|ICD9CM|AB|08.59|Adjust lid position NEC
C0176156|ICD9CM|HT|08.6|Reconstruction of eyelid with flaps or grafts
C0176157|ICD9CM|PT|08.61|Reconstruction of eyelid with skin flap or graft
C0176157|ICD9CM|AB|08.61|Lid reconst w skin graft
C0176158|ICD9CM|PT|08.62|Reconstruction of eyelid with mucous membrane flap or graft
C0176158|ICD9CM|AB|08.62|Lid reconst w muc graft
C0176159|ICD9CM|PT|08.69|Other reconstruction of eyelid with flaps or grafts
C0176159|ICD9CM|AB|08.69|Lid reconstr w graft NEC
C0176160|ICD9CM|HT|08.7|Other reconstruction of eyelid
C0176162|ICD9CM|PT|08.72|Other reconstruction of eyelid, partial-thickness
C0176162|ICD9CM|AB|08.72|Lid recons-part thic NEC
C0176163|ICD9CM|PT|08.74|Other reconstruction of eyelid, full-thickness
C0176163|ICD9CM|AB|08.74|Lid reconst-ful thic NEC
C0176165|ICD9CM|PT|08.81|Linear repair of laceration of eyelid or eyebrow
C0176165|ICD9CM|AB|08.81|Linear rep lid lacer
C0176167|ICD9CM|PT|08.83|Other repair of laceration of eyelid, partial-thickness
C0176167|ICD9CM|AB|08.83|Lid lacer rx-prt th NEC
C0176169|ICD9CM|PT|08.85|Other repair of laceration of eyelid, full-thickness
C0176169|ICD9CM|AB|08.85|Lid lac rx-ful thic NEC
C0176172|ICD9CM|HT|08.8|Other repair of eyelid
C0176172|ICD9CM|PT|08.89|Other eyelid repair
C0176172|ICD9CM|AB|08.89|Eyelid repair NEC
C0176173|ICD9CM|HT|08.9|Other operations on eyelids
C0176173|ICD9CM|PT|08.99|Other operations on eyelids
C0176173|ICD9CM|AB|08.99|Eyelid operation NEC
C0176174|ICD9CM|PT|08.93|Other epilation of eyelid
C0176174|ICD9CM|AB|08.93|Eyelid epilation NEC
C0176176|ICD9CM|PT|09.19|Other diagnostic procedures on lacrimal system
C0176176|ICD9CM|AB|09.19|Lacrimal sys dx proc NEC
C0176177|ICD9CM|HT|09.2|Excision of lesion or tissue of lacrimal gland
C0176178|ICD9CM|PT|09.21|Excision of lesion of lacrimal gland
C0176178|ICD9CM|AB|09.21|Excis les lacrimal gland
C0176179|ICD9CM|PT|09.22|Other partial dacryoadenectomy
C0176179|ICD9CM|AB|09.22|Part dacryoadenect NEC
C0176180|ICD9CM|PT|09.3|Other operations on lacrimal gland
C0176180|ICD9CM|AB|09.3|Other lacrimal gland ops
C0176182|ICD9CM|PT|09.49|Other manipulation of lacrimal passage
C0176182|ICD9CM|AB|09.49|Lac passage manip NEC
C0176183|ICD9CM|HT|09.5|Incision of lacrimal sac and passages
C0176184|ICD9CM|PT|09.59|Other incision of lacrimal passages
C0176184|ICD9CM|AB|09.59|Lacrim passage incis NEC
C0176185|ICD9CM|PT|09.6|Excision of lacrimal sac and passage
C0176185|ICD9CM|AB|09.6|Lacrim sac/passage excis
C0176186|ICD9CM|HT|09.7|Repair of canaliculus and punctum
C0176187|ICD9CM|PT|09.71|Correction of everted punctum
C0176187|ICD9CM|AB|09.71|Correct everted punctum
C0176188|ICD9CM|PT|09.72|Other repair of punctum
C0176188|ICD9CM|AB|09.72|Punctum repair NEC
C0176189|ICD9CM|PT|09.73|Repair of canaliculus
C0176189|ICD9CM|AB|09.73|Canaliculus repair
C0176190|ICD9CM|HT|09.8|Fistulization of lacrimal tract to nasal cavity
C0176191|ICD9CM|PT|09.83|Conjunctivorhinostomy with insertion of tube or stent
C0176191|ICD9CM|AB|09.83|Conjunctivorhinos w tube
C0176192|ICD9CM|HT|09.9|Other operations on lacrimal system
C0176192|ICD9CM|PT|09.99|Other operations on lacrimal system
C0176192|ICD9CM|AB|09.99|Lacrimal system op NEC
C0176193|ICD9CM|PT|10.1|Other incision of conjunctiva
C0176193|ICD9CM|AB|10.1|Conjunctiva incision NEC
C0176195|ICD9CM|PT|10.29|Other diagnostic procedures on conjunctiva
C0176195|ICD9CM|AB|10.29|Conjunctiva dx proc NEC
C0176196|ICD9CM|HT|10.3|Excision or destruction of lesion or tissue of conjunctiva
C0176197|ICD9CM|PT|10.31|Excision of lesion or tissue of conjunctiva
C0176197|ICD9CM|AB|10.31|Excise conjunctiv lesion
C0176198|ICD9CM|PT|10.33|Other destructive procedures on conjunctiva
C0176198|ICD9CM|AB|10.33|Oth conjunc destruc proc
C0176199|ICD9CM|PT|10.42|Reconstruction of conjunctival cul-de-sac with free graft
C0176199|ICD9CM|AB|10.42|Graft conjunc cul-de-sac
C0176200|ICD9CM|PT|10.43|Other reconstruction of conjunctival cul-de-sac
C0176200|ICD9CM|AB|10.43|Conjun cul-de-sac rx NEC
C0176201|ICD9CM|PT|10.44|Other free graft to conjunctiva
C0176201|ICD9CM|AB|10.44|Conjunc free graft NEC
C0176202|ICD9CM|PT|10.49|Other conjunctivoplasty
C0176202|ICD9CM|AB|10.49|Conjunctivoplasty NEC
C0176203|ICD9CM|PT|10.5|Lysis of adhesions of conjunctiva and eyelid
C0176203|ICD9CM|AB|10.5|Conjunc/lid adhesiolysis
C0176206|ICD9CM|PT|11.21|Scraping of cornea for smear or culture
C0176206|ICD9CM|AB|11.21|Corneal scrape for smear
C0176207|ICD9CM|PT|11.29|Other diagnostic procedures on cornea
C0176207|ICD9CM|AB|11.29|Corneal dx proc NEC
C0176209|ICD9CM|PT|11.39|Other excision of pterygium
C0176209|ICD9CM|AB|11.39|Pterygium excision NEC
C0176210|ICD9CM|HT|11.4|Excision or destruction of tissue or other lesion of cornea
C0176211|ICD9CM|PT|11.42|Thermocauterization of corneal lesion
C0176211|ICD9CM|AB|11.42|Thermocaut cornea lesion
C0176212|ICD9CM|PT|11.49|Other removal or destruction of corneal lesion
C0176212|ICD9CM|AB|11.49|Destruct cornea les NEC
C0176213|ICD9CM|PT|11.53|Repair of corneal laceration or wound with conjunctival flap
C0176213|ICD9CM|AB|11.53|Rx cornea lac w conj flp
C0176214|ICD9CM|PT|11.59|Other repair of cornea
C0176214|ICD9CM|AB|11.59|Corneal repair NEC
C0176215|ICD9CM|PT|11.62|Other lamellar keratoplasty
C0176215|ICD9CM|AB|11.62|Lamellar keratoplast NEC
C0176217|ICD9CM|AB|11.73|Keratoprosthesis
C0176217|ICD9CM|PT|11.73|Keratoprosthesis
C0176218|ICD9CM|HT|11.7|Other reconstructive and refractive surgery on cornea
C0176218|ICD9CM|PT|11.79|Other reconstructive and refractive surgery on cornea
C0176218|ICD9CM|AB|11.79|Cornea reconstruct NEC
C0176219|ICD9CM|PT|12.02|Removal of intraocular foreign body from anterior segment of eye without use of magnet
C0176219|ICD9CM|AB|12.02|Nonmag remov ant seg FB
C0176220|ICD9CM|HT|12.1|Iridotomy and simple iridectomy
C0176221|MTH|PN|NOCODE|Iridotomy NEC in ICD9CM_2014
C0176221|ICD9CM|PT|12.12|Other iridotomy
C0176221|ICD9CM|AB|12.12|Iridotomy NEC
C0176222|MTH|PN|NOCODE|Iridectomy NEC in ICD9CM_2014
C0176222|ICD9CM|PT|12.14|Other iridectomy
C0176222|ICD9CM|AB|12.14|Iridectomy NEC
C0176223|ICD9CM|HT|12.2|Diagnostic procedures on iris, ciliary body, sclera, and anterior chamber
C0176224|ICD9CM|HT|12.3|Iridoplasty and coreoplasty
C0176225|ICD9CM|PT|12.32|Lysis of other anterior synechiae
C0176225|ICD9CM|AB|12.32|Ant synechia lysis NEC
C0176226|MTH|PN|NOCODE|Iridoplasty NEC in ICD9CM_2014
C0176226|ICD9CM|PT|12.39|Other iridoplasty
C0176226|ICD9CM|AB|12.39|Iridoplasty NEC
C0176227|ICD9CM|HT|12.4|Excision or destruction of lesion of iris and ciliary body
C0176229|ICD9CM|PT|12.65|Other scleral fistulization with iridectomy
C0176229|ICD9CM|AB|12.65|Scler fistuliz w iridect
C0176230|ICD9CM|PT|12.69|Other scleral fistulizing procedure
C0176230|ICD9CM|AB|12.69|Scler fistulizing op NEC
C0176231|ICD9CM|HT|12.7|Other procedures for relief of elevated intraocular pressure
C0176232|ICD9CM|PT|12.79|Other glaucoma procedures
C0176232|ICD9CM|AB|12.79|Glaucoma procedure NEC
C0176235|ICD9CM|PT|12.84|Excision or destruction of lesion of sclera
C0176235|ICD9CM|AB|12.84|Destruct scleral lesion
C0176236|ICD9CM|PT|12.86|Other repair of scleral staphyloma
C0176236|ICD9CM|AB|12.86|Rep scler staphyloma NEC
C0176237|ICD9CM|PT|12.88|Other scleral reinforcement
C0176237|ICD9CM|AB|12.88|Sclera reinforcement NEC
C0176238|ICD9CM|PT|12.89|Other operations on sclera
C0176238|ICD9CM|AB|12.89|Scleral operation NEC
C0176239|ICD9CM|HT|12.9|Other operations on iris, ciliary body, and anterior chamber
C0176242|ICD9CM|PT|12.93|Removal or destruction of epithelial downgrowth from anterior chamber
C0176242|ICD9CM|AB|12.93|Remov epithel downgrowth
C0176243|ICD9CM|PT|12.97|Other operations on iris
C0176243|ICD9CM|AB|12.97|Iris operation NEC
C0176244|ICD9CM|PT|12.98|Other operations on ciliary body
C0176244|ICD9CM|AB|12.98|Ciliary body op NEC
C0176245|ICD9CM|PT|12.99|Other operations on anterior chamber
C0176245|ICD9CM|AB|12.99|Anterior chamber op NEC
C0176247|ICD9CM|HT|13.4|Extracapsular extraction of lens by fragmentation and aspiration technique
C0176248|ICD9CM|PT|13.42|Mechanical phacofragmentation and aspiration of cataract by posterior route
C0176248|ICD9CM|AB|13.42|Post catarac frag/aspir
C0176249|ICD9CM|PT|13.43|Mechanical phacofragmentation and other aspiration of cataract
C0176249|ICD9CM|AB|13.43|Cataract frag/aspir NEC
C0176250|ICD9CM|PT|13.64|Discission of secondary membrane [after cataract]
C0176250|ICD9CM|AB|13.64|After-catar discission
C0176254|ICD9CM|PT|13.71|Insertion of intraocular lens prosthesis at time of cataract extraction, one-stage
C0176254|ICD9CM|AB|13.71|Insert lens at catar ext
C0176256|ICD9CM|HT|13.9|Other operations on lens
C0176258|ICD9CM|HT|14.1|Diagnostic procedures on retina, choroid, vitreous, and posterior chamber
C0176259|ICD9CM|PT|14.19|Other diagnostic procedures on retina, choroid, vitreous, and posterior chamber
C0176259|ICD9CM|AB|14.19|Dx proc post seg NEC
C0176260|ICD9CM|HT|14.2|Destruction of lesion of retina and choroid
C0176261|ICD9CM|PT|14.25|Destruction of chorioretinal lesion by photocoagulation of unspecified type
C0176261|ICD9CM|AB|14.25|Chorioret les p/coag NOS
C0176262|ICD9CM|PT|14.29|Other destruction of chorioretinal lesion
C0176262|ICD9CM|AB|14.29|Chorioret les destr NEC
C0176263|ICD9CM|HT|14.3|Repair of retinal tear
C0176264|ICD9CM|PT|14.31|Repair of retinal tear by diathermy
C0176264|ICD9CM|AB|14.31|Retinal tear diathermy
C0176265|ICD9CM|PT|14.32|Repair of retinal tear by cryotherapy
C0176265|ICD9CM|AB|14.32|Retinal tear cryotherapy
C0176266|ICD9CM|PT|14.34|Repair of retinal tear by laser photocoagulation
C0176266|ICD9CM|AB|14.34|Retinal tear laser coag
C0176267|ICD9CM|PT|14.35|Repair of retinal tear by photocoagulation of unspecified type
C0176267|ICD9CM|AB|14.35|Retina tear photocoa NOS
C0176268|ICD9CM|PT|14.39|Other repair of retinal tear
C0176268|ICD9CM|AB|14.39|Retinal tear repair NEC
C0176269|ICD9CM|HT|14.4|Repair of retinal detachment with scleral buckling and implant
C0176270|ICD9CM|HT|14.5|Other repair of retinal detachment
C0176270|ICD9CM|PT|14.59|Other repair of retinal detachment
C0176270|ICD9CM|AB|14.59|Repair retina detach NEC
C0176271|ICD9CM|PT|14.51|Repair of retinal detachment with diathermy
C0176271|ICD9CM|AB|14.51|Detach retina-diathermy
C0176276|ICD9CM|PT|14.72|Other removal of vitreous
C0176276|ICD9CM|AB|14.72|Vitreous removal NEC
C0176278|ICD9CM|PT|14.9|Other operations on retina, choroid, and posterior chamber
C0176278|ICD9CM|AB|14.9|Other post segment ops
C0176279|ICD9CM|HT|15.0|Diagnostic procedures on extraocular muscles or tendons
C0176280|ICD9CM|PT|15.01|Biopsy of extraocular muscle or tendon
C0176280|ICD9CM|AB|15.01|Extraoc musc-tend biopsy
C0176281|ICD9CM|PT|15.09|Other diagnostic procedures on extraocular muscles and tendons
C0176281|ICD9CM|AB|15.09|Extraoc musc dx proc NEC
C0176282|ICD9CM|HT|15.1|Operations on one extraocular muscle involving temporary detachment from globe
C0176283|ICD9CM|PT|15.12|Advancement of one extraocular muscle
C0176283|ICD9CM|AB|15.12|1 extraoc muscl advance
C0176284|ICD9CM|PT|15.19|Other operations on one extraocular muscle involving temporary detachment from globe
C0176284|ICD9CM|AB|15.19|Xtraoc mus op/detach NEC
C0176285|ICD9CM|HT|15.2|Other operations on one extraocular muscle
C0176285|ICD9CM|PT|15.29|Other operations on one extraocular muscle
C0176285|ICD9CM|AB|15.29|Op on 1 extraoc musc NEC
C0176287|ICD9CM|PT|15.4|Other operations on two or more extraocular muscles, one or both eyes
C0176287|ICD9CM|AB|15.4|Oth op on >l extraoc mus
C0176288|ICD9CM|PT|15.7|Repair of injury of extraocular muscle
C0176288|ICD9CM|AB|15.7|Extraoc musc inj repair
C0176289|ICD9CM|PT|15.9|Other operations on extraocular muscles and tendons
C0176289|ICD9CM|AB|15.9|Oth extraoc mus-tend op
C0176290|ICD9CM|PT|16.02|Orbitotomy with insertion of orbital implant
C0176290|ICD9CM|AB|16.02|Orbitotomy w implant
C0176291|MTH|PN|NOCODE|ORBITOTOMY NEC in ICD9CM
C0176291|ICD9CM|AB|16.09|Orbitotomy NEC
C0176291|ICD9CM|PT|16.09|Other orbitotomy
C0176292|ICD9CM|HT|16.2|Diagnostic procedures on orbit and eyeball
C0176293|ICD9CM|PT|16.29|Other diagnostic procedures on orbit and eyeball
C0176293|ICD9CM|AB|16.29|Eyebal/orbit dx proc NEC
C0176294|ICD9CM|PT|16.39|Other evisceration of eyeball
C0176294|ICD9CM|AB|16.39|Eyeball evisceration NEC
C0176295|ICD9CM|PT|16.42|Enucleation of eyeball with other synchronous implant
C0176295|ICD9CM|AB|16.42|Eye enuc w implant NEC
C0176296|ICD9CM|PT|16.49|Other enucleation of eyeball
C0176296|ICD9CM|AB|16.49|Eyeball enucleation NEC
C0176297|ICD9CM|PT|16.59|Other exenteration of orbit
C0176297|ICD9CM|AB|16.59|Orbital exenteration NEC
C0176299|ICD9CM|PT|16.64|Other revision of enucleation socket
C0176299|ICD9CM|AB|16.64|Enuc socket revis NEC
C0176300|ICD9CM|PT|16.65|Secondary graft to exenteration cavity
C0176300|ICD9CM|AB|16.65|2ndry exent cavity graft
C0176301|ICD9CM|PT|16.66|Other revision of exenteration cavity
C0176301|ICD9CM|AB|16.66|Revis exenter cavity NEC
C0176302|ICD9CM|PT|16.69|Other secondary procedures after removal of eyeball
C0176302|ICD9CM|AB|16.69|2nd op post eye rem NEC
C0176303|ICD9CM|HT|16.7|Removal of ocular or orbital implant
C0176304|ICD9CM|HT|16.8|Repair of injury of eyeball and orbit
C0176306|ICD9CM|PT|16.82|Repair of rupture of eyeball
C0176306|ICD9CM|AB|16.82|Repair eyeball rupture
C0176307|ICD9CM|PT|16.89|Other repair of injury of eyeball or orbit
C0176307|ICD9CM|AB|16.89|Eye/orbit inj repair NEC
C0176308|ICD9CM|HT|16.9|Other operations on orbit and eyeball
C0176310|ICD9CM|PT|16.98|Other operations on orbit
C0176310|ICD9CM|AB|16.98|Operation on orbit NEC
C0176311|ICD9CM|PT|16.99|Other operations on eyeball
C0176311|ICD9CM|AB|16.99|Operation on eyeball NEC
C0176312|ICD9CM|PT|18.09|Other incision of external ear
C0176312|ICD9CM|AB|18.09|External ear incis NEC
C0176314|ICD9CM|PT|18.19|Other diagnostic procedures on external ear
C0176314|ICD9CM|AB|18.19|Ext ear diagnos proc NEC
C0176315|ICD9CM|HT|18.2|Excision or destruction of lesion of external ear
C0176316|ICD9CM|PT|18.21|Excision of preauricular sinus
C0176316|ICD9CM|AB|18.21|Preauricular sinus excis
C0176317|ICD9CM|PT|18.29|Excision or destruction of other lesion of external ear
C0176317|ICD9CM|AB|18.29|Destruct ext ear les NEC
C0176318|ICD9CM|HT|18.3|Other excision of external ear
C0176318|ICD9CM|PT|18.39|Other excision of external ear
C0176318|ICD9CM|AB|18.39|Excis external ear NEC
C0176321|ICD9CM|HT|18.7|Other plastic repair of external ear
C0176321|ICD9CM|PT|18.79|Other plastic repair of external ear
C0176321|ICD9CM|AB|18.79|Plastic rep ext ear NEC
C0176322|ICD9CM|PT|18.71|Construction of auricle of ear
C0176322|ICD9CM|AB|18.71|Construction ear auricle
C0176323|ICD9CM|PT|18.9|Other operations on external ear
C0176323|ICD9CM|AB|18.9|Other ext ear operations
C0176324|ICD9CM|PT|19.19|Other stapedectomy
C0176324|ICD9CM|AB|19.19|Stapedectomy NEC
C0176325|ICD9CM|PT|19.21|Revision of stapedectomy with incus replacement
C0176325|ICD9CM|AB|19.21|Rev stapdec w incus repl
C0176326|ICD9CM|PT|19.29|Other revision of stapedectomy
C0176326|ICD9CM|AB|19.29|Stapedectomy revis NEC
C0176327|ICD9CM|PT|19.3|Other operations on ossicular chain
C0176327|ICD9CM|AB|19.3|Ossicular chain op NEC
C0176328|ICD9CM|HT|19.5|Other tympanoplasty
C0176331|ICD9CM|PT|19.54|Type IV tympanoplasty
C0176331|ICD9CM|AB|19.54|Type 4 tympanoplasty
C0176332|ICD9CM|PT|19.55|Type V tympanoplasty
C0176332|ICD9CM|AB|19.55|Type 5 tympanoplasty
C0176333|ICD9CM|PT|19.9|Other repair of middle ear
C0176333|ICD9CM|AB|19.9|Middle ear repair NEC
C0176334|ICD9CM|PT|20.09|Other myringotomy
C0176334|ICD9CM|AB|20.09|Myringotomy NEC
C0176335|ICD9CM|PT|20.1|Removal of tympanostomy tube
C0176335|ICD9CM|AB|20.1|Tympanostomy tube remove
C0176336|ICD9CM|HT|20.2|Incision of mastoid and middle ear
C0176338|ICD9CM|HT|20.3|Diagnostic procedures on middle and inner ear
C0176339|ICD9CM|PT|20.32|Biopsy of middle and inner ear
C0176339|ICD9CM|AB|20.32|Mid & inner ear biopsy
C0176340|ICD9CM|PT|20.39|Other diagnostic procedures on middle and inner ear
C0176340|ICD9CM|AB|20.39|Mid/in ear dx proc NEC
C0176341|ICD9CM|AB|20.41|Simple mastoidectomy
C0176341|ICD9CM|PT|20.41|Simple mastoidectomy
C0176342|MTH|PN|NOCODE|Mastoidectomy NEC in ICD9CM_2014
C0176342|ICD9CM|PT|20.49|Other mastoidectomy
C0176342|ICD9CM|AB|20.49|Mastoidectomy NEC
C0176343|ICD9CM|HT|20.5|Other excision of middle ear
C0176343|ICD9CM|PT|20.59|Other excision of middle ear
C0176343|ICD9CM|AB|20.59|Middle ear excision NEC
C0176345|ICD9CM|HT|20.7|Incision, excision, and destruction of inner ear
C0176346|ICD9CM|PT|20.79|Other incision, excision, and destruction of inner ear
C0176346|ICD9CM|AB|20.79|Inc/exc/destr in ear NEC
C0176348|ICD9CM|PT|20.97|Implantation or replacement of cochlear prosthetic device, single channel
C0176348|ICD9CM|AB|20.97|Imp/rep schan coch pros
C0176349|ICD9CM|PT|20.98|Implantation or replacement of cochlear prosthetic device, multiple channel
C0176349|ICD9CM|AB|20.98|Imp/rep mchan cochl pros
C0176350|ICD9CM|PT|21.01|Control of epistaxis by anterior nasal packing
C0176350|ICD9CM|AB|21.01|Ant nasal pack for epist
C0176354|ICD9CM|PT|21.06|Control of epistaxis by ligation of the external carotid artery
C0176354|ICD9CM|AB|21.06|Ext carot art lig-epist
C0176355|ICD9CM|PT|21.07|Control of epistaxis by excision of nasal mucosa and skin grafting of septum and lateral nasal wall
C0176355|ICD9CM|AB|21.07|Nasal sept grft-epistax
C0176356|ICD9CM|PT|21.09|Control of epistaxis by other means
C0176356|ICD9CM|AB|21.09|Epistaxis control NEC
C0176357|ICD9CM|HT|21.2|Diagnostic procedures on nose
C0176358|ICD9CM|PT|21.22|Biopsy of nose
C0176358|ICD9CM|AB|21.22|Nasal biopsy
C0176359|ICD9CM|PT|21.29|Other diagnostic procedures on nose
C0176359|ICD9CM|AB|21.29|Nasal dx proc NEC
C0176360|ICD9CM|HT|21.3|Local excision or destruction of lesion of nose
C0176361|ICD9CM|PT|21.30|Excision or destruction of lesion of nose, not otherwise specified
C0176361|ICD9CM|AB|21.30|Nasal lesion excis NOS
C0176362|ICD9CM|PT|21.31|Local excision or destruction of intranasal lesion
C0176362|ICD9CM|AB|21.31|Intranas les destruction
C0176363|ICD9CM|PT|21.32|Local excision or destruction of other lesion of nose
C0176363|ICD9CM|AB|21.32|Nasal les destruct NEC
C0176364|ICD9CM|AB|21.4|Resection of nose
C0176364|ICD9CM|PT|21.4|Resection of nose
C0176365|ICD9CM|PT|21.61|Turbinectomy by diathermy or cryosurgery
C0176365|ICD9CM|AB|21.61|Diather/cryo turbinectom
C0176367|ICD9CM|PT|21.69|Other turbinectomy
C0176367|ICD9CM|AB|21.69|Turbinectomy NEC
C0176368|ICD9CM|HT|21.7|Reduction of nasal fracture
C0176369|ICD9CM|HT|21.8|Repair and plastic operations on the nose
C0176370|ICD9CM|PT|21.82|Closure of nasal fistula
C0176370|ICD9CM|AB|21.82|Nasal fistula closure
C0176371|ICD9CM|AB|21.85|Augmentation rhinoplasty
C0176371|ICD9CM|PT|21.85|Augmentation rhinoplasty
C0176372|ICD9CM|PT|21.88|Other septoplasty
C0176372|ICD9CM|AB|21.88|Septoplasty NEC
C0176373|ICD9CM|PT|21.89|Other repair and plastic operations on nose
C0176373|ICD9CM|AB|21.89|Nasal repair NEC
C0176374|ICD9CM|HT|21.9|Other operations on nose
C0176374|ICD9CM|PT|21.99|Other operations on nose
C0176374|ICD9CM|AB|21.99|Nasal operation NEC
C0176375|ICD9CM|PT|22.01|Puncture of nasal sinus for aspiration or lavage
C0176375|ICD9CM|AB|22.01|Sinus punct for lavage
C0176376|ICD9CM|PT|22.02|Aspiration or lavage of nasal sinus through natural ostium
C0176376|ICD9CM|AB|22.02|Sinus lavage thru ostium
C0176377|ICD9CM|HT|22.1|Diagnostic procedures on nasal sinus
C0176378|ICD9CM|PT|22.11|Closed [endoscopic] [needle] biopsy of nasal sinus
C0176378|ICD9CM|AB|22.11|Closed nasal sinus bx
C0176379|ICD9CM|PT|22.12|Open biopsy of nasal sinus
C0176379|ICD9CM|AB|22.12|Open biopsy nasal sinus
C0176380|ICD9CM|PT|22.19|Other diagnostic procedures on nasal sinuses
C0176380|ICD9CM|AB|22.19|Nasal sinus dx proc NEC
C0176381|ICD9CM|HT|22.3|External maxillary antrotomy
C0176382|ICD9CM|PT|22.39|Other external maxillary antrotomy
C0176382|ICD9CM|AB|22.39|Ext maxillary antrot NEC
C0176383|ICD9CM|HT|22.4|Frontal sinusotomy and sinusectomy
C0176384|ICD9CM|HT|22.5|Other nasal sinusotomy
C0176385|ICD9CM|PT|22.53|Incision of multiple nasal sinuses
C0176385|ICD9CM|AB|22.53|Multiple sinus incision
C0176386|ICD9CM|HT|22.6|Other nasal sinusectomy
C0176387|ICD9CM|PT|22.60|Sinusectomy, not otherwise specified
C0176387|ICD9CM|AB|22.60|Sinusectomy NOS
C0176388|ICD9CM|PT|22.62|Excision of lesion of maxillary sinus with other approach
C0176388|ICD9CM|AB|22.62|Exc max sinus lesion NEC
C0176389|ICD9CM|PT|22.79|Other repair of nasal sinus
C0176389|ICD9CM|AB|22.79|Nasal sinus repair NEC
C0176390|ICD9CM|PT|22.9|Other operations on nasal sinuses
C0176390|ICD9CM|AB|22.9|Other nasal sinus ops
C0176391|ICD9CM|HT|23.0|Forceps extraction of tooth
C0176392|ICD9CM|PT|23.09|Extraction of other tooth
C0176392|ICD9CM|AB|23.09|Tooth extraction NEC
C0176394|ICD9CM|PT|23.11|Removal of residual root
C0176394|ICD9CM|AB|23.11|Residual root removal
C0176395|ICD9CM|PT|23.19|Other surgical extraction of tooth
C0176395|ICD9CM|AB|23.19|Surg tooth extract NEC
C0176396|ICD9CM|PT|23.2|Restoration of tooth by filling
C0176396|ICD9CM|AB|23.2|Tooth restor by filling
C0176397|ICD9CM|PT|23.3|Restoration of tooth by inlay
C0176397|ICD9CM|AB|23.3|Tooth restorat by inlay
C0176398|ICD9CM|HT|23.4|Other dental restoration
C0176398|ICD9CM|PT|23.49|Other dental restoration
C0176398|ICD9CM|AB|23.49|Dental restoration NEC
C0176399|ICD9CM|PT|23.42|Insertion of fixed bridge
C0176399|ICD9CM|AB|23.42|Fixed bridge insertion
C0176402|ICD9CM|PT|23.71|Root canal therapy with irrigation
C0176402|ICD9CM|AB|23.71|Root canal w irrigation
C0176403|ICD9CM|PT|23.72|Root canal therapy with apicoectomy
C0176403|ICD9CM|HT|23.7|Apicoectomy and root canal therapy
C0176403|ICD9CM|AB|23.72|Root canal w apicoectomy
C0176404|ICD9CM|PT|24.0|Incision of gum or alveolar bone
C0176404|ICD9CM|AB|24.0|Gum or alveolar incision
C0176405|ICD9CM|HT|24.1|Diagnostic procedures on teeth, gums, and alveoli
C0176406|ICD9CM|PT|24.11|Biopsy of gum
C0176406|ICD9CM|AB|24.11|Gum biopsy
C0176407|ICD9CM|PT|24.12|Biopsy of alveolus
C0176407|ICD9CM|AB|24.12|Alveolus biopsy
C0176408|ICD9CM|PT|24.19|Other diagnostic procedures on teeth, gums, and alveoli
C0176408|ICD9CM|AB|24.19|Tooth & gum dx proc NEC
C0176409|ICD9CM|HT|24.3|Other operations on gum
C0176409|ICD9CM|PT|24.39|Other operations on gum
C0176409|ICD9CM|AB|24.39|Gum operation NEC
C0176410|ICD9CM|AB|24.32|Suture of gum laceration
C0176410|ICD9CM|PT|24.32|Suture of laceration of gum
C0176411|ICD9CM|PT|24.4|Excision of dental lesion of jaw
C0176411|ICD9CM|AB|24.4|Exc of dental les of jaw
C0176412|ICD9CM|AB|24.6|Exposure of tooth
C0176412|ICD9CM|PT|24.6|Exposure of tooth
C0176413|ICD9CM|PT|24.7|Application of orthodontic appliance
C0176413|ICD9CM|AB|24.7|Orthodon applianc applic
C0176414|ICD9CM|PT|24.8|Other orthodontic operation
C0176414|ICD9CM|AB|24.8|Other orthodontic operat
C0176415|ICD9CM|HT|25.0|Diagnostic procedures on tongue
C0176416|ICD9CM|PT|25.01|Closed [needle] biopsy of tongue
C0176416|ICD9CM|AB|25.01|Closed biopsy of tongue
C0176417|ICD9CM|AB|25.02|Open biopsy of tongue
C0176417|ICD9CM|PT|25.02|Open biopsy of tongue
C0176418|ICD9CM|PT|25.09|Other diagnostic procedures on tongue
C0176418|ICD9CM|AB|25.09|Tongue dx procedure NEC
C0176419|ICD9CM|PT|25.1|Excision or destruction of lesion or tissue of tongue
C0176419|ICD9CM|AB|25.1|Destruction tongue les
C0176420|ICD9CM|HT|25.5|Repair of tongue and glossoplasty
C0176421|ICD9CM|PT|25.59|Other repair and plastic operations on tongue
C0176421|ICD9CM|AB|25.59|Repair of tongue NEC
C0176422|ICD9CM|HT|25.9|Other operations on tongue
C0176422|ICD9CM|PT|25.99|Other operations on tongue
C0176422|ICD9CM|AB|25.99|Tongue operation NEC
C0176423|ICD9CM|AB|25.94|Other glossotomy
C0176423|ICD9CM|PT|25.94|Other glossotomy
C0176424|ICD9CM|PT|26.0|Incision of salivary gland or duct
C0176424|ICD9CM|AB|26.0|Incis salivary glnd/duct
C0176425|ICD9CM|HT|26.1|Diagnostic procedures on salivary glands and ducts
C0176427|ICD9CM|PT|26.12|Open biopsy of salivary gland or duct
C0176427|ICD9CM|AB|26.12|Open bx saliv gland/duct
C0176428|ICD9CM|PT|26.19|Other diagnostic procedures on salivary glands and ducts
C0176428|ICD9CM|AB|26.19|Saliv glnd dx proc NEC
C0176430|ICD9CM|PT|26.29|Other excision of salivary gland lesion
C0176430|ICD9CM|AB|26.29|Saliv lesion excis NEC
C0176431|ICD9CM|HT|26.4|Repair of salivary gland or duct
C0176433|ICD9CM|PT|27.0|Drainage of face and floor of mouth
C0176433|ICD9CM|AB|27.0|Drain face & mouth floor
C0176434|ICD9CM|HT|27.2|Diagnostic procedures on oral cavity
C0176435|ICD9CM|PT|27.21|Biopsy of bony palate
C0176435|ICD9CM|AB|27.21|Bony palate biopsy
C0176436|ICD9CM|PT|27.29|Other diagnostic procedures on oral cavity
C0176436|ICD9CM|AB|27.29|Oral cavity dx proc NEC
C0176437|ICD9CM|HT|27.3|Excision of lesion or tissue of bony palate
C0176438|ICD9CM|PT|27.31|Local excision or destruction of lesion or tissue of bony palate
C0176438|ICD9CM|AB|27.31|Loc exc bony palate les
C0176439|ICD9CM|PT|27.32|Wide excision or destruction of lesion or tissue of bony palate
C0176439|ICD9CM|AB|27.32|Wide exc bony palate les
C0176440|ICD9CM|HT|27.4|Excision of other parts of mouth
C0176442|ICD9CM|PT|27.42|Wide excision of lesion of lip
C0176442|ICD9CM|AB|27.42|Wide excision of lip les
C0176443|ICD9CM|PT|27.43|Other excision of lesion or tissue of lip
C0176443|ICD9CM|AB|27.43|Excision of lip les NEC
C0176444|ICD9CM|PT|27.49|Other excision of mouth
C0176444|ICD9CM|AB|27.49|Excision of mouth NEC
C0176445|ICD9CM|PT|27.51|Suture of laceration of lip
C0176445|ICD9CM|AB|27.51|Suture of lip laceration
C0176446|ICD9CM|PT|27.52|Suture of laceration of other part of mouth
C0176446|ICD9CM|AB|27.52|Suture of mouth lac NEC
C0176447|ICD9CM|PT|27.55|Full-thickness skin graft to lip and mouth
C0176447|ICD9CM|AB|27.55|Full-thick grft to mouth
C0176448|ICD9CM|PT|27.56|Other skin graft to lip and mouth
C0176448|ICD9CM|AB|27.56|Skin graft to mouth NEC
C0176449|ICD9CM|PT|27.59|Other plastic repair of mouth
C0176449|ICD9CM|AB|27.59|Mouth repair NEC
C0176450|ICD9CM|PT|27.69|Other plastic repair of palate
C0176450|ICD9CM|AB|27.69|Oth plastic repair palat
C0176453|ICD9CM|PT|27.99|Other operations on oral cavity
C0176453|ICD9CM|AB|27.99|Oral cavity ops NEC
C0176454|ICD9CM|HT|28.1|Diagnostic procedures on tonsils and adenoids
C0176455|ICD9CM|PT|28.11|Biopsy of tonsils and adenoids
C0176455|ICD9CM|AB|28.11|Tonsil&adenoid biopsy
C0176456|ICD9CM|PT|28.19|Other diagnostic procedures on tonsils and adenoids
C0176456|ICD9CM|AB|28.19|Tonsil&adenoid dx op NEC
C0176457|ICD9CM|PT|28.91|Removal of foreign body from tonsil and adenoid by incision
C0176457|ICD9CM|AB|28.91|Incis to remov tonsil FB
C0176458|ICD9CM|PT|28.92|Excision of lesion of tonsil and adenoid
C0176458|ICD9CM|AB|28.92|Excis tonsil/adenoid les
C0176459|ICD9CM|HT|29.1|Diagnostic procedures on pharynx
C0176460|ICD9CM|PT|29.19|Other diagnostic procedures on pharynx
C0176460|ICD9CM|AB|29.19|Pharyngeal dx proc NEC
C0176461|ICD9CM|PT|29.2|Excision of branchial cleft cyst or vestige
C0176461|ICD9CM|AB|29.2|Exc branchial cleft cyst
C0176464|ICD9CM|PT|29.39|Other excision or destruction of lesion or tissue of pharynx
C0176464|ICD9CM|AB|29.39|Excis/destr les phar NEC
C0176465|ICD9CM|PT|29.4|Plastic operation on pharynx
C0176465|ICD9CM|AB|29.4|Plastic op on pharynx
C0176466|ICD9CM|PT|29.52|Closure of branchial cleft fistula
C0176466|ICD9CM|AB|29.52|Clos branch cleft fistul
C0176467|ICD9CM|PT|29.53|Closure of other fistula of pharynx
C0176467|ICD9CM|AB|29.53|Clos pharynx fistula NEC
C0176469|ICD9CM|HT|30.0|Excision or destruction of lesion or tissue of larynx
C0176471|ICD9CM|PT|30.09|Other excision or destruction of lesion or tissue of larynx
C0176471|ICD9CM|AB|30.09|Destruct larynx les NEC
C0176474|ICD9CM|AB|30.4|Radical laryngectomy
C0176474|ICD9CM|PT|30.4|Radical laryngectomy
C0176475|ICD9CM|PT|31.29|Other permanent tracheostomy
C0176475|ICD9CM|AB|31.29|Other perm tracheostomy
C0176476|ICD9CM|PT|31.3|Other incision of larynx or trachea
C0176476|ICD9CM|AB|31.3|Incis larynx trachea NEC
C0176477|ICD9CM|HT|31.4|Diagnostic procedures on larynx and trachea
C0176478|ICD9CM|PT|31.41|Tracheoscopy through artificial stoma
C0176478|ICD9CM|AB|31.41|Tracheoscopy thru stoma
C0176481|ICD9CM|PT|31.45|Open biopsy of larynx or trachea
C0176481|ICD9CM|AB|31.45|Opn bx larynx or trachea
C0176482|ICD9CM|PT|31.48|Other diagnostic procedures on larynx
C0176482|ICD9CM|AB|31.48|Oth larynx dx procedure
C0176483|ICD9CM|PT|31.49|Other diagnostic procedures on trachea
C0176483|ICD9CM|AB|31.49|Oth trachea dx procedure
C0176484|ICD9CM|PT|31.5|Local excision or destruction of lesion or tissue of trachea
C0176484|ICD9CM|AB|31.5|Local destruc trach les
C0176486|ICD9CM|PT|31.62|Closure of fistula of larynx
C0176486|ICD9CM|AB|31.62|Laryngeal fistula clos
C0176487|ICD9CM|PT|31.64|Repair of laryngeal fracture
C0176487|ICD9CM|AB|31.64|Laryngeal fx repair
C0176488|ICD9CM|PT|31.69|Other repair of larynx
C0176488|ICD9CM|AB|31.69|Other laryngeal repair
C0176489|ICD9CM|HT|31.7|Repair and plastic operations on trachea
C0176490|ICD9CM|PT|31.73|Closure of other fistula of trachea
C0176490|ICD9CM|AB|31.73|Trachea fistula clos NEC
C0176491|ICD9CM|PT|31.75|Reconstruction of trachea and construction of artificial larynx
C0176491|ICD9CM|AB|31.75|Tracheal reconstruction
C0176492|ICD9CM|PT|31.79|Other repair and plastic operations on trachea
C0176492|ICD9CM|AB|31.79|Other tracheal repair
C0176493|ICD9CM|PT|31.92|Lysis of adhesions of trachea or larynx
C0176493|ICD9CM|AB|31.92|Lysis trach/larynx adhes
C0176494|ICD9CM|PT|31.93|Replacement of laryngeal or tracheal stent
C0176494|ICD9CM|AB|31.93|Replace trac/laryn stent
C0176495|ICD9CM|PT|31.94|Injection of locally-acting therapeutic substance into trachea
C0176495|ICD9CM|AB|31.94|Tracheal injection
C0176497|ICD9CM|PT|31.98|Other operations on larynx
C0176497|ICD9CM|AB|31.98|Oth laryngeal operation
C0176499|ICD9CM|HT|32.0|Local excision or destruction of lesion or tissue of bronchus
C0176500|ICD9CM|PT|32.01|Endoscopic excision or destruction of lesion or tissue of bronchus
C0176500|ICD9CM|AB|32.01|Endosc destruc bronc les
C0176501|ICD9CM|PT|32.09|Other local excision or destruction of lesion or tissue of bronchus
C0176501|ICD9CM|AB|32.09|Other destruc bronc les
C0176502|ICD9CM|PT|32.1|Other excision of bronchus
C0176502|ICD9CM|AB|32.1|Other bronchial excision
C0176503|ICD9CM|HT|32.2|Local excision or destruction of lesion or tissue of lung
C0176504|ICD9CM|PT|32.28|Endoscopic excision or destruction of lesion or tissue of lung
C0176504|ICD9CM|AB|32.28|Endosc destruc lung les
C0176505|ICD9CM|PT|32.29|Other local excision or destruction of lesion or tissue of lung
C0176505|ICD9CM|AB|32.29|Destroy loc lung les NEC
C0176507|ICD9CM|PT|32.6|Radical dissection of thoracic structures
C0176507|ICD9CM|AB|32.6|Rad dissec thorac struct
C0176509|ICD9CM|HT|33.2|Diagnostic procedures on lung and bronchus
C0176510|ICD9CM|PT|33.21|Bronchoscopy through artificial stoma
C0176510|ICD9CM|AB|33.21|Bronchoscopy thru stoma
C0176511|ICD9CM|PT|33.24|Closed [endoscopic] biopsy of bronchus
C0176511|ICD9CM|AB|33.24|Closed bronchial biopsy
C0176512|ICD9CM|AB|33.26|Closed lung biopsy
C0176512|ICD9CM|PT|33.26|Closed [percutaneous] [needle] biopsy of lung
C0176513|ICD9CM|PT|33.27|Closed endoscopic biopsy of lung
C0176513|ICD9CM|AB|33.27|Clos endoscopic lung bx
C0176514|ICD9CM|PT|33.28|Open biopsy of lung
C0176514|ICD9CM|AB|33.28|Open lung biopsy
C0176515|ICD9CM|PT|33.29|Other diagnostic procedures on lung or bronchus
C0176515|ICD9CM|AB|33.29|Bronch/lung dx proc NEC
C0176516|ICD9CM|PT|33.31|Destruction of phrenic nerve for collapse of lung
C0176516|ICD9CM|AB|33.31|Destr phren-lung collaps
C0176517|ICD9CM|PT|33.33|Pneumoperitoneum for collapse of lung
C0176517|ICD9CM|AB|33.33|Pneumoperit-lung collaps
C0176518|ICD9CM|HT|33.4|Repair and plastic operation on lung and bronchus
C0176520|ICD9CM|PT|33.48|Other repair and plastic operations on bronchus
C0176520|ICD9CM|AB|33.48|Bronchial repair NEC
C0176521|ICD9CM|PT|33.49|Other repair and plastic operations on lung
C0176521|ICD9CM|AB|33.49|Lung repair NEC
C0176524|ICD9CM|AB|33.93|Puncture of lung
C0176524|ICD9CM|PT|33.93|Puncture of lung
C0176525|ICD9CM|PT|33.98|Other operations on bronchus
C0176525|ICD9CM|AB|33.98|Bronchial operation NEC
C0176527|ICD9CM|HT|34.0|Incision of chest wall and pleura
C0176530|ICD9CM|HT|34.2|Diagnostic procedures on chest wall, pleura, mediastinum, and diaphragm
C0176532|ICD9CM|PT|34.25|Closed [percutaneous] [needle] biopsy of mediastinum
C0176532|ICD9CM|AB|34.25|Clos mediastinal biopsy
C0176533|ICD9CM|PT|34.28|Other diagnostic procedures on chest wall, pleura, and diaphragm
C0176533|ICD9CM|AB|34.28|Dx procedure thorax NEC
C0176534|ICD9CM|PT|34.29|Other diagnostic procedures on mediastinum
C0176534|ICD9CM|AB|34.29|Dx proc mediastinum NEC
C0176536|ICD9CM|PT|34.4|Excision or destruction of lesion of chest wall
C0176536|ICD9CM|AB|34.4|Destruct chest wall les
C0176537|ICD9CM|AB|34.51|Decortication of lung
C0176537|ICD9CM|PT|34.51|Decortication of lung
C0176538|ICD9CM|PT|34.59|Other excision of pleura
C0176538|ICD9CM|AB|34.59|Other pleural excision
C0176539|ICD9CM|PT|34.73|Closure of other fistula of thorax
C0176539|ICD9CM|AB|34.73|Clos thoracic fistul NEC
C0176543|ICD9CM|PT|34.81|Excision of lesion or tissue of diaphragm
C0176543|ICD9CM|AB|34.81|Excise diaphragm lesion
C0176544|ICD9CM|PT|34.84|Other repair of diaphragm
C0176544|ICD9CM|AB|34.84|Other diaphragm repair
C0176545|ICD9CM|PT|34.89|Other operations on diaphragm
C0176545|ICD9CM|AB|34.89|Diaphragm operation NEC
C0176548|ICD9CM|PT|35.00|Closed heart valvotomy, unspecified valve
C0176548|ICD9CM|AB|35.00|Closed valvotomy NOS
C0176554|ICD9CM|PT|35.10|Open heart valvuloplasty without replacement, unspecified valve
C0176554|ICD9CM|AB|35.10|Open valvuloplasty NOS
C0176559|ICD9CM|PT|35.31|Operations on papillary muscle
C0176559|ICD9CM|AB|35.31|Papillary muscle ops
C0176562|ICD9CM|PT|35.39|Operations on other structures adjacent to valves of heart
C0176562|ICD9CM|AB|35.39|Tiss adj to valv ops NEC
C0176563|ICD9CM|HT|35.4|Production of septal defect in heart
C0176564|ICD9CM|PT|35.41|Enlargement of existing atrial septal defect
C0176564|ICD9CM|AB|35.41|Enlarge existing sep def
C0176566|ICD9CM|HT|35.5|Repair of atrial and ventricular septa with prosthesis
C0176567|ICD9CM|PT|35.50|Repair of unspecified septal defect of heart with prosthesis
C0176567|ICD9CM|AB|35.50|Prosth rep hrt septa NOS
C0176569|ICD9CM|PT|35.52|Repair of atrial septal defect with prosthesis, closed technique
C0176569|ICD9CM|AB|35.52|Pros repair atria def-cl
C0176570|ICD9CM|HT|35.6|Repair of atrial and ventricular septa with tissue graft
C0176572|ICD9CM|HT|35.7|Other and unspecified repair of atrial and ventricular septa
C0176573|ICD9CM|PT|35.70|Other and unspecified repair of unspecified septal defect of heart
C0176573|ICD9CM|AB|35.70|Heart septa repair NOS
C0176574|ICD9CM|PT|35.71|Other and unspecified repair of atrial septal defect
C0176574|ICD9CM|AB|35.71|Atria septa def rep NEC
C0176575|ICD9CM|PT|35.72|Other and unspecified repair of ventricular septal defect
C0176575|ICD9CM|AB|35.72|Ventr septa def rep NEC
C0176576|ICD9CM|PT|35.73|Other and unspecified repair of endocardial cushion defect
C0176576|ICD9CM|AB|35.73|Endocar cushion rep NEC
C0176577|ICD9CM|HT|35.8|Total repair of certain congenital cardiac anomalies
C0176578|ICD9CM|PT|35.82|Total repair of total anomalous pulmonary venous connection
C0176578|ICD9CM|AB|35.82|Total repair of tapvc
C0176579|ICD9CM|HT|35.9|Other operations on valves and septa of heart
C0176580|ICD9CM|PT|35.94|Creation of conduit between atrium and pulmonary artery
C0176580|ICD9CM|AB|35.94|Conduit artium-pulm art
C0176581|ICD9CM|PT|35.98|Other operations on septa of heart
C0176581|ICD9CM|AB|35.98|Other heart septa ops
C0176582|ICD9CM|PT|35.99|Other operations on valves of heart
C0176582|ICD9CM|AB|35.99|Other heart valve ops
C0176585|ICD9CM|PT|36.03|Open chest coronary artery angioplasty
C0176585|ICD9CM|AB|36.03|Open coronry angioplasty
C0176587|ICD9CM|PT|36.09|Other removal of coronary artery obstruction
C0176587|ICD9CM|AB|36.09|Rem of cor art obstr NEC
C0176589|ICD9CM|PT|36.19|Other bypass anastomosis for heart revascularization
C0176589|ICD9CM|AB|36.19|Hrt revas byps anas NEC
C0176590|ICD9CM|HT|36.3|Other heart revascularization
C0176590|ICD9CM|PT|36.39|Other heart revascularization
C0176590|ICD9CM|AB|36.39|Oth heart revascular
C0176591|ICD9CM|HT|36.9|Other operations on vessels of heart
C0176591|ICD9CM|PT|36.99|Other operations on vessels of heart
C0176591|ICD9CM|AB|36.99|Heart vessel op NEC
C0176593|ICD9CM|HT|37.1|Cardiotomy and pericardiotomy
C0176594|ICD9CM|HT|37.2|Diagnostic procedures on heart and pericardium
C0176595|ICD9CM|PT|37.29|Other diagnostic procedures on heart and pericardium
C0176595|ICD9CM|AB|37.29|Hrt/pericar dx proc NEC
C0176596|ICD9CM|HT|37.3|Pericardiectomy and excision of lesion of heart
C0176597|ICD9CM|PT|37.33|Excision or destruction of other lesion or tissue of heart, open approach
C0176597|ICD9CM|AB|37.33|Exc/dest hrt lesion open
C0176599|ICD9CM|PT|37.61|Implant of pulsation balloon
C0176599|ICD9CM|AB|37.61|Pulsation balloon implan
C0176602|ICD9CM|HT|37.7|Insertion, revision, replacement, and removal of leads; insertion of temporary pacemaker system; or revision of cardiac device pocket
C0176604|ICD9CM|PT|37.71|Initial insertion of transvenous lead [electrode] into ventricle
C0176604|ICD9CM|AB|37.71|Int insert lead in vent
C0176607|ICD9CM|PT|37.74|Insertion or replacement of epicardial lead [electrode] into epicardium
C0176607|ICD9CM|AB|37.74|Int or repl lead epicar
C0176611|ICD9CM|PT|37.78|Insertion of temporary transvenous pacemaker system
C0176611|ICD9CM|AB|37.78|Inser temp pacemaker sys
C0176613|ICD9CM|HT|37.8|Insertion, replacement, removal, and revision of pacemaker device
C0176614|ICD9CM|PT|37.80|Insertion of permanent pacemaker, initial or replacement, type of device not specified
C0176614|ICD9CM|AB|37.80|Int or repl perm pacemkr
C0176616|ICD9CM|PT|37.85|Replacement of any type pacemaker device with single-chamber device, not specified as rate responsive
C0176616|ICD9CM|AB|37.85|Repl pacem w 1-cham, non
C0176617|ICD9CM|PT|37.89|Revision or removal of pacemaker device
C0176617|ICD9CM|AB|37.89|Revise or remove pacemak
C0176619|ICD9CM|PT|37.94|Implantation or replacement of automatic cardioverter/defibrillator, total system [AICD]
C0176619|ICD9CM|AB|37.94|Implt/repl carddefib tot
C0176621|ICD9CM|PT|37.97|Replacement of automatic cardioverter/defibrillator lead(s) only
C0176621|ICD9CM|AB|37.97|Repl cardiodefib leads
C0176622|ICD9CM|PT|38.01|Incision of vessel, intracranial vessels
C0176622|ICD9CM|AB|38.01|Intracran vessel incis
C0176623|ICD9CM|PT|38.02|Incision of vessel, other vessels of head and neck
C0176623|ICD9CM|AB|38.02|Head/neck ves incis NEC
C0176624|ICD9CM|PT|38.03|Incision of vessel, upper limb vessels
C0176624|ICD9CM|AB|38.03|Upper limb vessel incis
C0176625|ICD9CM|PT|38.05|Incision of vessel, other thoracic vessels
C0176625|ICD9CM|AB|38.05|Thoracic vessel inc NEC
C0176629|ICD9CM|PT|38.12|Endarterectomy, other vessels of head and neck
C0176629|ICD9CM|AB|38.12|Head & neck endarter NEC
C0176631|ICD9CM|PT|38.15|Endarterectomy, other thoracic vessels
C0176631|ICD9CM|AB|38.15|Thoracic endarterectomy
C0176633|ICD9CM|PT|38.29|Other diagnostic procedures on blood vessels
C0176633|ICD9CM|AB|38.29|Blood vessel dx proc NEC
C0176634|ICD9CM|PT|38.31|Resection of vessel with anastomosis, intracranial vessels
C0176634|ICD9CM|AB|38.31|Intracran ves resec-anas
C0176635|ICD9CM|PT|38.32|Resection of vessel with anastomosis, other vessels of head and neck
C0176635|ICD9CM|AB|38.32|Head/neck ves resec-anas
C0176636|ICD9CM|PT|38.33|Resection of vessel with anastomosis, upper limb vessels
C0176636|ICD9CM|AB|38.33|Arm vessel resect/anast
C0176637|ICD9CM|PT|38.35|Resection of vessel with anastomosis, other thoracic vessels
C0176637|ICD9CM|AB|38.35|Thor vessel resect/anast
C0176639|ICD9CM|PT|38.41|Resection of vessel with replacement, intracranial vessels
C0176639|ICD9CM|AB|38.41|Intracran ves resec-repl
C0176640|ICD9CM|PT|38.42|Resection of vessel with replacement, other vessels of head and neck
C0176640|ICD9CM|AB|38.42|Head/neck ves resec-repl
C0176641|ICD9CM|PT|38.43|Resection of vessel with replacement, upper limb vessels
C0176641|ICD9CM|AB|38.43|Arm ves resect w replace
C0176642|ICD9CM|PT|38.45|Resection of vessel with replacement, thoracic vessels
C0176642|ICD9CM|AB|38.45|Resect thorac ves w repl
C0176643|ICD9CM|PT|38.47|Resection of vessel with replacement, abdominal veins
C0176643|ICD9CM|AB|38.47|Abd vein resect w replac
C0176644|ICD9CM|PT|38.48|Resection of vessel with replacement, lower limb arteries
C0176644|ICD9CM|AB|38.48|Leg artery resec w repla
C0176645|ICD9CM|PT|38.49|Resection of vessel with replacement, lower limb veins
C0176645|ICD9CM|AB|38.49|Leg vein resect w replac
C0176647|ICD9CM|PT|38.51|Ligation and stripping of varicose veins, intracranial vessels
C0176647|ICD9CM|AB|38.51|Intcran var v lig-strip
C0176648|ICD9CM|PT|38.52|Ligation and stripping of varicose veins, other vessels of head and neck
C0176648|ICD9CM|AB|38.52|Head/neck var v lig-str
C0176649|ICD9CM|PT|38.53|Ligation and stripping of varicose veins, upper limb vessels
C0176649|ICD9CM|AB|38.53|Arm varicose v lig-strip
C0176650|ICD9CM|PT|38.55|Ligation and stripping of varicose veins, other thoracic vessels
C0176650|ICD9CM|AB|38.55|Thorac var v lig-strip
C0176651|ICD9CM|PT|38.57|Ligation and stripping of varicose veins, abdominal veins
C0176651|ICD9CM|AB|38.57|Abd varicos v liga-strip
C0176652|ICD9CM|PT|38.59|Ligation and stripping of varicose veins, lower limb veins
C0176652|ICD9CM|AB|38.59|Leg varicos v liga-strip
C0176653|ICD9CM|PT|38.61|Other excision of vessels, intracranial vessels
C0176653|ICD9CM|AB|38.61|Intracran vessel excis
C0176654|ICD9CM|PT|38.62|Other excision of vessels, other vessels of head and neck
C0176654|ICD9CM|AB|38.62|Head/neck vessel excis
C0176655|ICD9CM|PT|38.63|Other excision of vessels, upper limb vessels
C0176655|ICD9CM|AB|38.63|Arm vessel excision
C0176656|ICD9CM|AB|38.64|Excision of aorta
C0176656|ICD9CM|PT|38.64|Other excision of vessels, aorta, abdominal
C0176657|ICD9CM|PT|38.65|Other excision of vessels, thoracic vessels
C0176657|ICD9CM|AB|38.65|Thoracic vessel excision
C0176658|ICD9CM|PT|38.66|Other excision of vessels, abdominal arteries
C0176658|ICD9CM|AB|38.66|Abdominal artery excis
C0176659|ICD9CM|PT|38.67|Other excision of vessels, abdominal veins
C0176659|ICD9CM|AB|38.67|Abdominal vein excision
C0176660|ICD9CM|PT|38.68|Other excision of vessels, lower limb arteries
C0176660|ICD9CM|AB|38.68|Leg artery excision
C0176661|ICD9CM|PT|38.69|Other excision of vessels, lower limb veins
C0176661|ICD9CM|AB|38.69|Leg vein excision
C0176662|ICD9CM|HT|38.8|Other surgical occlusion of vessels
C0176663|ICD9CM|PT|38.81|Other surgical occlusion of vessels, intracranial vessels
C0176663|ICD9CM|AB|38.81|Occlus intracran ves NEC
C0176664|ICD9CM|PT|38.82|Other surgical occlusion of vessels, other vessels of head and neck
C0176664|ICD9CM|AB|38.82|Occlus head/neck ves NEC
C0176665|ICD9CM|PT|38.83|Other surgical occlusion of vessels, upper limb vessels
C0176665|ICD9CM|AB|38.83|Occlude arm vessel NEC
C0176666|ICD9CM|PT|38.84|Other surgical occlusion of vessels, aorta, abdominal
C0176666|ICD9CM|AB|38.84|Occlude aorta NEC
C0176667|ICD9CM|PT|38.85|Other surgical occlusion of vessels, thoracic vessels
C0176667|ICD9CM|AB|38.85|Occlude thoracic ves NEC
C0176668|ICD9CM|PT|38.86|Other surgical occlusion of vessels, abdominal arteries
C0176668|ICD9CM|AB|38.86|Occlude abd artery NEC
C0176669|ICD9CM|PT|38.87|Other surgical occlusion of vessels, abdominal veins
C0176669|ICD9CM|AB|38.87|Occlude abd vein NEC
C0176670|ICD9CM|PT|38.88|Other surgical occlusion of vessels, lower limb arteries
C0176670|ICD9CM|AB|38.88|Occlude leg artery NEC
C0176671|ICD9CM|PT|38.89|Other surgical occlusion of vessels, lower limb veins
C0176671|ICD9CM|AB|38.89|Occlude leg vein NEC
C0176672|ICD9CM|HT|38.9|Puncture of vessel
C0176674|ICD9CM|PT|38.98|Other puncture of artery
C0176674|ICD9CM|AB|38.98|Arterial puncture NEC
C0176675|ICD9CM|PT|38.99|Other puncture of vein
C0176675|ICD9CM|AB|38.99|Venous puncture NEC
C0176677|ICD9CM|HT|39.2|Other shunt or vascular bypass
C0176678|ICD9CM|PT|39.22|Aorta-subclavian-carotid bypass
C0176678|ICD9CM|AB|39.22|Aorta-subclv-carot bypas
C0176679|ICD9CM|PT|39.23|Other intrathoracic vascular shunt or bypass
C0176679|ICD9CM|AB|39.23|Intrathoracic shunt NEC
C0176680|ICD9CM|AB|39.24|Aorta-renal bypass
C0176680|ICD9CM|PT|39.24|Aorta-renal bypass
C0176681|ICD9CM|PT|39.26|Other intra-abdominal vascular shunt or bypass
C0176681|ICD9CM|AB|39.26|Intra-abdomin shunt NEC
C0176682|ICD9CM|PT|39.28|Extracranial-intracranial (EC-IC) vascular bypass
C0176682|ICD9CM|AB|39.28|Extracran-intracr bypass
C0176683|ICD9CM|HT|39.3|Suture of vessel
C0176685|ICD9CM|PT|39.49|Other revision of vascular procedure
C0176685|ICD9CM|AB|39.49|Vasc proc revision NEC
C0176686|ICD9CM|PT|39.52|Other repair of aneurysm
C0176686|ICD9CM|AB|39.52|Aneurysm repair NEC
C0176688|ICD9CM|PT|39.56|Repair of blood vessel with tissue patch graft
C0176688|ICD9CM|AB|39.56|Repair vess w tis patch
C0176689|ICD9CM|PT|39.57|Repair of blood vessel with synthetic patch graft
C0176689|ICD9CM|AB|39.57|Rep vess w synth patch
C0176690|ICD9CM|PT|39.58|Repair of blood vessel with unspecified type of patch graft
C0176690|ICD9CM|AB|39.58|Repair vess w patch NOS
C0176692|ICD9CM|PT|39.66|Percutaneous cardiopulmonary bypass
C0176692|ICD9CM|AB|39.66|Per cardiopulmon bypass
C0176693|ICD9CM|HT|39.8|Operations on carotid body, carotid sinus and other vascular bodies
C0176694|ICD9CM|AB|39.91|Freeing of vessel
C0176694|ICD9CM|PT|39.91|Freeing of vessel
C0176695|ICD9CM|PT|39.94|Replacement of vessel-to-vessel cannula
C0176695|ICD9CM|AB|39.94|Replac ves-to-ves cannul
C0176696|ICD9CM|PT|40.0|Incision of lymphatic structures
C0176696|ICD9CM|AB|40.0|Incis lymphatic structur
C0176697|ICD9CM|HT|40.1|Diagnostic procedures on lymphatic structures
C0176698|ICD9CM|PT|40.19|Other diagnostic procedures on lymphatic structures
C0176698|ICD9CM|AB|40.19|Lymphatic diag proc NEC
C0176699|ICD9CM|HT|40.2|Simple excision of lymphatic structure
C0176700|ICD9CM|PT|40.29|Simple excision of other lymphatic structure
C0176700|ICD9CM|AB|40.29|Simp exc lymph struc NEC
C0176703|ICD9CM|HT|40.5|Radical excision of other lymph nodes
C0176703|ICD9CM|PT|40.59|Radical excision of other lymph nodes
C0176703|ICD9CM|AB|40.59|Rad node dissection NEC
C0176706|ICD9CM|PT|40.69|Other operations on thoracic duct
C0176706|ICD9CM|AB|40.69|Thoracic duct op NEC
C0176708|ICD9CM|PT|41.02|Allogeneic bone marrow transplant with purging
C0176708|ICD9CM|AB|41.02|Alo bone marrow trnsplnt
C0176709|ICD9CM|PT|41.03|Allogeneic bone marrow transplant without purging
C0176709|ICD9CM|AB|41.03|Allogrft bone marrow NOS
C0176710|ICD9CM|AB|41.1|Puncture of spleen
C0176710|ICD9CM|PT|41.1|Puncture of spleen
C0176711|ICD9CM|HT|41.3|Diagnostic procedures on bone marrow and spleen
C0176712|ICD9CM|PT|41.32|Closed [aspiration] [percutaneous] biopsy of spleen
C0176712|ICD9CM|AB|41.32|Closed spleen biopsy
C0176713|ICD9CM|PT|41.38|Other diagnostic procedures on bone marrow
C0176713|ICD9CM|AB|41.38|Marrow diagnost proc NEC
C0176714|ICD9CM|PT|41.39|Other diagnostic procedures on spleen
C0176714|ICD9CM|AB|41.39|Spleen diagnost proc NEC
C0176715|ICD9CM|HT|41.4|Excision or destruction of lesion or tissue of spleen
C0176717|ICD9CM|HT|41.9|Other operations on spleen and bone marrow
C0176720|ICD9CM|PT|41.99|Other operations on spleen
C0176720|ICD9CM|AB|41.99|Spleen operation NEC
C0176721|ICD9CM|PT|42.09|Other incision of esophagus
C0176721|ICD9CM|AB|42.09|Esophageal incision NEC
C0176722|ICD9CM|PT|42.19|Other external fistulization of esophagus
C0176722|ICD9CM|AB|42.19|Ext fistulizat esoph NEC
C0176723|ICD9CM|HT|42.2|Diagnostic procedures on esophagus
C0176724|ICD9CM|PT|42.21|Operative esophagoscopy by incision
C0176724|ICD9CM|AB|42.21|Esophagoscopy by incis
C0176725|ICD9CM|PT|42.23|Other esophagoscopy
C0176725|ICD9CM|AB|42.23|Esophagoscopy NEC
C0176727|ICD9CM|PT|42.29|Other diagnostic procedures on esophagus
C0176727|ICD9CM|AB|42.29|Esophageal dx proc NEC
C0176728|ICD9CM|HT|42.3|Local excision or destruction of lesion or tissue of esophagus
C0176729|ICD9CM|PT|42.31|Local excision of esophageal diverticulum
C0176729|ICD9CM|AB|42.31|Loc excis esoph divertic
C0176730|ICD9CM|PT|42.32|Local excision of other lesion or tissue of esophagus
C0176730|ICD9CM|AB|42.32|Local excis esophag NEC
C0176731|ICD9CM|PT|42.33|Endoscopic excision or destruction of lesion or tissue of esophagus
C0176731|ICD9CM|AB|42.33|Endosc destruc esoph les
C0176732|ICD9CM|PT|42.39|Other destruction of lesion or tissue of esophagus
C0176732|ICD9CM|AB|42.39|Destruct esophag les NEC
C0176733|ICD9CM|HT|42.5|Intrathoracic anastomosis of esophagus
C0176734|ICD9CM|PT|42.51|Intrathoracic esophagoesophagostomy
C0176734|ICD9CM|AB|42.51|Thorac esophagoesophagos
C0176735|ICD9CM|PT|42.54|Other intrathoracic esophagoenterostomy
C0176735|ICD9CM|AB|42.54|Thorac esophagoenter NEC
C0176736|ICD9CM|PT|42.56|Other intrathoracic esophagocolostomy
C0176736|ICD9CM|AB|42.56|Thorac esophagocolos NEC
C0176737|ICD9CM|PT|42.59|Other intrathoracic anastomosis of esophagus
C0176737|ICD9CM|AB|42.59|Thorac esophag anast NEC
C0176738|ICD9CM|HT|42.6|Antesternal anastomosis of esophagus
C0176739|ICD9CM|PT|42.61|Antesternal esophagoesophagostomy
C0176739|ICD9CM|AB|42.61|Stern esophagoesophagost
C0176740|ICD9CM|PT|42.62|Antesternal esophagogastrostomy
C0176740|ICD9CM|AB|42.62|Stern esophagogastrostom
C0176741|ICD9CM|PT|42.63|Antesternal esophageal anastomosis with interposition of small bowel
C0176741|ICD9CM|AB|42.63|Stern sm bowel interpos
C0176742|ICD9CM|PT|42.64|Other antesternal esophagoenterostomy
C0176742|ICD9CM|AB|42.64|Stern esophagoenter NEC
C0176743|ICD9CM|PT|42.65|Antesternal esophageal anastomosis with interposition of colon
C0176743|ICD9CM|AB|42.65|Stern lg bowel interpos
C0176744|ICD9CM|PT|42.66|Other antesternal esophagocolostomy
C0176744|ICD9CM|AB|42.66|Stern esophagocolos NEC
C0176745|ICD9CM|PT|42.68|Other antesternal esophageal anastomosis with interposition
C0176745|ICD9CM|AB|42.68|Stern interposition NEC
C0176746|ICD9CM|PT|42.69|Other antesternal anastomosis of esophagus
C0176746|ICD9CM|AB|42.69|Stern esophag anast NEC
C0176747|ICD9CM|PT|42.81|Insertion of permanent tube into esophagus
C0176747|ICD9CM|AB|42.81|Insert perm tube esophag
C0176748|ICD9CM|PT|42.86|Production of subcutaneous tunnel without esophageal anastomosis
C0176748|ICD9CM|AB|42.86|Prod subq tunnel no anas
C0176749|ICD9CM|PT|42.87|Other graft of esophagus
C0176749|ICD9CM|AB|42.87|Esophageal graft NEC
C0176750|ICD9CM|HT|42.9|Other operations on esophagus
C0176751|ICD9CM|PT|43.11|Percutaneous [endoscopic] gastrostomy [PEG]
C0176751|ICD9CM|AB|43.11|Percu endosc gastrostomy
C0176752|ICD9CM|AB|43.19|Other gastrostomy
C0176752|ICD9CM|PT|43.19|Other gastrostomy
C0176753|ICD9CM|HT|43.4|Local excision or destruction of lesion or tissue of stomach
C0176754|ICD9CM|PT|43.41|Endoscopic excision or destruction of lesion or tissue of stomach
C0176754|ICD9CM|AB|43.41|Endosc destr stomach les
C0176755|ICD9CM|PT|43.42|Local excision of other lesion or tissue of stomach
C0176755|ICD9CM|AB|43.42|Local gastr excision NEC
C0176756|ICD9CM|PT|43.49|Other destruction of lesion or tissue of stomach
C0176756|ICD9CM|AB|43.49|Local gastr destruct NEC
C0176757|ICD9CM|PT|43.5|Partial gastrectomy with anastomosis to esophagus
C0176757|ICD9CM|AB|43.5|Proximal gastrectomy
C0176758|ICD9CM|PT|43.6|Partial gastrectomy with anastomosis to duodenum
C0176758|ICD9CM|AB|43.6|Distal gastrectomy
C0176759|ICD9CM|PT|43.99|Other total gastrectomy
C0176759|ICD9CM|AB|43.99|Total gastrectomy NEC
C0176760|ICD9CM|PT|44.03|Other selective vagotomy
C0176760|ICD9CM|AB|44.03|Selective vagotomy NEC
C0176761|ICD9CM|HT|44.1|Diagnostic procedures on stomach
C0176763|ICD9CM|PT|44.19|Other diagnostic procedures on stomach
C0176763|ICD9CM|AB|44.19|Gastric diagnos proc NEC
C0176764|ICD9CM|PT|44.21|Dilation of pylorus by incision
C0176764|ICD9CM|AB|44.21|Dilate pylorus, incision
C0176765|ICD9CM|AB|44.29|Other pyloroplasty
C0176765|ICD9CM|PT|44.29|Other pyloroplasty
C0176766|ICD9CM|HT|44.4|Control of hemorrhage and suture of ulcer of stomach or duodenum
C0176767|ICD9CM|AB|44.40|Suture peptic ulcer NOS
C0176767|ICD9CM|PT|44.40|Suture of peptic ulcer, not otherwise specified
C0176768|ICD9CM|PT|44.41|Suture of gastric ulcer site
C0176768|ICD9CM|AB|44.41|Sut gastric ulcer site
C0176770|ICD9CM|PT|44.43|Endoscopic control of gastric or duodenal bleeding
C0176770|ICD9CM|AB|44.43|Endosc control gast hem
C0176771|ICD9CM|PT|44.44|Transcatheter embolization for gastric or duodenal bleeding
C0176771|ICD9CM|AB|44.44|Transcath embo gast hem
C0176772|ICD9CM|PT|44.49|Other control of hemorrhage of stomach or duodenum
C0176772|ICD9CM|AB|44.49|Other control gast hem
C0176773|ICD9CM|PT|44.5|Revision of gastric anastomosis
C0176773|ICD9CM|AB|44.5|Revision gastric anastom
C0176775|ICD9CM|PT|44.63|Closure of other gastric fistula
C0176775|ICD9CM|AB|44.63|Close gastric fistul NEC
C0176776|ICD9CM|PT|44.66|Other procedures for creation of esophagogastric sphincteric competence
C0176776|ICD9CM|AB|44.66|Creat esophagastr sphinc
C0176777|ICD9CM|PT|44.92|Intraoperative manipulation of stomach
C0176777|ICD9CM|AB|44.92|Intraop gastric manipul
C0176780|ICD9CM|PT|45.02|Other incision of small intestine
C0176780|ICD9CM|AB|45.02|Small bowel incision NEC
C0176781|ICD9CM|HT|45.1|Diagnostic procedures on small intestine
C0176782|ICD9CM|PT|45.11|Transabdominal endoscopy of small intestine
C0176782|ICD9CM|AB|45.11|Transab sm bowel endosc
C0176784|ICD9CM|PT|45.16|Esophagogastroduodenoscopy [EGD] with closed biopsy
C0176784|ICD9CM|AB|45.16|Egd with closed biopsy
C0176785|ICD9CM|PT|45.19|Other diagnostic procedures on small intestine
C0176785|ICD9CM|AB|45.19|Sm bowel dx proc NEC
C0176789|ICD9CM|PT|45.28|Other diagnostic procedures on large intestine
C0176789|ICD9CM|AB|45.28|Lg bowel dx proced NEC
C0176790|ICD9CM|HT|45.3|Local excision or destruction of lesion or tissue of small intestine
C0176791|ICD9CM|PT|45.30|Endoscopic excision or destruction of lesion of duodenum
C0176791|ICD9CM|AB|45.30|Endosc destru duoden les
C0176792|ICD9CM|PT|45.31|Other local excision of lesion of duodenum
C0176792|ICD9CM|AB|45.31|Oth excise duodenum les
C0176793|ICD9CM|PT|45.32|Other destruction of lesion of duodenum
C0176793|ICD9CM|AB|45.32|Destruct duoden les NEC
C0176794|ICD9CM|PT|45.33|Local excision of lesion or tissue of small intestine, except duodenum
C0176794|ICD9CM|AB|45.33|Local excis sm bowel NEC
C0176795|ICD9CM|PT|45.34|Other destruction of lesion of small intestine, except duodenum
C0176795|ICD9CM|AB|45.34|Destr sm bowel les NEC
C0176796|ICD9CM|HT|45.4|Local excision or destruction of lesion or tissue of large intestine
C0176797|ICD9CM|PT|45.41|Excision of lesion or tissue of large intestine
C0176797|ICD9CM|AB|45.41|Excise lg intestine les
C0176799|ICD9CM|PT|45.49|Other destruction of lesion of large intestine
C0176799|ICD9CM|AB|45.49|Destruc lg bowel les NEC
C0176801|ICD9CM|PT|45.51|Isolation of segment of small intestine
C0176801|ICD9CM|AB|45.51|Sm bowel segment isolat
C0176802|ICD9CM|PT|45.52|Isolation of segment of large intestine
C0176802|ICD9CM|AB|45.52|Lg bowel segment isolat
C0176803|ICD9CM|HT|45.6|Other excision of small intestine
C0176804|ICD9CM|PT|45.62|Other partial resection of small intestine
C0176804|ICD9CM|AB|45.62|Part sm bowel resect NEC
C0176806|ICD9CM|HT|45.8|Total intra-abdominal colectomy
C0176808|ICD9CM|PT|45.93|Other small-to-large intestinal anastomosis
C0176808|ICD9CM|AB|45.93|Small-to-large bowel NEC
C0176809|ICD9CM|PT|45.95|Anastomosis to anus
C0176809|ICD9CM|AB|45.95|Anal anastomosis
C0176811|ICD9CM|PT|46.23|Other permanent ileostomy
C0176811|ICD9CM|AB|46.23|Permanent ileostomy NEC
C0176812|ICD9CM|PT|46.31|Delayed opening of other enterostomy
C0176812|ICD9CM|AB|46.31|Delay opening enterostom
C0176813|ICD9CM|PT|46.32|Percutaneous (endoscopic) jejunostomy [PEJ]
C0176813|ICD9CM|AB|46.32|Percu endosc jejunostomy
C0176816|ICD9CM|PT|46.43|Other revision of stoma of large intestine
C0176816|ICD9CM|AB|46.43|Lg bowel stoma revis NEC
C0176817|ICD9CM|PT|46.62|Other fixation of small intestine
C0176817|ICD9CM|AB|46.62|Small bowel fixation NEC
C0176818|ICD9CM|PT|46.64|Other fixation of large intestine
C0176818|ICD9CM|AB|46.64|Large bowel fixation NEC
C0176819|ICD9CM|HT|46.7|Other repair of intestine
C0176819|ICD9CM|PT|46.79|Other repair of intestine
C0176819|ICD9CM|AB|46.79|Repair of intestine NEC
C0176821|ICD9CM|PT|46.73|Suture of laceration of small intestine, except duodenum
C0176821|ICD9CM|AB|46.73|Small bowel suture NEC
C0176822|ICD9CM|PT|46.74|Closure of fistula of small intestine, except duodenum
C0176822|ICD9CM|AB|46.74|Close sm bowel fist NEC
C0176823|ICD9CM|PT|46.75|Suture of laceration of large intestine
C0176823|ICD9CM|AB|46.75|Suture lg bowel lacerat
C0176824|ICD9CM|HT|46.8|Dilation and manipulation of intestine
C0176825|ICD9CM|AB|46.85|Dilation of intestine
C0176825|ICD9CM|PT|46.85|Dilation of intestine
C0176826|ICD9CM|AB|46.91|Myotomy of sigmoid colon
C0176826|ICD9CM|PT|46.91|Myotomy of sigmoid colon
C0176827|ICD9CM|PT|46.92|Myotomy of other parts of colon
C0176827|ICD9CM|AB|46.92|Myotomy of colon NEC
C0176828|ICD9CM|PT|46.95|Local perfusion of small intestine
C0176828|ICD9CM|AB|46.95|Local sm bowel perfusion
C0176829|ICD9CM|PT|46.96|Local perfusion of large intestine
C0176829|ICD9CM|AB|46.96|Local lg bowel perfusion
C0176830|ICD9CM|PT|47.2|Drainage of appendiceal abscess
C0176830|ICD9CM|AB|47.2|Drain appendiceal absc
C0176831|ICD9CM|HT|47.9|Other operations on appendix
C0176831|ICD9CM|PT|47.99|Other operations on appendix
C0176831|ICD9CM|AB|47.99|Appendiceal ops NEC
C0176832|ICD9CM|HT|48.2|Diagnostic procedures on rectum, rectosigmoid and perirectal tissue
C0176833|ICD9CM|PT|48.21|Transabdominal proctosigmoidoscopy
C0176833|ICD9CM|AB|48.21|Transab proctosigmoidosc
C0176835|ICD9CM|AB|48.25|Open rectal biopsy
C0176835|ICD9CM|PT|48.25|Open biopsy of rectum
C0176836|ICD9CM|PT|48.26|Biopsy of perirectal tissue
C0176836|ICD9CM|AB|48.26|Perirectal tissue biopsy
C0176837|ICD9CM|PT|48.29|Other diagnostic procedures on rectum, rectosigmoid and perirectal tissue
C0176837|ICD9CM|AB|48.29|Rect/perirect dx op NEC
C0176838|ICD9CM|HT|48.3|Local excision or destruction of lesion or tissue of rectum
C0176839|ICD9CM|PT|48.31|Radical electrocoagulation of rectal lesion or tissue
C0176839|ICD9CM|AB|48.31|Rad electrocoag-rect les
C0176840|ICD9CM|PT|48.32|Other electrocoagulation of rectal lesion or tissue
C0176840|ICD9CM|AB|48.32|Electrocoag rect les NEC
C0176841|ICD9CM|PT|48.33|Destruction of rectal lesion or tissue by laser
C0176841|ICD9CM|AB|48.33|Laser destruc rectal les
C0176842|ICD9CM|PT|48.34|Destruction of rectal lesion or tissue by cryosurgery
C0176842|ICD9CM|AB|48.34|Cryosurg destr rect les
C0176843|ICD9CM|PT|48.35|Local excision of rectal lesion or tissue
C0176843|ICD9CM|AB|48.35|Local excis rectal les
C0176844|ICD9CM|HT|48.4|Pull-through resection of rectum
C0176845|ICD9CM|PT|48.49|Other pull-through resection of rectum
C0176845|ICD9CM|AB|48.49|Pull-thru rect resec NEC
C0176847|ICD9CM|HT|48.6|Other resection of rectum
C0176847|ICD9CM|PT|48.69|Other resection of rectum
C0176847|ICD9CM|AB|48.69|Rectal resection NEC
C0176848|ICD9CM|PT|48.62|Anterior resection of rectum with synchronous colostomy
C0176848|ICD9CM|AB|48.62|Ant rect resect w colost
C0176849|ICD9CM|PT|48.63|Other anterior resection of rectum
C0176849|ICD9CM|AB|48.63|Anterior rect resect NEC
C0176850|ICD9CM|PT|48.65|Duhamel resection of rectum
C0176850|ICD9CM|AB|48.65|Duhamel rectal resection
C0176851|ICD9CM|PT|48.73|Closure of other rectal fistula
C0176851|ICD9CM|AB|48.73|Close rectal fist NEC
C0176853|ICD9CM|PT|48.76|Other proctopexy
C0176853|ICD9CM|AB|48.76|Proctopexy NEC
C0176854|ICD9CM|PT|48.79|Other repair of rectum
C0176854|ICD9CM|AB|48.79|Repair of rectum NEC
C0176855|ICD9CM|HT|48.8|Incision or excision of perirectal tissue or lesion
C0176856|ICD9CM|HT|48.9|Other operations on rectum and perirectal tissue
C0176856|ICD9CM|PT|48.99|Other operations on rectum and perirectal tissue
C0176856|ICD9CM|AB|48.99|Rectal perirect op NEC
C0176857|ICD9CM|HT|49.0|Incision or excision of perianal tissue
C0176858|ICD9CM|PT|49.01|Incision of perianal abscess
C0176858|ICD9CM|AB|49.01|Incis perianal abscess
C0176859|ICD9CM|PT|49.02|Other incision of perianal tissue
C0176859|ICD9CM|AB|49.02|Perianal incision NEC
C0176860|ICD9CM|PT|49.04|Other excision of perianal tissue
C0176860|ICD9CM|AB|49.04|Perianal excision NEC
C0176861|ICD9CM|HT|49.1|Incision or excision of anal fistula
C0176862|ICD9CM|HT|49.2|Diagnostic procedures on anus and perianal tissue
C0176863|ICD9CM|PT|49.29|Other diagnostic procedures on anus and perianal tissue
C0176863|ICD9CM|AB|49.29|Anal/perian dx proc NEC
C0176864|ICD9CM|PT|49.39|Other local excision or destruction of lesion or tissue of anus
C0176864|ICD9CM|HT|49.3|Local excision or destruction of other lesion or tissue of anus
C0176864|ICD9CM|AB|49.39|Other destruc anus les
C0176865|ICD9CM|PT|49.31|Endoscopic excision or destruction of lesion or tissue of anus
C0176865|ICD9CM|AB|49.31|Endosc destruc anus les
C0176866|ICD9CM|HT|49.4|Procedures on hemorrhoids
C0176867|ICD9CM|PT|49.41|Reduction of hemorrhoids
C0176867|ICD9CM|AB|49.41|Hemorrhoid reduction
C0176869|ICD9CM|PT|49.49|Other procedures on hemorrhoids
C0176869|ICD9CM|AB|49.49|Hemorrhoid procedure NEC
C0176870|ICD9CM|HT|49.5|Division of anal sphincter
C0176871|ICD9CM|PT|49.59|Other anal sphincterotomy
C0176871|ICD9CM|AB|49.59|Anal sphincterotomy NEC
C0176872|ICD9CM|AB|49.6|Excision of anus
C0176872|ICD9CM|PT|49.6|Excision of anus
C0176873|ICD9CM|PT|49.79|Other repair of anal sphincter
C0176873|ICD9CM|AB|49.79|Anal sphinct repair NEC
C0176874|ICD9CM|HT|49.9|Other operations on anus
C0176874|ICD9CM|PT|49.99|Other operations on anus
C0176874|ICD9CM|AB|49.99|Anal operation NEC
C0176876|ICD9CM|PT|49.93|Other incision of anus
C0176876|ICD9CM|AB|49.93|Anal incision NEC
C0176877|ICD9CM|PT|49.94|Reduction of anal prolapse
C0176877|ICD9CM|AB|49.94|Reduction anal prolapse
C0176879|ICD9CM|PT|50.11|Closed (percutaneous) [needle] biopsy of liver
C0176879|ICD9CM|AB|50.11|Closed liver biopsy
C0176880|ICD9CM|PT|50.19|Other diagnostic procedures on liver
C0176880|ICD9CM|AB|50.19|Hepatic dx proc NEC
C0176881|ICD9CM|HT|50.2|Local excision or destruction of liver tissue or lesion
C0176882|ICD9CM|PT|50.21|Marsupialization of lesion of liver
C0176882|ICD9CM|AB|50.21|Marsupializat liver les
C0176883|ICD9CM|PT|50.29|Other destruction of lesion of liver
C0176883|ICD9CM|AB|50.29|Destruc hepatic les NEC
C0176884|ICD9CM|PT|50.51|Auxiliary liver transplant
C0176884|ICD9CM|AB|50.51|Auxiliary liver transpl
C0176885|ICD9CM|PT|50.61|Closure of laceration of liver
C0176885|ICD9CM|AB|50.61|Closure liver lacerat
C0176886|ICD9CM|PT|50.69|Other repair of liver
C0176886|ICD9CM|AB|50.69|Liver repair NEC
C0176887|ICD9CM|HT|50.9|Other operations on liver
C0176887|ICD9CM|PT|50.99|Other operations on liver
C0176887|ICD9CM|AB|50.99|Liver operation NEC
C0176888|ICD9CM|PT|50.92|Extracorporeal hepatic assistance
C0176888|ICD9CM|AB|50.92|Extracorpor hepat Assis
C0176889|ICD9CM|PT|50.93|Localized perfusion of liver
C0176889|ICD9CM|AB|50.93|Local perfusion liver
C0176890|ICD9CM|PT|50.94|Other injection of therapeutic substance into liver
C0176890|ICD9CM|AB|50.94|Hepatic injection NEC
C0176891|ICD9CM|HT|51.0|Cholecystotomy and cholecystostomy
C0176893|ICD9CM|AB|51.02|Trocar cholecystostomy
C0176893|ICD9CM|PT|51.02|Trocar cholecystostomy
C0176894|ICD9CM|PT|51.04|Other cholecystotomy
C0176894|ICD9CM|AB|51.04|Cholecystotomy NEC
C0176895|ICD9CM|HT|51.1|Diagnostic procedures on biliary tract
C0176899|ICD9CM|PT|51.13|Open biopsy of gallbladder or bile ducts
C0176899|ICD9CM|AB|51.13|Open biliary tract bx
C0176900|ICD9CM|PT|51.14|Other closed [endoscopic] biopsy of biliary duct or sphincter of Oddi
C0176900|ICD9CM|AB|51.14|Clo endosc bx bile duct
C0176901|ICD9CM|PT|51.19|Other diagnostic procedures on biliary tract
C0176901|ICD9CM|AB|51.19|Biliary tr dx proc NEC
C0176902|ICD9CM|HT|51.3|Anastomosis of gallbladder or bile duct
C0176904|ICD9CM|PT|51.35|Other gallbladder anastomosis
C0176904|ICD9CM|AB|51.35|Gallbladder anastom NEC
C0176905|ICD9CM|PT|51.39|Other bile duct anastomosis
C0176905|ICD9CM|AB|51.39|Bile duct anastomos NEC
C0176906|ICD9CM|HT|51.4|Incision of bile duct for relief of obstruction
C0176908|ICD9CM|PT|51.42|Common duct exploration for relief of other obstruction
C0176908|ICD9CM|AB|51.42|Cde for obstruction NEC
C0176909|ICD9CM|PT|51.49|Incision of other bile ducts for relief of obstruction
C0176909|ICD9CM|AB|51.49|Incis obstr bile duc NEC
C0176910|ICD9CM|HT|51.5|Other incision of bile duct
C0176912|ICD9CM|HT|51.6|Local excision or destruction of lesion or tissue of biliary ducts and sphincter of Oddi
C0176914|ICD9CM|PT|51.63|Other excision of common duct
C0176914|ICD9CM|AB|51.63|Common duct excis NEC
C0176915|ICD9CM|PT|51.64|Endoscopic excision or destruction of lesion of biliary ducts or sphincter of Oddi
C0176915|ICD9CM|AB|51.64|Endosc destru bile les
C0176916|ICD9CM|PT|51.69|Excision of other bile duct
C0176916|ICD9CM|AB|51.69|Bile duct excision NEC
C0176917|ICD9CM|PT|51.79|Repair of other bile ducts
C0176917|ICD9CM|AB|51.79|Bile duct repair NEC
C0176918|ICD9CM|HT|51.8|Other operations on biliary ducts and sphincter of Oddi
C0176919|ICD9CM|PT|51.82|Pancreatic sphincterotomy
C0176919|ICD9CM|AB|51.82|Pancreat sphincterotom
C0176920|ICD9CM|PT|51.83|Pancreatic sphincteroplasty
C0176920|ICD9CM|AB|51.83|Pancreat sphincteroplas
C0176921|ICD9CM|PT|51.84|Endoscopic dilation of ampulla and biliary duct
C0176921|ICD9CM|AB|51.84|Endosc dilation ampulla
C0176923|ICD9CM|PT|51.86|Endoscopic insertion of nasobiliary drainage tube
C0176923|ICD9CM|AB|51.86|Endosc inser nasobil tub
C0176924|ICD9CM|PT|51.87|Endoscopic insertion of stent (tube) into bile duct
C0176924|ICD9CM|AB|51.87|Endosc inser stent bile
C0176925|ICD9CM|PT|51.88|Endoscopic removal of stone(s) from biliary tract
C0176925|ICD9CM|AB|51.88|Endosc remove bile stone
C0176926|ICD9CM|PT|51.89|Other operations on sphincter of Oddi
C0176926|ICD9CM|AB|51.89|Sphinct of oddi op NEC
C0176928|ICD9CM|PT|51.93|Closure of other biliary fistula
C0176928|ICD9CM|AB|51.93|Clos biliary fistul NEC
C0176929|ICD9CM|PT|51.98|Other percutaneous procedures on biliary tract
C0176929|ICD9CM|AB|51.98|Oth perc proc bil trct
C0176930|ICD9CM|PT|52.01|Drainage of pancreatic cyst by catheter
C0176930|ICD9CM|AB|52.01|Cath drain-pancreat cyst
C0176931|ICD9CM|PT|52.09|Other pancreatotomy
C0176931|ICD9CM|AB|52.09|Pancreatotomy NEC
C0176932|ICD9CM|HT|52.1|Diagnostic procedures on pancreas
C0176935|ICD9CM|PT|52.14|Closed [endoscopic] biopsy of pancreatic duct
C0176935|ICD9CM|AB|52.14|Clo endosc bx pancre duc
C0176936|ICD9CM|PT|52.19|Other diagnostic procedures on pancreas
C0176936|ICD9CM|AB|52.19|Pancreatic dx proc NEC
C0176937|ICD9CM|HT|52.2|Local excision or destruction of pancreas and pancreatic duct
C0176938|ICD9CM|PT|52.21|Endoscopic excision or destruction of lesion or tissue of pancreatic duct
C0176938|ICD9CM|AB|52.21|Endosc destr pancrea les
C0176939|ICD9CM|PT|52.22|Other excision or destruction of lesion or tissue of pancreas or pancreatic duct
C0176939|ICD9CM|AB|52.22|Other destru pancrea les
C0176940|ICD9CM|AB|52.52|Distal pancreatectomy
C0176940|ICD9CM|PT|52.52|Distal pancreatectomy
C0176941|ICD9CM|PT|52.53|Radical subtotal pancreatectomy
C0176941|ICD9CM|AB|52.53|Rad subtot pancreatectom
C0176945|ICD9CM|PT|52.92|Cannulation of pancreatic duct
C0176945|ICD9CM|AB|52.92|Cannulation pancrea duc
C0176948|ICD9CM|PT|52.95|Other repair of pancreas
C0176948|ICD9CM|AB|52.95|Pancreatic repair NEC
C0176955|ICD9CM|PT|53.29|Other unilateral femoral herniorrhaphy
C0176955|ICD9CM|AB|53.29|Unil femor hern rep NEC
C0176957|ICD9CM|PT|53.39|Other bilateral femoral herniorrhaphy
C0176957|ICD9CM|AB|53.39|Bil fem hern repair NEC
C0176959|ICD9CM|HT|53.5|Repair of other hernia of anterior abdominal wall (without graft or prosthesis)
C0176961|ICD9CM|PT|53.59|Repair of other hernia of anterior abdominal wall
C0176961|ICD9CM|AB|53.59|Abd wall hern repair NEC
C0176962|ICD9CM|HT|53.6|Repair of other hernia of anterior abdominal wall with graft or prosthesis
C0176967|ICD9CM|AB|53.9|Other hernia repair
C0176967|ICD9CM|PT|53.9|Other hernia repair
C0176969|ICD9CM|HT|54.2|Diagnostic procedures of abdominal region
C0176972|ICD9CM|PT|54.29|Other diagnostic procedures on abdominal region
C0176972|ICD9CM|AB|54.29|Abd region dx proc NEC
C0176973|ICD9CM|PT|54.3|Excision or destruction of lesion or tissue of abdominal wall or umbilicus
C0176973|ICD9CM|AB|54.3|Destruct abd wall lesion
C0176974|ICD9CM|PT|54.4|Excision or destruction of peritoneal tissue
C0176974|ICD9CM|AB|54.4|Destruct peritoneal tiss
C0176977|ICD9CM|PT|54.63|Other suture of abdominal wall
C0176977|ICD9CM|AB|54.63|Abd wall suture NEC
C0176978|ICD9CM|HT|54.7|Other repair of abdominal wall and peritoneum
C0176979|ICD9CM|PT|54.72|Other repair of abdominal wall
C0176979|ICD9CM|AB|54.72|Abdomen wall repair NEC
C0176980|ICD9CM|PT|54.73|Other repair of peritoneum
C0176980|ICD9CM|AB|54.73|Peritoneal repair NEC
C0176981|ICD9CM|PT|54.74|Other repair of omentum
C0176981|ICD9CM|AB|54.74|Omental repair NEC
C0176982|ICD9CM|PT|54.75|Other repair of mesentery
C0176982|ICD9CM|AB|54.75|Mesenteric repair NEC
C0176984|ICD9CM|HT|55.0|Nephrotomy and nephrostomy
C0176985|ICD9CM|PT|55.04|Percutaneous nephrostomy with fragmentation
C0176985|ICD9CM|AB|55.04|Percu nephrostmy w frag
C0176986|ICD9CM|HT|55.1|Pyelotomy and pyelostomy
C0176989|ICD9CM|HT|55.2|Diagnostic procedures on kidney
C0176990|ICD9CM|AB|55.22|Pyeloscopy
C0176990|ICD9CM|PT|55.22|Pyeloscopy
C0176992|ICD9CM|PT|55.29|Other diagnostic procedures on kidney
C0176992|ICD9CM|AB|55.29|Renal diagnost proc NEC
C0176993|ICD9CM|HT|55.3|Local excision or destruction of lesion or tissue of kidney
C0176994|ICD9CM|PT|55.31|Marsupialization of kidney lesion
C0176994|ICD9CM|AB|55.31|Renal les marsupializat
C0176995|ICD9CM|PT|55.39|Other local destruction or excision of renal lesion or tissue
C0176995|ICD9CM|AB|55.39|Loc destr renal les NEC
C0176996|ICD9CM|HT|55.5|Complete nephrectomy
C0176997|ICD9CM|PT|55.53|Removal of transplanted or rejected kidney
C0176997|ICD9CM|AB|55.53|Rejected kidney nephrect
C0176998|ICD9CM|PT|55.81|Suture of laceration of kidney
C0176998|ICD9CM|AB|55.81|Suture kidney laceration
C0176999|ICD9CM|PT|55.82|Closure of nephrostomy and pyelostomy
C0176999|ICD9CM|AB|55.82|Close nephrost & pyelost
C0177000|ICD9CM|PT|55.83|Closure of other fistula of kidney
C0177000|ICD9CM|AB|55.83|Close renal fistula NEC
C0177002|ICD9CM|AB|55.86|Renal anastomosis
C0177002|ICD9CM|PT|55.86|Anastomosis of kidney
C0177004|ICD9CM|PT|55.96|Other injection of therapeutic substance into kidney
C0177004|ICD9CM|AB|55.96|Renal injection NEC
C0177005|ICD9CM|PT|55.97|Implantation or replacement of mechanical kidney
C0177005|ICD9CM|AB|55.97|Implant mechanic kidney
C0177006|ICD9CM|HT|56.3|Diagnostic procedures on ureter
C0177007|ICD9CM|PT|56.32|Closed percutaneous biopsy of ureter
C0177007|ICD9CM|AB|56.32|Closed ureteral biopsy
C0177008|ICD9CM|PT|56.33|Closed endoscopic biopsy of ureter
C0177008|ICD9CM|AB|56.33|Clos endosc ureteral bx
C0177009|ICD9CM|PT|56.34|Open biopsy of ureter
C0177009|ICD9CM|AB|56.34|Open ureteral biopsy
C0177011|ICD9CM|PT|56.39|Other diagnostic procedures on ureter
C0177011|ICD9CM|AB|56.39|Ureteral dx procedur NEC
C0177012|ICD9CM|HT|56.5|Cutaneous uretero-ileostomy
C0177014|ICD9CM|HT|56.6|Other external urinary diversion
C0177015|ICD9CM|PT|56.62|Revision of other cutaneous ureterostomy
C0177015|ICD9CM|AB|56.62|Revis cutan ureteros NEC
C0177018|ICD9CM|PT|56.84|Closure of other fistula of ureter
C0177018|ICD9CM|AB|56.84|Close ureter fistula NEC
C0177019|ICD9CM|PT|56.86|Removal of ligature from ureter
C0177019|ICD9CM|AB|56.86|Remove ureteral ligature
C0177020|ICD9CM|PT|56.89|Other repair of ureter
C0177020|ICD9CM|AB|56.89|Repair of ureter NEC
C0177022|ICD9CM|HT|57.1|Cystotomy and cystostomy
C0177023|ICD9CM|PT|57.11|Percutaneous aspiration of bladder
C0177023|ICD9CM|AB|57.11|Percutan bladder aspirat
C0177024|ICD9CM|PT|57.12|Lysis of intraluminal adhesions with incision into bladder
C0177024|ICD9CM|AB|57.12|Cystotomy & adhesiolysis
C0177025|ICD9CM|AB|57.17|Percutaneous cystostomy
C0177025|ICD9CM|PT|57.17|Percutaneous cystostomy
C0177026|ICD9CM|PT|57.18|Other suprapubic cystostomy
C0177026|ICD9CM|AB|57.18|Other suprapu cystostomy
C0177027|ICD9CM|PT|57.19|Other cystotomy
C0177027|ICD9CM|AB|57.19|Cystotomy NEC
C0177028|ICD9CM|PT|57.22|Revision or closure of vesicostomy
C0177028|ICD9CM|AB|57.22|Revise clo vesicostomy
C0177029|ICD9CM|HT|57.3|Diagnostic procedures on bladder
C0177030|ICD9CM|PT|57.31|Cystoscopy through artificial stoma
C0177030|ICD9CM|AB|57.31|Cystoscopy thru stoma
C0177032|ICD9CM|PT|57.34|Open biopsy of bladder
C0177032|ICD9CM|AB|57.34|Open bladder biopsy
C0177033|ICD9CM|PT|57.39|Other diagnostic procedures on bladder
C0177033|ICD9CM|AB|57.39|Bladder diagnos proc NEC
C0177034|ICD9CM|HT|57.4|Transurethral excision or destruction of bladder tissue
C0177035|ICD9CM|PT|57.41|Transurethral lysis of intraluminal adhesions
C0177035|ICD9CM|AB|57.41|Tu adhesiolysis bladder
C0177036|ICD9CM|PT|57.49|Other transurethral excision or destruction of lesion or tissue of bladder
C0177036|ICD9CM|AB|57.49|Tu destruc bladd les NEC
C0177037|ICD9CM|HT|57.5|Other excision or destruction of bladder tissue
C0177038|ICD9CM|AB|57.51|Excision of urachus
C0177038|ICD9CM|PT|57.51|Excision of urachus
C0177039|ICD9CM|PT|57.59|Open excision or destruction of other lesion or tissue of bladder
C0177039|ICD9CM|AB|57.59|Bladder les destruct NEC
C0177041|ICD9CM|PT|57.79|Other total cystectomy
C0177041|ICD9CM|AB|57.79|Total cystectomy NEC
C0177044|ICD9CM|PT|57.84|Repair of other fistula of bladder
C0177044|ICD9CM|AB|57.84|Vesic fistula repair NEC
C0177045|ICD9CM|PT|57.88|Other anastomosis of bladder
C0177045|ICD9CM|AB|57.88|Bladder anastomosis NEC
C0177046|ICD9CM|PT|57.89|Other repair of bladder
C0177046|ICD9CM|HT|57.8|Other repair of urinary bladder
C0177046|ICD9CM|AB|57.89|Bladder repair NEC
C0177047|ICD9CM|AB|57.91|Bladder sphincterotomy
C0177047|ICD9CM|PT|57.91|Sphincterotomy of bladder
C0177049|ICD9CM|PT|57.94|Insertion of indwelling urinary catheter
C0177049|ICD9CM|AB|57.94|Insert indwelling cath
C0177050|ICD9CM|PT|57.95|Replacement of indwelling urinary catheter
C0177050|ICD9CM|AB|57.95|Replace indwelling cath
C0177051|ICD9CM|PT|57.96|Implantation of electronic bladder stimulator
C0177051|ICD9CM|AB|57.96|Implant bladder stimulat
C0177052|ICD9CM|PT|57.97|Replacement of electronic bladder stimulator
C0177052|ICD9CM|AB|57.97|Replace bladder stimulat
C0177053|ICD9CM|HT|58.2|Diagnostic procedures on urethra
C0177054|ICD9CM|PT|58.22|Other urethroscopy
C0177054|ICD9CM|AB|58.22|Urethroscopy NEC
C0177055|ICD9CM|PT|58.29|Other diagnostic procedures on urethra and periurethral tissue
C0177055|ICD9CM|AB|58.29|Urethral dx proc NEC
C0177056|ICD9CM|HT|58.3|Excision or destruction of lesion or tissue of urethra
C0177057|ICD9CM|PT|58.31|Endoscopic excision or destruction of lesion or tissue of urethra
C0177057|ICD9CM|AB|58.31|Endosc destr urethra les
C0177058|ICD9CM|PT|58.39|Other local excision or destruction of lesion or tissue of urethra
C0177058|ICD9CM|AB|58.39|Other destru urethra les
C0177059|ICD9CM|PT|58.43|Closure of other fistula of urethra
C0177059|ICD9CM|AB|58.43|Close ureth fistula NEC
C0177060|ICD9CM|PT|58.45|Repair of hypospadias or epispadias
C0177060|ICD9CM|AB|58.45|Hypo-epispadius repair
C0177061|ICD9CM|PT|58.46|Other reconstruction of urethra
C0177061|ICD9CM|AB|58.46|Ureth reconstruction NEC
C0177063|ICD9CM|PT|58.49|Other repair of urethra
C0177063|ICD9CM|AB|58.49|Urethral repair NEC
C0177065|ICD9CM|HT|59.0|Dissection of retroperitoneal tissue
C0177067|ICD9CM|PT|59.02|Other lysis of perirenal or periureteral adhesions
C0177067|ICD9CM|AB|59.02|Periren adhesiolys NEC
C0177068|ICD9CM|PT|59.09|Other incision of perirenal or periureteral tissue
C0177068|ICD9CM|AB|59.09|Periren/ureter incis NEC
C0177069|ICD9CM|PT|59.19|Other incision of perivesical tissue
C0177069|ICD9CM|AB|59.19|Perivesical incision NEC
C0177070|ICD9CM|HT|59.2|Diagnostic procedures on perirenal and perivesical tissue
C0177071|ICD9CM|PT|59.21|Biopsy of perirenal or perivesical tissue
C0177071|ICD9CM|AB|59.21|Periren/ureteral biopsy
C0177072|ICD9CM|PT|59.29|Other diagnostic procedures on perirenal tissue, perivesical tissue, and retroperitoneum
C0177072|ICD9CM|AB|59.29|Periren/uret dx proc NEC
C0177074|ICD9CM|PT|59.5|Retropubic urethral suspension
C0177074|ICD9CM|AB|59.5|Retropubic ureth suspens
C0177076|ICD9CM|HT|59.7|Other repair of urinary stress incontinence
C0177076|ICD9CM|PT|59.79|Other repair of urinary stress incontinence
C0177076|ICD9CM|AB|59.79|Urin incontin repair NEC
C0177077|ICD9CM|PT|59.91|Excision of perirenal or perivesical tissue
C0177077|ICD9CM|AB|59.91|Periren/vesicle excision
C0177078|ICD9CM|PT|59.92|Other operations on perirenal or perivesical tissue
C0177078|ICD9CM|AB|59.92|Periren/vesicle op NEC
C0177080|ICD9CM|HT|60.1|Diagnostic procedures on prostate and seminal vesicles
C0177082|ICD9CM|PT|60.12|Open biopsy of prostate
C0177082|ICD9CM|AB|60.12|Open prostatic biopsy
C0177084|ICD9CM|PT|60.14|Open biopsy of seminal vesicles
C0177084|ICD9CM|AB|60.14|Open seminal vesicles bx
C0177085|ICD9CM|PT|60.15|Biopsy of periprostatic tissue
C0177085|ICD9CM|AB|60.15|Periprostatic biopsy
C0177086|ICD9CM|PT|60.18|Other diagnostic procedures on prostate and periprostatic tissue
C0177086|ICD9CM|AB|60.18|Prostatic dx proced NEC
C0177087|ICD9CM|PT|60.19|Other diagnostic procedures on seminal vesicles
C0177087|ICD9CM|AB|60.19|Semin ves dx proced NEC
C0177088|ICD9CM|PT|60.61|Local excision of lesion of prostate
C0177088|ICD9CM|AB|60.61|Los excis prostatic les
C0177091|ICD9CM|HT|60.8|Incision or excision of periprostatic tissue
C0177092|ICD9CM|PT|60.91|Percutaneous aspiration of prostate
C0177092|ICD9CM|AB|60.91|Percut prostatic aspirat
C0177094|ICD9CM|PT|60.94|Control of (postoperative) hemorrhage of prostate
C0177094|ICD9CM|AB|60.94|Control prostate hemorr
C0177096|ICD9CM|PT|61.0|Incision and drainage of scrotum and tunica vaginalis
C0177096|ICD9CM|AB|61.0|Scrotum & tunica i & d
C0177097|ICD9CM|HT|61.1|Diagnostic procedures on scrotum and tunica vaginalis
C0177098|ICD9CM|PT|61.11|Biopsy of scrotum or tunica vaginalis
C0177098|ICD9CM|AB|61.11|Scrotum & tunica biopsy
C0177101|ICD9CM|PT|61.3|Excision or destruction of lesion or tissue of scrotum
C0177101|ICD9CM|AB|61.3|Scrotal les destruction
C0177102|ICD9CM|HT|61.4|Repair of scrotum and tunica vaginalis
C0177105|ICD9CM|PT|61.49|Other repair of scrotum and tunica vaginalis
C0177105|ICD9CM|AB|61.49|Scrotum/tunic repair NEC
C0177106|ICD9CM|PT|61.91|Percutaneous aspiration of tunica vaginalis
C0177106|ICD9CM|AB|61.91|Percut tunica aspiration
C0177107|ICD9CM|PT|61.92|Excision of lesion of tunica vaginalis other than hydrocele
C0177107|ICD9CM|AB|61.92|Excision tunica les NEC
C0177108|ICD9CM|HT|62.1|Diagnostic procedures on testes
C0177109|ICD9CM|PT|62.11|Closed [percutaneous] [needle] biopsy of testis
C0177109|ICD9CM|AB|62.11|Closed testicular biopsy
C0177110|ICD9CM|PT|62.12|Open biopsy of testis
C0177110|ICD9CM|AB|62.12|Open testicular biopsy
C0177111|ICD9CM|PT|62.19|Other diagnostic procedures on testes
C0177111|ICD9CM|AB|62.19|Testes dx procedure NEC
C0177112|ICD9CM|PT|62.2|Excision or destruction of testicular lesion
C0177112|ICD9CM|AB|62.2|Testicular les destruct
C0177114|ICD9CM|PT|62.69|Other repair of testis
C0177114|ICD9CM|AB|62.69|Testicular repair NEC
C0177115|ICD9CM|PT|62.91|Aspiration of testis
C0177115|ICD9CM|AB|62.91|Aspiration of testes
C0177116|ICD9CM|HT|63.0|Diagnostic procedures on spermatic cord, epididymis, and vas deferens
C0177117|ICD9CM|PT|63.01|Biopsy of spermatic cord, epididymis, or vas deferens
C0177117|ICD9CM|AB|63.01|Spermatic cord/vas biops
C0177118|ICD9CM|PT|63.09|Other diagnostic procedures on spermatic cord, epididymis, and vas deferens
C0177118|ICD9CM|AB|63.09|Spermat cord/vas dx NEC
C0177119|ICD9CM|PT|63.1|Excision of varicocele and hydrocele of spermatic cord
C0177119|ICD9CM|AB|63.1|Exc spermatic varicocele
C0177120|ICD9CM|PT|63.2|Excision of cyst of epididymis
C0177120|ICD9CM|AB|63.2|Excise epididymis cyst
C0177121|ICD9CM|PT|63.3|Excision of other lesion or tissue of spermatic cord and epididymis
C0177121|ICD9CM|AB|63.3|Excise cord/epid les NEC
C0177124|ICD9CM|PT|63.52|Reduction of torsion of testis or spermatic cord
C0177124|ICD9CM|AB|63.52|Reduction torsion testes
C0177125|ICD9CM|PT|63.53|Transplantation of spermatic cord
C0177125|ICD9CM|AB|63.53|Transplant spermat cord
C0177126|ICD9CM|PT|63.59|Other repair of spermatic cord and epididymis
C0177126|ICD9CM|AB|63.59|Cord & epidid repair NEC
C0177127|ICD9CM|HT|63.7|Vasectomy and ligation of vas deferens
C0177129|ICD9CM|HT|63.8|Repair of vas deferens and epididymis
C0177130|ICD9CM|PT|63.81|Suture of laceration of vas deferens and epididymis
C0177130|ICD9CM|AB|63.81|Suture vas & epidid lac
C0177133|ICD9CM|PT|63.89|Other repair of vas deferens and epididymis
C0177133|ICD9CM|AB|63.89|Vas & epididy repair NEC
C0177134|ICD9CM|HT|63.9|Other operations on spermatic cord, epididymis, and vas deferens
C0177135|ICD9CM|PT|63.99|Other operations on spermatic card, epididymis, and vas deferens
C0177135|ICD9CM|AB|63.99|Cord/epid/vas ops NEC
C0177136|ICD9CM|HT|64.1|Diagnostic procedures on the penis
C0177137|ICD9CM|PT|64.11|Biopsy of penis
C0177137|ICD9CM|AB|64.11|Penile biopsy
C0177138|ICD9CM|PT|64.19|Other diagnostic procedures on penis
C0177138|ICD9CM|AB|64.19|Penile diagnost proc NEC
C0177139|ICD9CM|PT|64.2|Local excision or destruction of lesion of penis
C0177139|ICD9CM|AB|64.2|Local excis penile les
C0177140|ICD9CM|HT|64.4|Repair and plastic operation on penis
C0177141|ICD9CM|AB|64.42|Release of chordee
C0177141|ICD9CM|PT|64.42|Release of chordee
C0177142|ICD9CM|AB|64.43|Construction of penis
C0177142|ICD9CM|PT|64.43|Construction of penis
C0177143|ICD9CM|PT|64.49|Other repair of penis
C0177143|ICD9CM|AB|64.49|Penile repair NEC
C0177145|ICD9CM|PT|64.91|Dorsal or lateral slit of prepuce
C0177145|ICD9CM|AB|64.91|Dorsal/lat slit prepuce
C0177147|ICD9CM|PT|64.95|Insertion or replacement of non-inflatable penile prosthesis
C0177147|ICD9CM|AB|64.95|Ins noninfl penis prosth
C0177149|ICD9CM|PT|64.97|Insertion or replacement of inflatable penile prosthesis
C0177149|ICD9CM|AB|64.97|Ins inflate penis prosth
C0177150|ICD9CM|PT|64.98|Other operations on penis
C0177150|ICD9CM|AB|64.98|Penile operation NEC
C0177152|ICD9CM|PT|65.11|Aspiration biopsy of ovary
C0177152|ICD9CM|AB|65.11|Ovarian aspirat biopsy
C0177153|ICD9CM|PT|65.12|Other biopsy of ovary
C0177153|ICD9CM|AB|65.12|Ovarian biopsy NEC
C0177154|ICD9CM|PT|65.19|Other diagnostic procedures on ovaries
C0177154|ICD9CM|AB|65.19|Ovarian dx procedure NEC
C0177155|ICD9CM|HT|65.2|Local excision or destruction of ovarian lesion or tissue
C0177156|ICD9CM|PT|65.22|Wedge resection of ovary
C0177156|ICD9CM|AB|65.22|Ovarian wedge resection
C0177157|ICD9CM|PT|65.29|Other local excision or destruction of ovary
C0177157|ICD9CM|AB|65.29|Local destr ova les NEC
C0177161|ICD9CM|PT|65.79|Other repair of ovary
C0177161|ICD9CM|AB|65.79|Repair of ovary NEC
C0177163|ICD9CM|HT|66.1|Diagnostic procedures on fallopian tubes
C0177164|ICD9CM|PT|66.19|Other diagnostic procedures on fallopian tubes
C0177164|ICD9CM|AB|66.19|Fallop tube dx proc NEC
C0177165|ICD9CM|HT|66.2|Bilateral endoscopic destruction or occlusion of fallopian tubes
C0177166|ICD9CM|PT|66.29|Other bilateral endoscopic destruction or occlusion of fallopian tubes
C0177166|ICD9CM|AB|66.29|Bilat endos occ tube NEC
C0177167|ICD9CM|PT|66.31|Other bilateral ligation and crushing of fallopian tubes
C0177167|ICD9CM|AB|66.31|Bilat tubal crushing NEC
C0177168|ICD9CM|PT|66.32|Other bilateral ligation and division of fallopian tubes
C0177168|ICD9CM|AB|66.32|Bilat tubal division NEC
C0177169|ICD9CM|PT|66.4|Total unilateral salpingectomy
C0177169|ICD9CM|AB|66.4|Total unilat salpingect
C0177172|ICD9CM|PT|66.52|Removal of remaining fallopian tube
C0177172|ICD9CM|AB|66.52|Remove solitary fal tube
C0177173|ICD9CM|HT|66.6|Other salpingectomy
C0177175|ICD9CM|PT|66.62|Salpingectomy with removal of tubal pregnancy
C0177175|ICD9CM|AB|66.62|Remov tube & ectop preg
C0177176|ICD9CM|PT|66.69|Other partial salpingectomy
C0177176|ICD9CM|AB|66.69|Partial salpingectom NEC
C0177177|ICD9CM|PT|66.71|Simple suture of fallopian tube
C0177177|ICD9CM|AB|66.71|Simpl suture fallop tube
C0177178|ICD9CM|AB|66.74|Salpingo-uterostomy
C0177178|ICD9CM|PT|66.74|Salpingo-uterostomy
C0177179|ICD9CM|PT|66.79|Other repair of fallopian tube
C0177179|ICD9CM|AB|66.79|Fallop tube repair NEC
C0177180|ICD9CM|PT|66.92|Unilateral destruction or occlusion of fallopian tube
C0177180|ICD9CM|AB|66.92|Unilat fallop tube destr
C0177181|ICD9CM|PT|66.93|Implantation or replacement of prosthesis of fallopian tube
C0177181|ICD9CM|AB|66.93|Impl fallop tube prosth
C0177182|ICD9CM|PT|66.94|Removal of prosthesis of fallopian tube
C0177182|ICD9CM|AB|66.94|Remov fallop tube prosth
C0177183|ICD9CM|PT|66.95|Insufflation of therapeutic agent into fallopian tubes
C0177183|ICD9CM|AB|66.95|Blow therapeut into tube
C0177185|ICD9CM|HT|67.1|Diagnostic procedures on cervix
C0177186|ICD9CM|PT|67.12|Other cervical biopsy
C0177186|ICD9CM|AB|67.12|Cervical biopsy NEC
C0177187|ICD9CM|PT|67.19|Other diagnostic procedures on cervix
C0177187|ICD9CM|AB|67.19|Cervical dx procedur NEC
C0177189|ICD9CM|HT|67.3|Other excision or destruction of lesion or tissue of cervix
C0177189|ICD9CM|PT|67.39|Other excision or destruction of lesion or tissue of cervix
C0177189|ICD9CM|AB|67.39|Cervical les destruc NEC
C0177190|ICD9CM|PT|67.31|Marsupialization of cervical cyst
C0177190|ICD9CM|AB|67.31|Cervical cyst marsupial
C0177192|ICD9CM|PT|67.33|Destruction of lesion of cervix by cryosurgery
C0177192|ICD9CM|AB|67.33|Cervical les cryotherapy
C0177195|ICD9CM|PT|68.11|Digital examination of uterus
C0177195|ICD9CM|AB|68.11|Digital exam of uterus
C0177196|ICD9CM|PT|68.15|Closed biopsy of uterine ligaments
C0177196|ICD9CM|AB|68.15|Clos uterine ligament bx
C0177197|ICD9CM|PT|68.16|Closed biopsy of uterus
C0177197|ICD9CM|AB|68.16|Closed uterine biopsy
C0177198|ICD9CM|PT|68.19|Other diagnostic procedures on uterus and supporting structures
C0177198|ICD9CM|AB|68.19|Uterus/adnex dx proc NEC
C0177199|ICD9CM|HT|68.2|Excision or destruction of lesion or tissue of uterus
C0177200|ICD9CM|PT|68.22|Incision or excision of congenital septum of uterus
C0177200|ICD9CM|AB|68.22|Incision uterine septum
C0177201|ICD9CM|PT|68.29|Other excision or destruction of lesion of uterus
C0177201|ICD9CM|AB|68.29|Uterine les destruct NEC
C0177204|ICD9CM|PT|69.02|Dilation and curettage following delivery or abortion
C0177204|ICD9CM|AB|69.02|D & C post delivery
C0177205|ICD9CM|HT|69.1|Excision or destruction of lesion or tissue of uterus and supporting structures
C0177206|ICD9CM|PT|69.19|Other excision or destruction of uterus and supporting structures
C0177206|ICD9CM|AB|69.19|Destruc uter support NEC
C0177207|ICD9CM|HT|69.2|Repair of uterine supporting structures
C0177209|ICD9CM|PT|69.22|Other uterine suspension
C0177209|ICD9CM|AB|69.22|Uterine suspension NEC
C0177210|ICD9CM|PT|69.23|Vaginal repair of chronic inversion of uterus
C0177210|ICD9CM|AB|69.23|Vag repair invers uterus
C0177211|ICD9CM|PT|69.29|Other repair of uterus and supporting structures
C0177211|ICD9CM|AB|69.29|Uterus/adnexa repair NEC
C0177213|ICD9CM|PT|69.49|Other repair of uterus
C0177213|ICD9CM|AB|69.49|Uterine repair NEC
C0177214|ICD9CM|HT|69.5|Aspiration curettage of uterus
C0177215|ICD9CM|PT|69.52|Aspiration curettage following delivery or abortion
C0177215|ICD9CM|AB|69.52|Aspirat curet-post deliv
C0177216|ICD9CM|PT|69.59|Other aspiration curettage of uterus
C0177216|ICD9CM|AB|69.59|Aspir curett uterus NEC
C0177218|ICD9CM|HT|69.9|Other operations on uterus, cervix, and supporting structures
C0177219|ICD9CM|AB|69.93|Insertion of laminaria
C0177219|ICD9CM|PT|69.93|Insertion of laminaria
C0177220|ICD9CM|PT|69.94|Manual replacement of inverted uterus
C0177220|ICD9CM|AB|69.94|Man replace invert uter
C0177221|ICD9CM|PT|69.97|Removal of other penetrating foreign body from cervix
C0177221|ICD9CM|AB|69.97|Remove penetrat cerv FB
C0177222|ICD9CM|PT|69.98|Other operations on supporting structures of uterus
C0177222|ICD9CM|AB|69.98|Uterine support op NEC
C0177223|ICD9CM|PT|69.99|Other operations on cervix and uterus
C0177223|ICD9CM|AB|69.99|Uterine operation NEC
C0177224|ICD9CM|HT|70.1|Incision of vagina and cul-de-sac
C0177225|ICD9CM|PT|70.13|Lysis of intraluminal adhesions of vagina
C0177225|ICD9CM|AB|70.13|Intralum vag adhesiolys
C0177226|ICD9CM|PT|70.14|Other vaginotomy
C0177226|ICD9CM|AB|70.14|Vaginotomy NEC
C0177227|ICD9CM|HT|70.2|Diagnostic procedures on vagina and cul-de-sac
C0177228|ICD9CM|PT|70.29|Other diagnostic procedures on vagina and cul-de-sac
C0177228|ICD9CM|AB|70.29|Vagin/cul-de-sac dx NEC
C0177229|ICD9CM|HT|70.3|Local excision or destruction of vagina and cul-de-sac
C0177230|ICD9CM|PT|70.32|Excision or destruction of lesion of cul-de-sac
C0177230|ICD9CM|AB|70.32|Excis cul-de-sac lesion
C0177232|ICD9CM|HT|70.6|Vaginal construction and reconstruction
C0177234|ICD9CM|PT|70.74|Repair of other vaginoenteric fistula
C0177234|ICD9CM|AB|70.74|Rep vaginoent fistul NEC
C0177235|ICD9CM|PT|70.75|Repair of other fistula of vagina
C0177235|ICD9CM|AB|70.75|Repair vag fistula NEC
C0177236|ICD9CM|HT|70.9|Other operations on vagina and cul-de-sac
C0177237|ICD9CM|PT|70.91|Other operations on vagina
C0177237|ICD9CM|AB|70.91|Vaginal operation NEC
C0177238|ICD9CM|PT|70.92|Other operations on cul-de-sac
C0177238|ICD9CM|AB|70.92|Cul-de-sac operation NEC
C0177239|ICD9CM|HT|71.0|Incision of vulva and perineum
C0177241|ICD9CM|PT|71.09|Other incision of vulva and perineum
C0177241|ICD9CM|AB|71.09|Incis vulva/perineum NEC
C0177242|ICD9CM|HT|71.1|Diagnostic procedures on vulva
C0177243|ICD9CM|PT|71.19|Other diagnostic procedures on vulva
C0177243|ICD9CM|AB|71.19|Vulvar diagnos proc NEC
C0177245|ICD9CM|PT|71.21|Percutaneous aspiration of Bartholin's gland (cyst)
C0177245|ICD9CM|AB|71.21|Percutan bartholin aspir
C0177246|ICD9CM|PT|71.22|Incision of Bartholin's gland (cyst)
C0177246|ICD9CM|AB|71.22|Incise bartholin's gland
C0177248|ICD9CM|PT|71.24|Excision or other destruction of Bartholin's gland (cyst)
C0177248|ICD9CM|AB|71.24|Destruc bartholin gland
C0177249|ICD9CM|PT|71.29|Other operations on Bartholin's gland
C0177249|ICD9CM|AB|71.29|Bartholin's gland op NEC
C0177250|ICD9CM|PT|71.3|Other local excision or destruction of vulva and perineum
C0177250|ICD9CM|AB|71.3|Local vulvar excis NEC
C0177252|ICD9CM|AB|71.5|Radical vulvectomy
C0177252|ICD9CM|PT|71.5|Radical vulvectomy
C0177253|ICD9CM|HT|71.6|Other vulvectomy
C0177254|ICD9CM|HT|71.7|Repair of vulva and perineum
C0177255|ICD9CM|PT|71.71|Suture of laceration of vulva or perineum
C0177255|ICD9CM|AB|71.71|Suture vulvar laceration
C0177256|ICD9CM|PT|71.72|Repair of fistula of vulva or perineum
C0177256|ICD9CM|AB|71.72|Repair vulvar fistula
C0177257|ICD9CM|PT|71.79|Other repair of vulva and perineum
C0177257|ICD9CM|AB|71.79|Vulvar/perin repair NEC
C0177258|ICD9CM|PT|71.8|Other operations on vulva
C0177258|ICD9CM|AB|71.8|Other vulvar operations
C0177260|ICD9CM|PT|72.1|Low forceps operation with episiotomy
C0177260|ICD9CM|AB|72.1|Low forceps w episiotomy
C0177261|ICD9CM|PT|72.21|Mid forceps operation with episiotomy
C0177261|ICD9CM|AB|72.21|Mid forceps w episiotomy
C0177262|ICD9CM|PT|72.29|Other mid forceps operation
C0177262|ICD9CM|AB|72.29|Mid forceps op NEC
C0177263|ICD9CM|PT|72.31|High forceps operation with episiotomy
C0177263|ICD9CM|AB|72.31|High forceps w episiot
C0177264|ICD9CM|PT|72.39|Other high forceps operation
C0177264|ICD9CM|AB|72.39|High forceps op NEC
C0177265|ICD9CM|PT|72.4|Forceps rotation of fetal head
C0177265|ICD9CM|AB|72.4|Forceps rotat fetal head
C0177267|ICD9CM|PT|72.52|Other partial breech extraction
C0177267|ICD9CM|AB|72.52|Part breech extract NEC
C0177269|ICD9CM|PT|72.54|Other total breech extraction
C0177269|ICD9CM|AB|72.54|Tot breech extrac NEC
C0177270|ICD9CM|PT|72.71|Vacuum extraction with episiotomy
C0177270|ICD9CM|AB|72.71|Vacuum ext del w episiot
C0177271|ICD9CM|PT|72.8|Other specified instrumental delivery
C0177271|ICD9CM|AB|72.8|Instrument delivery NEC
C0177274|ICD9CM|PT|73.09|Other artificial rupture of membranes
C0177274|ICD9CM|AB|73.09|Artif rupt membranes NEC
C0177275|ICD9CM|PT|73.1|Other surgical induction of labor
C0177275|ICD9CM|AB|73.1|Surg induct labor NEC
C0177276|ICD9CM|HT|73.5|Manually assisted delivery
C0177277|ICD9CM|PT|73.59|Other manually assisted delivery
C0177277|ICD9CM|AB|73.59|Manual assist deliv NEC
C0177279|ICD9CM|HT|73.9|Other operations assisting delivery
C0177279|ICD9CM|PT|73.99|Other operations assisting delivery
C0177279|ICD9CM|AB|73.99|Ops assisting deliv NEC
C0177283|ICD9CM|HT|75.3|Other intrauterine operations on fetus and amnion
C0177284|ICD9CM|AB|75.32|Fetal ekg
C0177284|ICD9CM|PT|75.32|Fetal EKG (scalp)
C0177285|ICD9CM|PT|75.33|Fetal blood sampling and biopsy
C0177285|ICD9CM|AB|75.33|Fetal blood sample/bx
C0177286|ICD9CM|PT|75.35|Other diagnostic procedures on fetus and amnion
C0177286|ICD9CM|AB|75.35|Dx proc fetus/amnion NEC
C0177287|ICD9CM|PT|75.36|Correction of fetal defect
C0177287|ICD9CM|AB|75.36|Correction fetal defect
C0177288|ICD9CM|PT|75.51|Repair of current obstetric laceration of cervix
C0177288|ICD9CM|AB|75.51|Repair ob lacerat cervix
C0177290|ICD9CM|PT|75.61|Repair of current obstetric laceration of bladder and urethra
C0177290|ICD9CM|AB|75.61|Repair ob lac blad/ureth
C0177291|ICD9CM|PT|75.8|Obstetric tamponade of uterus or vagina
C0177291|ICD9CM|AB|75.8|Ob tamponade uterus/vag
C0177293|ICD9CM|PT|75.92|Evacuation of other hematoma of vulva or vagina
C0177293|ICD9CM|AB|75.92|Evac ob hemat vulva/vag
C0177294|ICD9CM|PT|75.93|Surgical correction of inverted uterus
C0177294|ICD9CM|AB|75.93|Surg corr invert uterus
C0177296|ICD9CM|PT|76.09|Other incision of facial bone
C0177296|ICD9CM|AB|76.09|Facial bone incision NEC
C0177297|ICD9CM|HT|76.1|Diagnostic procedures on facial bones and joints
C0177298|ICD9CM|PT|76.11|Biopsy of facial bone
C0177298|ICD9CM|AB|76.11|Facial bone biopsy
C0177299|ICD9CM|PT|76.19|Other diagnostic procedures on facial bones and joints
C0177299|ICD9CM|AB|76.19|Facial bone dx proc NEC
C0177300|ICD9CM|PT|76.2|Local excision or destruction of lesion of facial bone
C0177300|ICD9CM|AB|76.2|Destruct facial bone les
C0177301|ICD9CM|PT|76.39|Partial ostectomy of other facial bone
C0177301|ICD9CM|AB|76.39|Part facial ostectom NEC
C0177302|ICD9CM|HT|76.4|Excision and reconstruction of facial bones
C0177303|ICD9CM|PT|76.42|Other total mandibulectomy
C0177303|ICD9CM|AB|76.42|Total mandibulectomy NEC
C0177304|ICD9CM|PT|76.43|Other reconstruction of mandible
C0177304|ICD9CM|AB|76.43|Mandibular reconst NEC
C0177305|ICD9CM|PT|76.44|Total ostectomy of other facial bone with synchronous reconstruction
C0177305|ICD9CM|AB|76.44|Tot face ostect w recons
C0177306|ICD9CM|PT|76.45|Other total ostectomy of other facial bone
C0177306|ICD9CM|AB|76.45|Tot face bone ostect NEC
C0177307|ICD9CM|PT|76.46|Other reconstruction of other facial bone
C0177307|ICD9CM|AB|76.46|Facial bone reconstr NEC
C0177308|ICD9CM|HT|76.6|Other facial bone repair and orthognathic surgery
C0177312|ICD9CM|PT|76.64|Other orthognathic surgery on mandible
C0177312|ICD9CM|AB|76.64|Mand orthognathic op NEC
C0177315|ICD9CM|PT|76.69|Other facial bone repair
C0177315|ICD9CM|AB|76.69|Facial bone repair NEC
C0177318|ICD9CM|PT|76.78|Other closed reduction of facial fracture
C0177318|ICD9CM|AB|76.78|Cl reduct facial fx NEC
C0177319|ICD9CM|PT|76.79|Other open reduction of facial fracture
C0177319|ICD9CM|AB|76.79|Open reduct face fx NEC
C0177320|ICD9CM|PT|76.95|Other manipulation of temporomandibular joint
C0177320|ICD9CM|AB|76.95|Tm manipulation NEC
C0177321|ICD9CM|PT|77.01|Sequestrectomy, scapula, clavicle, and thorax [ribs and sternum]
C0177321|ICD9CM|AB|77.01|Chest cage sequestrec
C0177322|ICD9CM|PT|77.02|Sequestrectomy, humerus
C0177322|ICD9CM|AB|77.02|Humerus sequestrectomy
C0177323|ICD9CM|PT|77.03|Sequestrectomy, radius and ulna
C0177323|ICD9CM|AB|77.03|Radius & ulna sequestrec
C0177324|ICD9CM|PT|77.04|Sequestrectomy, carpals and metacarpals
C0177324|ICD9CM|AB|77.04|Metacarp/carp sequestrec
C0177325|ICD9CM|PT|77.08|Sequestrectomy, tarsals and metatarsals
C0177325|ICD9CM|AB|77.08|Metatar/tar sequestrec
C0177326|ICD9CM|PT|77.09|Sequestrectomy, other bones
C0177326|ICD9CM|AB|77.09|Sequestrectomy NEC
C0177327|ICD9CM|HT|77.1|Other incision of bone without division
C0177328|ICD9CM|PT|77.11|Other incision of bone without division, scapula, clavicle, and thorax [ribs and sternum]
C0177328|ICD9CM|AB|77.11|Other chest cage incis
C0177329|ICD9CM|PT|77.12|Other incision of bone without division, humerus
C0177329|ICD9CM|AB|77.12|Other humerus incision
C0177330|ICD9CM|PT|77.13|Other incision of bone without division, radius and ulna
C0177330|ICD9CM|AB|77.13|Other radius/ulna incis
C0177331|ICD9CM|PT|77.14|Other incision of bone without division, carpals and metacarpals
C0177331|ICD9CM|AB|77.14|Oth metacarp/carp incis
C0177332|ICD9CM|PT|77.15|Other incision of bone without division, femur
C0177332|ICD9CM|AB|77.15|Other femoral incision
C0177333|ICD9CM|PT|77.16|Other incision of bone without division, patella
C0177333|ICD9CM|AB|77.16|Other patellar incision
C0177334|ICD9CM|PT|77.17|Other incision of bone without division, tibia and fibula
C0177334|ICD9CM|AB|77.17|Other tibia/fibula incis
C0177335|ICD9CM|PT|77.18|Other incision of bone without division, tarsals and metatarsals
C0177335|ICD9CM|AB|77.18|Oth metatars/tars incis
C0177336|ICD9CM|PT|77.19|Other incision of bone without division, other bones
C0177336|ICD9CM|AB|77.19|Bone incis w/o div NEC
C0177337|ICD9CM|PT|77.21|Wedge osteotomy, scapula, clavicle, and thorax [ribs and sternum]
C0177337|ICD9CM|AB|77.21|Chest cage wedg osteotom
C0177338|ICD9CM|PT|77.27|Wedge osteotomy, tibia and fibula
C0177338|ICD9CM|AB|77.27|Tibia/fibul wedg osteot
C0177339|ICD9CM|PT|77.29|Wedge osteotomy, other bones
C0177339|ICD9CM|AB|77.29|Wedge osteotomy NEC
C0177340|ICD9CM|PT|77.31|Other division of bone, scapula, clavicle, and thorax [ribs and sternum]
C0177340|ICD9CM|AB|77.31|Chest cage bone div NEC
C0177341|ICD9CM|PT|77.32|Other division of bone, humerus
C0177341|ICD9CM|AB|77.32|Humerus division NEC
C0177342|ICD9CM|PT|77.33|Other division of bone, radius and ulna
C0177342|ICD9CM|AB|77.33|Radius/ulna division NEC
C0177343|ICD9CM|PT|77.34|Other division of bone, carpals and metacarpals
C0177343|ICD9CM|AB|77.34|Metacar/car division NEC
C0177344|ICD9CM|PT|77.35|Other division of bone, femur
C0177344|ICD9CM|AB|77.35|Femoral division NEC
C0177345|ICD9CM|PT|77.36|Other division of bone, patella
C0177345|ICD9CM|AB|77.36|Patellar division NEC
C0177346|ICD9CM|PT|77.37|Other division of bone, tibia and fibula
C0177346|ICD9CM|AB|77.37|Tibia/fibula div NEC
C0177347|ICD9CM|PT|77.38|Other division of bone, tarsals and metatarsals
C0177347|ICD9CM|AB|77.38|Metatar/tar division NEC
C0177348|ICD9CM|PT|77.41|Biopsy of bone, scapula, clavicle, and thorax [ribs and sternum]
C0177348|ICD9CM|AB|77.41|Chest cage bone biopsy
C0177349|ICD9CM|PT|77.44|Biopsy of bone, carpals and metacarpals
C0177349|ICD9CM|AB|77.44|Metacarpal/carpal biopsy
C0177350|ICD9CM|PT|77.47|Biopsy of bone, tibia and fibula
C0177350|ICD9CM|AB|77.47|Tibia & fibula biopsy
C0177351|MTH|PN|NOCODE|Bone biopsy NEC in ICD9CM_2014
C0177351|ICD9CM|AB|77.49|Bone biopsy NEC
C0177351|ICD9CM|PT|77.49|Biopsy of bone, other bones
C0177352|ICD9CM|HT|77.5|Excision and repair of bunion and other toe deformities
C0177354|ICD9CM|PT|77.58|Other excision, fusion and repair of toes
C0177354|ICD9CM|AB|77.58|Oth exc, fus, repair toe
C0177355|ICD9CM|PT|77.59|Other bunionectomy
C0177355|ICD9CM|AB|77.59|Bunionectomy NEC
C0177356|ICD9CM|HT|77.6|Local excision of lesion or tissue of bone
C0177357|ICD9CM|PT|77.61|Local excision of lesion or tissue of bone, scapula, clavicle, and thorax [ribs and sternum]
C0177357|ICD9CM|AB|77.61|Exc chest cage bone les
C0177358|ICD9CM|PT|77.64|Local excision of lesion or tissue of bone, carpals and metacarpals
C0177358|ICD9CM|AB|77.64|Loc exc les metacar/car
C0177359|ICD9CM|PT|77.68|Local excision of lesion or tissue of bone, tarsals and metatarsals
C0177359|ICD9CM|AB|77.68|Loc exc les metatar/tar
C0177360|ICD9CM|PT|77.69|Local excision of lesion or tissue of bone, other bones
C0177360|ICD9CM|AB|77.69|Loc exc bone lesion NEC
C0177361|ICD9CM|PT|77.71|Excision of bone for graft, scapula, clavicle, and thorax [ribs and sternum]
C0177361|ICD9CM|AB|77.71|Ex chest cage bone-gft
C0177362|ICD9CM|PT|77.79|Excision of bone for graft, other bones
C0177362|ICD9CM|AB|77.79|Excise bone for gft NEC
C0177364|ICD9CM|PT|77.81|Other partial ostectomy, scapula, clavicle, and thorax [ribs and sternum]
C0177364|ICD9CM|AB|77.81|Oth chest cage ostectomy
C0177365|ICD9CM|PT|77.82|Other partial ostectomy, humerus
C0177365|ICD9CM|AB|77.82|Partial humerectomy NEC
C0177366|ICD9CM|PT|77.83|Other partial ostectomy, radius and ulna
C0177366|ICD9CM|AB|77.83|Part ostect-radius/ulna
C0177367|ICD9CM|PT|77.84|Other partial ostectomy, carpals and metacarpals
C0177367|ICD9CM|AB|77.84|Part ostect-metacar/car
C0177368|ICD9CM|PT|77.85|Other partial ostectomy, femur
C0177368|ICD9CM|AB|77.85|Part ostectomy-femur
C0177369|ICD9CM|PT|77.86|Other partial ostectomy, patella
C0177369|ICD9CM|AB|77.86|Partial patellectomy
C0177370|ICD9CM|PT|77.87|Other partial ostectomy, tibia and fibula
C0177370|ICD9CM|AB|77.87|Part ostect-tibia/fibula
C0177371|ICD9CM|PT|77.88|Other partial ostectomy, tarsals and metatarsals
C0177371|ICD9CM|AB|77.88|Part ostect-metatar/tar
C0177372|ICD9CM|PT|77.89|Other partial ostectomy, other bones
C0177372|ICD9CM|AB|77.89|Partial ostectomy NEC
C0177373|ICD9CM|PT|77.91|Total ostectomy, scapula, clavicle, and thorax [ribs and sternum]
C0177373|ICD9CM|AB|77.91|Tot chest cage ostectomy
C0177374|ICD9CM|PT|77.99|Total ostectomy, other bones
C0177374|ICD9CM|AB|77.99|Total ostectomy NEC
C0177375|ICD9CM|PT|78.01|Bone graft, scapula, clavicle, and thorax [ribs and sternum]
C0177375|ICD9CM|AB|78.01|Bone graft to chest cage
C0177377|ICD9CM|PT|78.04|Bone graft, carpals and metacarpals
C0177377|ICD9CM|AB|78.04|Bone grft to metacar/car
C0177378|ICD9CM|PT|78.07|Bone graft, tibia and fibula
C0177378|ICD9CM|AB|78.07|Bone graft-tibia/fibula
C0177379|ICD9CM|PT|78.08|Bone graft, tarsals and metatarsals
C0177379|ICD9CM|AB|78.08|Bone graft-metatar/tar
C0177380|ICD9CM|PT|78.09|Bone graft, other bones
C0177380|ICD9CM|AB|78.09|Bone graft NEC
C0177382|ICD9CM|PT|78.11|Application of external fixator device, scapula, clavicle, and thorax [ribs and sternum]
C0177382|ICD9CM|AB|78.11|Appl ext fix-chest cage
C0177383|ICD9CM|PT|78.12|Application of external fixator device, humerus
C0177383|ICD9CM|AB|78.12|Applic ext fix-humerus
C0177384|ICD9CM|PT|78.13|Application of external fixator device, radius and ulna
C0177384|ICD9CM|AB|78.13|Appl ext fix-radius/ulna
C0177385|ICD9CM|PT|78.14|Application of external fixator device, carpals and metacarpals
C0177385|ICD9CM|AB|78.14|Appl ext fix-metacar/car
C0177386|ICD9CM|PT|78.15|Application of external fixator device, femur
C0177386|ICD9CM|AB|78.15|Applic ext fix dev-femur
C0177387|ICD9CM|PT|78.16|Application of external fixator device, patella
C0177387|ICD9CM|AB|78.16|Appl ext fix dev-patella
C0177388|ICD9CM|PT|78.17|Application of external fixator device, tibia and fibula
C0177388|ICD9CM|AB|78.17|Appl ext fix-tib/fibula
C0177389|ICD9CM|PT|78.18|Application of external fixator device, tarsals and metatarsals
C0177389|ICD9CM|AB|78.18|Appl ext fix-metatar/tar
C0177390|ICD9CM|PT|78.19|Application of external fixator device, other bones
C0177390|ICD9CM|AB|78.19|Applic ext fix dev NEC
C0177391|ICD9CM|HT|78.2|Limb shortening procedures
C0177392|ICD9CM|PT|78.22|Limb shortening procedures, humerus
C0177392|ICD9CM|AB|78.22|Limb short proc-humerus
C0177393|ICD9CM|PT|78.23|Limb shortening procedures, radius and ulna
C0177393|ICD9CM|AB|78.23|Limb shorten-radius/ulna
C0177394|ICD9CM|PT|78.24|Limb shortening procedures, carpals and metacarpals
C0177394|ICD9CM|AB|78.24|Limb shorten-metacar/car
C0177395|ICD9CM|PT|78.25|Limb shortening procedures, femur
C0177395|ICD9CM|AB|78.25|Limb short proc-femur
C0177396|ICD9CM|PT|78.27|Limb shortening procedures, tibia and fibula
C0177396|ICD9CM|AB|78.27|Limb shorten-tib/fibula
C0177397|ICD9CM|PT|78.28|Limb shortening procedures, tarsals and metatarsals
C0177397|ICD9CM|AB|78.28|Limb shorten-metatar/tar
C0177398|ICD9CM|PT|78.29|Limb shortening procedures, other bones
C0177398|ICD9CM|AB|78.29|Limb shorten proc NEC
C0177400|ICD9CM|PT|78.32|Limb lengthening procedures, humerus
C0177400|ICD9CM|AB|78.32|Limb length proc-humerus
C0177401|ICD9CM|PT|78.33|Limb lengthening procedures, radius and ulna
C0177401|ICD9CM|AB|78.33|Limb length-radius/ulna
C0177402|ICD9CM|PT|78.34|Limb lengthening procedures, carpals and metacarpals
C0177402|ICD9CM|AB|78.34|Limb length-metacar/car
C0177403|ICD9CM|PT|78.35|Limb lengthening procedures, femur
C0177403|ICD9CM|AB|78.35|Limb length proc-femur
C0177404|ICD9CM|PT|78.37|Limb lengthening procedures, tibia and fibula
C0177404|ICD9CM|AB|78.37|Limb lengthen-tib/fibula
C0177405|ICD9CM|PT|78.38|Limb lengthening procedures, tarsals and metatarsals
C0177405|ICD9CM|AB|78.38|Limb lengthn-metatar/tar
C0177406|ICD9CM|PT|78.39|Limb lengthening procedures, other bones
C0177406|ICD9CM|AB|78.39|Limb lengthen proc NEC
C0177408|ICD9CM|PT|78.41|Other repair or plastic operations on bone, scapula, clavicle, and thorax [ribs and sternum]
C0177408|ICD9CM|AB|78.41|Oth chest cage rep/plast
C0177409|ICD9CM|PT|78.42|Other repair or plastic operations on bone, humerus
C0177409|ICD9CM|AB|78.42|Oth humerus repair/plast
C0177410|ICD9CM|PT|78.43|Other repair or plastic operations on bone, radius and ulna
C0177410|ICD9CM|AB|78.43|Oth rad/uln repair/plast
C0177411|ICD9CM|PT|78.44|Other repair or plastic operations on bone, carpals and metacarpals
C0177411|ICD9CM|AB|78.44|Oth metac/carp rep/plast
C0177412|ICD9CM|PT|78.45|Other repair or plastic operations on bone, femur
C0177412|ICD9CM|AB|78.45|Oth femur repair/plastic
C0177413|ICD9CM|PT|78.46|Other repair or plastic operations on bone, patella
C0177413|ICD9CM|AB|78.46|Oth patella repair/plast
C0177414|ICD9CM|PT|78.47|Other repair or plastic operations on bone, tibia and fibula
C0177414|ICD9CM|AB|78.47|Oth tib/fib repair/plast
C0177415|ICD9CM|PT|78.48|Other repair or plastic operations on bone, tarsals and metatarsals
C0177415|ICD9CM|AB|78.48|Oth meta/tar repa/plast
C0177416|ICD9CM|PT|78.49|Other repair or plastic operations on bone, other bones
C0177416|ICD9CM|AB|78.49|Oth bone repa/plast NEC
C0177417|ICD9CM|PT|78.51|Internal fixation of bone without fracture reduction, scapula, clavicle, and thorax [ribs and sternum]
C0177417|ICD9CM|AB|78.51|Int fixation-chest cage
C0177418|ICD9CM|PT|78.59|Internal fixation of bone without fracture reduction, other bones
C0177418|ICD9CM|AB|78.59|Int fix-no fx reduct NEC
C0177421|ICD9CM|PT|78.61|Removal of implanted devices from bone, scapula, clavicle, and thorax [ribs and sternum]
C0177421|ICD9CM|AB|78.61|Remov imp dev-chest cage
C0177422|ICD9CM|PT|78.62|Removal of implanted devices from bone, humerus
C0177422|ICD9CM|AB|78.62|Remove impl dev-humerus
C0177423|ICD9CM|PT|78.63|Removal of implanted devices from bone, radius and ulna
C0177423|ICD9CM|AB|78.63|Remov imp dev-radius/uln
C0177424|ICD9CM|PT|78.64|Removal of implanted devices from bone, carpals and metacarpals
C0177424|ICD9CM|AB|78.64|Remov imp dev-metac/carp
C0177425|ICD9CM|PT|78.65|Removal of implanted devices from bone, femur
C0177425|ICD9CM|AB|78.65|Remove imp device-femur
C0177426|ICD9CM|PT|78.66|Removal of implanted devices from bone, patella
C0177426|ICD9CM|AB|78.66|Remov imp device-patella
C0177427|ICD9CM|PT|78.67|Removal of implanted devices from bone, tibia and fibula
C0177427|ICD9CM|AB|78.67|Remov imp dev-tib/fibula
C0177428|ICD9CM|PT|78.68|Removal of implanted devices from bone, tarsals and metatarsals
C0177428|ICD9CM|AB|78.68|Remove imp dev-metat/tar
C0177429|ICD9CM|PT|78.69|Removal of implanted devices from bone, other bones
C0177429|ICD9CM|AB|78.69|Remove impl device NEC
C0177430|ICD9CM|PT|78.71|Osteoclasis, scapula, clavicle, and thorax [ribs and sternum]
C0177430|ICD9CM|AB|78.71|Osteoclasis-chest cage
C0177431|ICD9CM|PT|78.73|Osteoclasis, radius and ulna
C0177431|ICD9CM|AB|78.73|Osteoclasis-radius/ulna
C0177432|ICD9CM|PT|78.74|Osteoclasis, carpals and metacarpals
C0177432|ICD9CM|AB|78.74|Osteoclasis-metacar/car
C0177433|ICD9CM|PT|78.78|Osteoclasis, tarsals and metatarsals
C0177433|ICD9CM|AB|78.78|Osteoclasis-metatar/tar
C0177434|ICD9CM|PT|78.79|Osteoclasis, other bones
C0177434|ICD9CM|AB|78.79|Osteoclasis NEC
C0177446|ICD9CM|PT|78.91|Insertion of bone growth stimulator, scapula, clavicle and thorax [ribs and sternum]
C0177446|ICD9CM|AB|78.91|Insert bone stimul-chest
C0177447|ICD9CM|PT|78.99|Insertion of bone growth stimulator, other bones
C0177447|ICD9CM|AB|78.99|Insert bone stimul NEC
C0177457|ICD9CM|PT|79.22|Open reduction of fracture without internal fixation, radius and ulna
C0177457|ICD9CM|AB|79.22|Open reduc-radius/uln fx
C0177458|ICD9CM|PT|79.23|Open reduction of fracture without internal fixation, carpals and metacarpals
C0177458|ICD9CM|AB|79.23|Open reduc-metac/car fx
C0177459|ICD9CM|PT|79.24|Open reduction of fracture without internal fixation, phalanges of hand
C0177459|ICD9CM|AB|79.24|Open reduction-finger fx
C0177460|ICD9CM|PT|79.25|Open reduction of fracture without internal fixation, femur
C0177460|ICD9CM|AB|79.25|Open reduction-femur fx
C0177461|ICD9CM|PT|79.26|Open reduction of fracture without internal fixation, tibia and fibula
C0177461|ICD9CM|AB|79.26|Open reduc-tibia/fib fx
C0177462|ICD9CM|PT|79.27|Open reduction of fracture without internal fixation, tarsals and metatarsals
C0177462|ICD9CM|AB|79.27|Open reduc-metat/tars fx
C0177463|ICD9CM|PT|79.28|Open reduction of fracture without internal fixation, phalanges of foot
C0177463|ICD9CM|AB|79.28|Open reduction-toe fx
C0177464|ICD9CM|PT|79.29|Open reduction of fracture without internal fixation, other specified bone
C0177464|ICD9CM|AB|79.29|Open fx reduction NEC
C0177465|ICD9CM|PT|79.39|Open reduction of fracture with internal fixation, other specified bone
C0177465|ICD9CM|AB|79.39|Opn fx red w int fix NEC
C0177466|ICD9CM|PT|79.49|Closed reduction of separated epiphysis, other specified bone
C0177466|ICD9CM|AB|79.49|Cls reduc-sep epiphy NEC
C0177468|ICD9CM|PT|79.59|Open reduction of separated epiphysis, other specified bone
C0177468|ICD9CM|AB|79.59|Open red-sep epiphy NEC
C0177469|ICD9CM|HT|79.6|Debridement of open fracture site
C0177469|ICD9CM|PT|79.60|Debridement of open fracture, unspecified site
C0177469|ICD9CM|AB|79.60|Open fx site debride NOS
C0177470|ICD9CM|PT|79.63|Debridement of open fracture site, carpals and metacarpals
C0177470|ICD9CM|AB|79.63|Debrid opn fx-metac/car
C0177472|ICD9CM|PT|79.69|Debridement of open fracture site, other specified bone
C0177472|ICD9CM|AB|79.69|Open fx site debride NEC
C0177473|ICD9CM|PT|79.70|Closed reduction of dislocation of unspecified site
C0177473|ICD9CM|AB|79.70|Cl reduc disloc NOS
C0177474|ICD9CM|PT|79.74|Closed reduction of dislocation of hand and finger
C0177474|ICD9CM|AB|79.74|Cl reduc disloc-hand/fng
C0177475|ICD9CM|PT|79.75|Closed reduction of dislocation of hip
C0177475|ICD9CM|AB|79.75|Cl reduc disloc-hip
C0177476|ICD9CM|PT|79.79|Closed reduction of dislocation of other specified sites
C0177476|ICD9CM|AB|79.79|Cl reduc dislocation NEC
C0177477|ICD9CM|PT|79.80|Open reduction of dislocation of unspecified site
C0177477|ICD9CM|AB|79.80|Open reduc-dislocat NOS
C0177478|ICD9CM|PT|79.84|Open reduction of dislocation of hand and finger
C0177478|ICD9CM|AB|79.84|Opn reduc disloc-hand
C0177479|ICD9CM|PT|79.89|Open reduction of dislocation of other specified sites
C0177479|ICD9CM|AB|79.89|Open reduc-dislocat NEC
C0177482|ICD9CM|PT|79.92|Unspecified operation on bone injury, radius and ulna
C0177482|ICD9CM|AB|79.92|Radius/ulna inj op NOS
C0177489|ICD9CM|PT|79.99|Unspecified operation on bone injury, other specified bone
C0177489|ICD9CM|AB|79.99|Unspec op-bone inj NEC
C0177493|ICD9CM|HT|80.1|Other arthrotomy
C0177494|ICD9CM|PT|80.11|Other arthrotomy, shoulder
C0177494|ICD9CM|AB|80.11|Oth arthrotomy-shoulder
C0177495|ICD9CM|PT|80.12|Other arthrotomy, elbow
C0177495|ICD9CM|AB|80.12|Oth arthrotomy-elbow
C0177496|ICD9CM|PT|80.13|Other arthrotomy, wrist
C0177496|ICD9CM|AB|80.13|Oth arthrotomy-wrist
C0177497|ICD9CM|PT|80.14|Other arthrotomy, hand and finger
C0177497|ICD9CM|AB|80.14|Oth arthrotomy-hand/fngr
C0177498|ICD9CM|PT|80.15|Other arthrotomy, hip
C0177498|ICD9CM|AB|80.15|Oth arthrotomy-hip
C0177499|ICD9CM|PT|80.16|Other arthrotomy, knee
C0177499|ICD9CM|AB|80.16|Oth arthrotomy-knee
C0177500|ICD9CM|PT|80.17|Other arthrotomy, ankle
C0177500|ICD9CM|AB|80.17|Oth arthrotomy-ankle
C0177501|ICD9CM|PT|80.18|Other arthrotomy, foot and toe
C0177501|ICD9CM|AB|80.18|Oth arthrotomy-foot/toe
C0177502|ICD9CM|PT|80.19|Other arthrotomy, other specified sites
C0177502|ICD9CM|AB|80.19|Other arthrotomy NEC
C0177503|ICD9CM|PT|80.24|Arthroscopy, hand and finger
C0177503|ICD9CM|AB|80.24|Hand & finger arthroscop
C0177504|ICD9CM|PT|80.28|Arthroscopy, foot and toe
C0177504|ICD9CM|AB|80.28|Foot & toe arthroscopy
C0177505|ICD9CM|AB|80.35|Hip joint biopsy
C0177505|ICD9CM|PT|80.35|Biopsy of joint structure, hip
C0177506|ICD9CM|PT|80.39|Biopsy of joint structure, other specified sites
C0177506|ICD9CM|AB|80.39|Joint biopsy NEC
C0177507|ICD9CM|HT|80.4|Division of joint capsule, ligament, or cartilage
C0177508|ICD9CM|PT|80.41|Division of joint capsule, ligament, or cartilage, shoulder
C0177508|ICD9CM|AB|80.41|Shoulder struct division
C0177509|ICD9CM|PT|80.42|Division of joint capsule, ligament, or cartilage, elbow
C0177509|ICD9CM|AB|80.42|Elbow structure division
C0177510|ICD9CM|PT|80.43|Division of joint capsule, ligament, or cartilage, wrist
C0177510|ICD9CM|AB|80.43|Wrist structure division
C0177511|ICD9CM|PT|80.44|Division of joint capsule, ligament, or cartilage, hand and finger
C0177511|ICD9CM|AB|80.44|Hand joint struct divis
C0177512|ICD9CM|PT|80.45|Division of joint capsule, ligament, or cartilage, hip
C0177512|ICD9CM|AB|80.45|Hip structure division
C0177513|ICD9CM|PT|80.46|Division of joint capsule, ligament, or cartilage, knee
C0177513|ICD9CM|AB|80.46|Knee structure division
C0177514|ICD9CM|PT|80.47|Division of joint capsule, ligament, or cartilage, ankle
C0177514|ICD9CM|AB|80.47|Ankle structure division
C0177515|ICD9CM|PT|80.48|Division of joint capsule, ligament, or cartilage, foot and toe
C0177515|ICD9CM|AB|80.48|Foot joint struct divis
C0177516|ICD9CM|PT|80.49|Division of joint capsule, ligament, or cartilage, other specified sites
C0177516|ICD9CM|AB|80.49|Jt structur division NEC
C0177518|ICD9CM|PT|80.59|Other destruction of intervertebral disc
C0177518|ICD9CM|AB|80.59|Oth exc/dest intvrt disc
C0177519|ICD9CM|PT|80.74|Synovectomy, hand and finger
C0177519|ICD9CM|AB|80.74|Hand synovectomy
C0177520|ICD9CM|PT|80.79|Synovectomy, other specified sites
C0177520|ICD9CM|AB|80.79|Synovectomy-site NEC
C0177521|ICD9CM|HT|80.8|Other local excision or destruction of lesion of joint
C0177522|ICD9CM|PT|80.81|Other local excision or destruction of lesion of joint, shoulder
C0177522|ICD9CM|AB|80.81|Destruc-shoulder les NEC
C0177523|ICD9CM|PT|80.82|Other local excision or destruction of lesion of joint, elbow
C0177523|ICD9CM|AB|80.82|Destruc-elbow lesion NEC
C0177524|ICD9CM|PT|80.83|Other local excision or destruction of lesion of joint, wrist
C0177524|ICD9CM|AB|80.83|Destruc-wrist lesion NEC
C0177525|ICD9CM|PT|80.84|Other local excision or destruction of lesion of joint, hand and finger
C0177525|ICD9CM|AB|80.84|Destruc-hand jt les NEC
C0177526|ICD9CM|PT|80.85|Other local excision or destruction of lesion of joint, hip
C0177526|ICD9CM|AB|80.85|Destruct-hip lesion NEC
C0177527|ICD9CM|PT|80.86|Other local excision or destruction of lesion of joint, knee
C0177527|ICD9CM|AB|80.86|Destruct-knee lesion NEC
C0177528|ICD9CM|PT|80.87|Other local excision or destruction of lesion of joint, ankle
C0177528|ICD9CM|AB|80.87|Destruc-ankle lesion NEC
C0177529|ICD9CM|PT|80.88|Other local excision or destruction of lesion of joint, foot and toe
C0177529|ICD9CM|AB|80.88|Destruc-foot jt les NEC
C0177530|ICD9CM|PT|80.89|Other local excision or destruction of lesion of joint, other specified sites
C0177530|ICD9CM|AB|80.89|Destruct joint les NEC
C0177531|ICD9CM|HT|80.9|Other excision of joint
C0177532|ICD9CM|PT|80.91|Other excision of joint, shoulder
C0177532|ICD9CM|AB|80.91|Excision of shoulder NEC
C0177533|ICD9CM|PT|80.92|Other excision of joint, elbow
C0177533|ICD9CM|AB|80.92|Excision of elbow NEC
C0177534|ICD9CM|PT|80.93|Other excision of joint, wrist
C0177534|ICD9CM|AB|80.93|Excision of wrist NEC
C0177535|ICD9CM|PT|80.94|Other excision of joint, hand and finger
C0177535|ICD9CM|AB|80.94|Excision hand joint NEC
C0177536|ICD9CM|PT|80.95|Other excision of joint, hip
C0177536|ICD9CM|AB|80.95|Excision of hip NEC
C0177537|ICD9CM|PT|80.96|Other excision of joint, knee
C0177537|ICD9CM|AB|80.96|Excision of knee NEC
C0177538|ICD9CM|PT|80.97|Other excision of joint, ankle
C0177538|ICD9CM|AB|80.97|Excision of ankle NEC
C0177539|ICD9CM|PT|80.98|Other excision of joint, foot and toe
C0177539|ICD9CM|AB|80.98|Excision foot joint NEC
C0177540|MTH|PN|NOCODE|Excision of joint NEC in ICD9CM_2014
C0177540|ICD9CM|PT|80.99|Other excision of joint, other specified sites
C0177540|ICD9CM|AB|80.99|Excision of joint NEC
C0177542|ICD9CM|PT|81.02|Other cervical fusion of the anterior column, anterior technique
C0177542|ICD9CM|AB|81.02|Oth cerv fusion ant/ant
C0177543|ICD9CM|PT|81.03|Other cervical fusion of the posterior column, posterior technique
C0177543|ICD9CM|AB|81.03|Ot cerv fusion post/post
C0177553|ICD9CM|AB|81.17|Other fusion of foot
C0177553|ICD9CM|PT|81.17|Other fusion of foot
C0177554|ICD9CM|HT|81.2|Arthrodesis of other joint
C0177557|ICD9CM|HT|81.4|Other repair of joint of lower extremity
C0177558|ICD9CM|AB|81.44|Patellar stabilization
C0177558|ICD9CM|PT|81.44|Patellar stabilization
C0177559|ICD9CM|PT|81.45|Other repair of the cruciate ligaments
C0177559|ICD9CM|AB|81.45|Cruciate lig repair NEC
C0177560|ICD9CM|PT|81.46|Other repair of the collateral ligaments
C0177560|ICD9CM|AB|81.46|Collaterl lig repair NEC
C0177561|ICD9CM|AB|81.47|Other repair of knee
C0177561|ICD9CM|PT|81.47|Other repair of knee
C0177562|ICD9CM|AB|81.49|Other repair of ankle
C0177562|ICD9CM|PT|81.49|Other repair of ankle
C0177563|ICD9CM|HT|81.5|Joint replacement of lower extremity
C0177565|ICD9CM|HT|81.7|Arthroplasty and repair of hand, fingers, and wrist
C0177566|ICD9CM|PT|81.72|Arthroplasty of metacarpophalangeal and interphalangeal joint without implant
C0177566|ICD9CM|AB|81.72|Arthroplasty metacar w/o
C0177567|ICD9CM|PT|81.74|Arthroplasty of carpocarpal or carpometacarpal joint with implant
C0177567|ICD9CM|AB|81.74|Arthroplasty carpal wit
C0177568|ICD9CM|PT|81.75|Arthroplasty of carpocarpal or carpometacarpal joint without implant
C0177568|ICD9CM|AB|81.75|Arthroplasty carpal w/o
C0177569|ICD9CM|PT|81.79|Other repair of hand, fingers, and wrist
C0177569|ICD9CM|AB|81.79|Oth repair han/fin/wris
C0177570|ICD9CM|HT|81.8|Arthroplasty and repair of shoulder and elbow
C0177571|ICD9CM|PT|81.83|Other repair of shoulder
C0177571|ICD9CM|AB|81.83|Shoulder arthroplast NEC
C0177572|ICD9CM|PT|81.85|Other repair of elbow
C0177572|ICD9CM|AB|81.85|Elbow arthroplasty NEC
C0177573|ICD9CM|PT|81.92|Injection of therapeutic substance into joint or ligament
C0177573|ICD9CM|AB|81.92|Injection into joint
C0177574|ICD9CM|PT|81.93|Suture of capsule or ligament of upper extremity
C0177574|ICD9CM|AB|81.93|Sutur capsul/ligamen arm
C0177575|ICD9CM|PT|81.94|Suture of capsule or ligament of ankle and foot
C0177575|ICD9CM|AB|81.94|Suture capsul/lig ank/ft
C0177576|ICD9CM|PT|81.95|Suture of capsule or ligament of other lower extremity
C0177576|ICD9CM|AB|81.95|Sutur capsul/lig leg NEC
C0177577|ICD9CM|PT|81.98|Other diagnostic procedures on joint structures
C0177577|ICD9CM|AB|81.98|Other joint dx procedure
C0177578|ICD9CM|HT|82.0|Incision of muscle, tendon, fascia, and bursa of hand
C0177579|ICD9CM|PT|82.04|Incision and drainage of palmar or thenar space
C0177579|ICD9CM|AB|82.04|I & d palmar/thenar spac
C0177580|ICD9CM|PT|82.09|Other incision of soft tissue of hand
C0177580|ICD9CM|AB|82.09|Inc soft tissue hand NEC
C0177581|ICD9CM|HT|82.1|Division of muscle, tendon, and fascia of hand
C0177582|ICD9CM|PT|82.19|Other division of soft tissue of hand
C0177582|ICD9CM|AB|82.19|Div soft tissue hand NEC
C0177583|ICD9CM|HT|82.2|Excision of lesion of muscle, tendon, and fascia of hand
C0177584|ICD9CM|PT|82.29|Excision of other lesion of soft tissue of hand
C0177584|ICD9CM|AB|82.29|Exc les sft tiss hnd NEC
C0177585|ICD9CM|PT|82.33|Other tenonectomy of hand
C0177585|ICD9CM|AB|82.33|Hand tenonectomy NEC
C0177586|ICD9CM|PT|82.34|Excision of muscle or fascia of hand for graft
C0177586|ICD9CM|AB|82.34|Exc hnd mus/fas for grft
C0177587|ICD9CM|PT|82.35|Other fasciectomy of hand
C0177587|ICD9CM|AB|82.35|Hand fasciectomy NEC
C0177588|ICD9CM|AB|82.36|Other myectomy of hand
C0177588|ICD9CM|PT|82.36|Other myectomy of hand
C0177589|ICD9CM|HT|82.4|Suture of muscle, tendon, and fascia of hand
C0177591|ICD9CM|PT|82.43|Delayed suture of other tendon of hand
C0177591|ICD9CM|AB|82.43|Delay sut hand tend NEC
C0177592|ICD9CM|PT|82.44|Other suture of flexor tendon of hand
C0177592|ICD9CM|AB|82.44|Sutur flex tend hand NEC
C0177593|ICD9CM|PT|82.45|Other suture of other tendon of hand
C0177593|ICD9CM|AB|82.45|Suture hand tendon NEC
C0177594|ICD9CM|PT|82.46|Suture of muscle or fascia of hand
C0177594|ICD9CM|AB|82.46|Suture hand muscle/fasc
C0177595|ICD9CM|HT|82.5|Transplantation of muscle and tendon of hand
C0177596|ICD9CM|PT|82.55|Other change in hand muscle or tendon length
C0177596|ICD9CM|AB|82.55|Chng hnd mus/ten lng NEC
C0177597|ICD9CM|PT|82.56|Other hand tendon transfer or transplantation
C0177597|ICD9CM|AB|82.56|Transplant hand tend NEC
C0177598|ICD9CM|PT|82.57|Other hand tendon transposition
C0177598|ICD9CM|AB|82.57|Transposit hand tend NEC
C0177599|ICD9CM|PT|82.58|Other hand muscle transfer or transplantation
C0177599|ICD9CM|AB|82.58|Transplant hand musc NEC
C0177600|ICD9CM|PT|82.59|Other hand muscle transposition
C0177600|ICD9CM|AB|82.59|Transposit hand musc NEC
C0177601|ICD9CM|HT|82.6|Reconstruction of thumb
C0177602|ICD9CM|PT|82.61|Pollicization operation carrying over nerves and blood supply
C0177602|ICD9CM|AB|82.61|Pollicization operation
C0177603|ICD9CM|PT|82.69|Other reconstruction of thumb
C0177603|ICD9CM|AB|82.69|Thumb reconstruction NEC
C0177605|ICD9CM|PT|82.72|Plastic operation on hand with graft of muscle or fascia
C0177605|ICD9CM|AB|82.72|Plast op hnd-mus/fas grf
C0177606|ICD9CM|PT|82.79|Plastic operation on hand with other graft or implant
C0177606|ICD9CM|AB|82.79|Plast op hand w grft NEC
C0177608|ICD9CM|AB|82.85|Other tenodesis of hand
C0177608|ICD9CM|PT|82.85|Other tenodesis of hand
C0177609|ICD9CM|AB|82.86|Other tenoplasty of hand
C0177609|ICD9CM|PT|82.86|Other tenoplasty of hand
C0177610|ICD9CM|HT|82.9|Other operations on muscle, tendon, and fascia of hand
C0177610|ICD9CM|PT|82.99|Other operations on muscle, tendon, and fascia of hand
C0177610|ICD9CM|AB|82.99|Hand mus/ten/fas/ops NEC
C0177611|ICD9CM|PT|82.93|Aspiration of other soft tissue of hand
C0177611|ICD9CM|AB|82.93|Aspir soft tiss hand NEC
C0177612|ICD9CM|PT|82.96|Other injection of locally-acting therapeutic substance into soft tissue of hand
C0177612|ICD9CM|AB|82.96|Hand sft tissu injec NEC
C0177613|ICD9CM|HT|83.0|Incision of muscle, tendon, fascia, and bursa
C0177614|ICD9CM|PT|83.09|Other incision of soft tissue
C0177614|ICD9CM|AB|83.09|Soft tissue incision NEC
C0177615|ICD9CM|HT|83.1|Division of muscle, tendon, and fascia
C0177616|ICD9CM|AB|83.13|Other tenotomy
C0177616|ICD9CM|PT|83.13|Other tenotomy
C0177617|ICD9CM|PT|83.19|Other division of soft tissue
C0177617|ICD9CM|AB|83.19|Soft tissue division NEC
C0177618|ICD9CM|HT|83.2|Diagnostic procedures on muscle, tendon, fascia, and bursa, including that of hand
C0177619|ICD9CM|PT|83.29|Other diagnostic procedures on muscle, tendon, fascia, and bursa, including that of hand
C0177619|ICD9CM|AB|83.29|Soft tissue dx proc NEC
C0177620|ICD9CM|HT|83.3|Excision of lesion of muscle, tendon, fascia, and bursa
C0177621|ICD9CM|PT|83.39|Excision of lesion of other soft tissue
C0177621|ICD9CM|AB|83.39|Exc les soft tissue NEC
C0177622|ICD9CM|HT|83.4|Other excision of muscle, tendon, and fascia
C0177623|ICD9CM|AB|83.42|Other tenonectomy
C0177623|ICD9CM|PT|83.42|Other tenonectomy
C0177625|ICD9CM|AB|83.44|Other fasciectomy
C0177625|ICD9CM|PT|83.44|Other fasciectomy
C0177626|ICD9CM|AB|83.45|Other myectomy
C0177626|ICD9CM|PT|83.45|Other myectomy
C0177627|ICD9CM|PT|83.49|Other excision of soft tissue
C0177627|ICD9CM|AB|83.49|Other soft tissue excis
C0177628|ICD9CM|HT|83.6|Suture of muscle, tendon, and fascia
C0177629|ICD9CM|AB|83.64|Other suture of tendon
C0177629|ICD9CM|PT|83.64|Other suture of tendon
C0177630|ICD9CM|PT|83.65|Other suture of muscle or fascia
C0177630|ICD9CM|AB|83.65|Other muscle/fasc suture
C0177631|ICD9CM|HT|83.7|Reconstruction of muscle and tendon
C0177632|ICD9CM|PT|83.76|Other tendon transposition
C0177632|ICD9CM|AB|83.76|Other tendon transposit
C0177633|ICD9CM|PT|83.77|Muscle transfer or transplantation
C0177633|ICD9CM|AB|83.77|Muscle trnsfr/transplant
C0177634|ICD9CM|PT|83.79|Other muscle transposition
C0177634|ICD9CM|AB|83.79|Other muscle transposit
C0177635|ICD9CM|HT|83.8|Other plastic operations on muscle, tendon, and fascia
C0177636|ICD9CM|PT|83.82|Graft of muscle or fascia
C0177636|ICD9CM|AB|83.82|Muscle or fascia graft
C0177637|ICD9CM|PT|83.85|Other change in muscle or tendon length
C0177637|ICD9CM|AB|83.85|Musc/tend lng change NEC
C0177638|ICD9CM|PT|83.87|Other plastic operations on muscle
C0177638|ICD9CM|AB|83.87|Other plastic ops muscle
C0177639|ICD9CM|PT|83.88|Other plastic operations on tendon
C0177639|ICD9CM|AB|83.88|Other plastic ops tendon
C0177640|ICD9CM|PT|83.89|Other plastic operations on fascia
C0177640|ICD9CM|AB|83.89|Other plastic ops fascia
C0177641|ICD9CM|HT|83.9|Other operations on muscle, tendon, fascia, and bursa
C0177641|ICD9CM|PT|83.99|Other operations on muscle, tendon, fascia, and bursa
C0177641|ICD9CM|AB|83.99|Mus/ten/fas/bur op NEC
C0177642|ICD9CM|PT|83.91|Lysis of adhesions of muscle, tendon, fascia, and bursa
C0177642|ICD9CM|AB|83.91|Adhesiolysis mus/ten/fas
C0177643|ICD9CM|PT|83.92|Insertion or replacement of skeletal muscle stimulator
C0177643|ICD9CM|AB|83.92|Insert skel musc stimula
C0177644|ICD9CM|PT|83.95|Aspiration of other soft tissue
C0177644|ICD9CM|AB|83.95|Soft tissue aspirat NEC
C0177645|ICD9CM|PT|83.98|Injection of locally acting therapeutic substance into other soft tissue
C0177645|ICD9CM|AB|83.98|Soft tissue inject NEC
C0177646|ICD9CM|PT|84.01|Amputation and disarticulation of finger
C0177646|ICD9CM|AB|84.01|Finger amputation
C0177649|ICD9CM|PT|84.15|Other amputation below knee
C0177649|ICD9CM|AB|84.15|Below knee amputat NEC
C0177650|ICD9CM|AB|84.21|Thumb reattachment
C0177650|ICD9CM|PT|84.21|Thumb reattachment
C0177652|ICD9CM|PT|84.23|Forearm, wrist, or hand reattachment
C0177652|ICD9CM|AB|84.23|Forearm/wrist/hand reatt
C0177654|ICD9CM|AB|84.25|Toe reattachment
C0177654|ICD9CM|PT|84.25|Toe reattachment
C0177656|ICD9CM|PT|84.27|Lower leg or ankle reattachment
C0177656|ICD9CM|AB|84.27|Lower leg/ankle reattach
C0177657|ICD9CM|AB|84.28|Thigh reattachment
C0177657|ICD9CM|PT|84.28|Thigh reattachment
C0177658|ICD9CM|PT|84.29|Other reattachment of extremity
C0177658|ICD9CM|AB|84.29|Reattachment NEC
C0177660|ICD9CM|PT|84.41|Fitting of prosthesis of upper arm and shoulder
C0177660|ICD9CM|AB|84.41|Fit up arm/should prosth
C0177661|ICD9CM|PT|84.42|Fitting of prosthesis of lower arm and hand
C0177661|ICD9CM|AB|84.42|Fit lo arm/hand prosthes
C0177662|ICD9CM|AB|84.43|Fit arm prosthesis NOS
C0177662|ICD9CM|PT|84.43|Fitting of prosthesis of arm, not otherwise specified
C0177663|ICD9CM|HT|84.9|Other operations on musculoskeletal system
C0177663|ICD9CM|PT|84.99|Other operations on musculoskeletal system
C0177663|ICD9CM|HT|84|Other procedures on musculoskeletal system
C0177663|ICD9CM|AB|84.99|Musculoskeletal op NEC
C0177664|ICD9CM|PT|84.92|Separation of equal conjoined twins
C0177664|ICD9CM|AB|84.92|Separat equal join twin
C0177666|ICD9CM|PT|85.11|Closed [percutaneous] [needle] biopsy of breast
C0177666|ICD9CM|AB|85.11|Closed breast biopsy
C0177667|ICD9CM|PT|85.12|Open biopsy of breast
C0177667|ICD9CM|AB|85.12|Open breast biopsy
C0177668|ICD9CM|PT|85.19|Other diagnostic procedures on breast
C0177668|ICD9CM|AB|85.19|Breast dx procedure NEC
C0177671|ICD9CM|HT|85.3|Reduction mammoplasty and subcutaneous mammectomy
C0177672|ICD9CM|PT|85.36|Other bilateral subcutaneous mammectomy
C0177672|ICD9CM|AB|85.36|Bilat subq mammectom NEC
C0177674|ICD9CM|PT|85.51|Unilateral injection into breast for augmentation
C0177674|ICD9CM|AB|85.51|Unil breast injec-augmen
C0177675|ICD9CM|PT|85.52|Bilateral injection into breast for augmentation
C0177675|ICD9CM|AB|85.52|Bil breast injec-augment
C0177676|ICD9CM|HT|85.7|Total reconstruction of breast
C0177677|ICD9CM|HT|85.8|Other repair and plastic operations on breast
C0177678|ICD9CM|PT|85.87|Other repair or reconstruction of nipple
C0177678|ICD9CM|AB|85.87|Nipple repair NEC
C0177679|ICD9CM|PT|85.89|Other mammoplasty
C0177679|ICD9CM|AB|85.89|Mammoplasty NEC
C0177680|ICD9CM|HT|85.9|Other operations on the breast
C0177680|ICD9CM|PT|85.99|Other operations on the breast
C0177680|ICD9CM|AB|85.99|Breast operation NEC
C0177682|ICD9CM|PT|85.95|Insertion of breast tissue expander
C0177682|ICD9CM|AB|85.95|Inser breast tissu expan
C0177684|ICD9CM|HT|86.0|Incision of skin and subcutaneous tissue
C0177685|ICD9CM|PT|86.01|Aspiration of skin and subcutaneous tissue
C0177685|ICD9CM|AB|86.01|Aspiration skin & subq
C0177686|ICD9CM|PT|86.02|Injection or tattooing of skin lesion or defect
C0177686|ICD9CM|AB|86.02|Skin defect tattooing
C0177687|ICD9CM|PT|86.03|Incision of pilonidal sinus or cyst
C0177687|ICD9CM|AB|86.03|Incision pilonidal sinus
C0177688|ICD9CM|PT|86.04|Other incision with drainage of skin and subcutaneous tissue
C0177688|ICD9CM|AB|86.04|Other skin & subq i & d
C0177690|ICD9CM|PT|86.06|Insertion of totally implantable infusion pump
C0177690|ICD9CM|AB|86.06|Insert infusion pump
C0177691|ICD9CM|PT|86.07|Insertion of totally implantable vascular access device [VAD]
C0177691|ICD9CM|AB|86.07|Insert vasc access dev
C0177692|ICD9CM|PT|86.09|Other incision of skin and subcutaneous tissue
C0177692|ICD9CM|AB|86.09|Skin & subq incision NEC
C0177693|ICD9CM|HT|86.1|Diagnostic procedures on skin and subcutaneous tissue
C0177695|ICD9CM|PT|86.19|Other diagnostic procedures on skin and subcutaneous tissue
C0177695|ICD9CM|AB|86.19|Skin & subq dx proc NEC
C0177696|ICD9CM|HT|86.2|Excision or destruction of lesion or tissue of skin and subcutaneous tissue
C0177697|ICD9CM|PT|86.22|Excisional debridement of wound, infection, or burn
C0177697|ICD9CM|AB|86.22|Exc wound debridement
C0177698|ICD9CM|PT|86.23|Removal of nail, nail bed, or nail fold
C0177698|ICD9CM|AB|86.23|Nail removal
C0177699|ICD9CM|AB|86.24|Skin chemosurgery
C0177699|ICD9CM|PT|86.24|Chemosurgery of skin
C0177701|ICD9CM|PT|86.28|Nonexcisional debridement of wound, infection or burn
C0177701|ICD9CM|AB|86.28|Nonexcis debridement wnd
C0177702|ICD9CM|PT|86.3|Other local excision or destruction of lesion or tissue of skin and subcutaneous tissue
C0177702|ICD9CM|AB|86.3|Other local destruc skin
C0177705|ICD9CM|PT|86.61|Full-thickness skin graft to hand
C0177705|ICD9CM|AB|86.61|Full-thick hand skin grf
C0177706|ICD9CM|PT|86.62|Other skin graft to hand
C0177706|ICD9CM|AB|86.62|Hand skin graft NEC
C0177707|ICD9CM|PT|86.63|Full-thickness skin graft to other sites
C0177707|ICD9CM|AB|86.63|Full-thick skin grft NEC
C0177710|ICD9CM|PT|86.71|Cutting and preparation of pedicle grafts or flaps
C0177710|ICD9CM|AB|86.71|Cut & prep pedicle graft
C0177712|ICD9CM|PT|86.73|Attachment of pedicle or flap graft to hand
C0177712|ICD9CM|AB|86.73|Attach pedicle to hand
C0177713|ICD9CM|PT|86.74|Attachment of pedicle or flap graft to other sites
C0177713|ICD9CM|AB|86.74|Attach pedicle graft NEC
C0177714|ICD9CM|PT|86.75|Revision of pedicle or flap graft
C0177714|ICD9CM|AB|86.75|Revision of pedicle grft
C0177715|ICD9CM|HT|86.8|Other repair and reconstruction of skin and subcutaneous tissue
C0177715|ICD9CM|PT|86.89|Other repair and reconstruction of skin and subcutaneous tissue
C0177715|ICD9CM|AB|86.89|Skin repair & plasty NEC
C0177716|ICD9CM|PT|86.84|Relaxation of scar or web contracture of skin
C0177716|ICD9CM|AB|86.84|Relaxation of scar
C0177717|ICD9CM|HT|86.9|Other operations on skin and subcutaneous tissue
C0177717|ICD9CM|PT|86.99|Other operations on skin and subcutaneous tissue
C0177717|ICD9CM|AB|86.99|Skin & subq op NEC
C0177718|ICD9CM|PT|86.92|Electrolysis and other epilation of skin
C0177718|ICD9CM|AB|86.92|Epilation of skin
C0177719|ICD9CM|PT|87.04|Other tomography of head
C0177719|ICD9CM|AB|87.04|Head tomography NEC
C0177721|ICD9CM|AB|87.07|Contrast laryngogram
C0177721|ICD9CM|PT|87.07|Contrast laryngogram
C0177722|ICD9CM|PT|87.09|Other soft tissue x-ray of face, head, and neck
C0177722|ICD9CM|AB|87.09|Head soft tiss x-ray NEC
C0177723|ICD9CM|HT|87.1|Other x-ray of face, head, and neck
C0177726|ICD9CM|PT|87.16|Other x-ray of facial bones
C0177726|ICD9CM|AB|87.16|Facial bone x-ray NEC
C0177727|ICD9CM|PT|87.22|Other x-ray of cervical spine
C0177727|ICD9CM|AB|87.22|Cervical spine x-ray NEC
C0177728|ICD9CM|PT|87.23|Other x-ray of thoracic spine
C0177728|ICD9CM|AB|87.23|Thoracic spine x-ray NEC
C0177729|ICD9CM|PT|87.24|Other x-ray of lumbosacral spine
C0177729|ICD9CM|AB|87.24|Lumbosac spine x-ray NEC
C0177730|ICD9CM|PT|87.29|Other x-ray of spine
C0177730|ICD9CM|AB|87.29|Spinal x-ray NEC
C0177732|ICD9CM|PT|87.35|Contrast radiogram of mammary ducts
C0177732|ICD9CM|AB|87.35|Contr mammary ductogram
C0177733|ICD9CM|PT|87.39|Other soft tissue x-ray of chest wall
C0177733|ICD9CM|AB|87.39|Thorax sft tiss xray NEC
C0177735|ICD9CM|PT|87.42|Other tomography of thorax
C0177735|ICD9CM|AB|87.42|Thoracic tomography NEC
C0177737|ICD9CM|PT|87.49|Other chest x-ray
C0177737|ICD9CM|HT|87.4|Other x-ray of thorax
C0177737|ICD9CM|AB|87.49|Chest x-ray NEC
C0177738|ICD9CM|HT|87.5|Biliary tract x-ray
C0177739|ICD9CM|PT|87.51|Percutaneous hepatic cholangiogram
C0177739|ICD9CM|AB|87.51|Perc hepat Cholangiogram
C0177740|ICD9CM|PT|87.59|Other biliary tract x-ray
C0177740|ICD9CM|AB|87.59|Biliary tract x-ray NEC
C0177741|ICD9CM|HT|87.6|Other x-ray of digestive system
C0177742|ICD9CM|PT|87.65|Other x-ray of intestine
C0177742|ICD9CM|AB|87.65|Intestinal x-ray NEC
C0177743|ICD9CM|PT|87.69|Other digestive tract x-ray
C0177743|ICD9CM|AB|87.69|Digestive tract xray NEC
C0177745|ICD9CM|PT|87.72|Other nephrotomogram
C0177745|ICD9CM|AB|87.72|Nephrotomogram NEC
C0177746|ICD9CM|AB|87.75|Percutaneous pyelogram
C0177746|ICD9CM|PT|87.75|Percutaneous pyelogram
C0177747|ICD9CM|PT|87.77|Other cystogram
C0177747|ICD9CM|AB|87.77|Cystogram NEC
C0177749|ICD9CM|PT|87.79|Other x-ray of the urinary system
C0177749|ICD9CM|AB|87.79|Urinary system x-ray NEC
C0177750|ICD9CM|PT|87.82|Gas contrast hysterosalpingogram
C0177750|ICD9CM|AB|87.82|Gas hysterosalpingogram
C0177751|ICD9CM|PT|87.83|Opaque dye contrast hysterosalpingogram
C0177751|ICD9CM|AB|87.83|Dye hysterosalpingogram
C0177752|ICD9CM|PT|87.85|Other x-ray of fallopian tubes and uterus
C0177752|ICD9CM|AB|87.85|Tube & uterus x-ray NEC
C0177753|ICD9CM|PT|87.89|Other x-ray of female genital organs
C0177753|ICD9CM|AB|87.89|Female genital x-ray NEC
C0177754|ICD9CM|HT|87.9|X-ray of male genital organs
C0177755|ICD9CM|PT|87.91|Contrast seminal vesiculogram
C0177755|ICD9CM|AB|87.91|Contr semin vesiculogram
C0177756|ICD9CM|PT|87.92|Other x-ray of prostate and seminal vesicles
C0177756|ICD9CM|AB|87.92|Prostat/sem ves xray NEC
C0177757|ICD9CM|AB|87.93|Contrast epididymogram
C0177757|ICD9CM|PT|87.93|Contrast epididymogram
C0177758|ICD9CM|AB|87.94|Contrast vasogram
C0177758|ICD9CM|PT|87.94|Contrast vasogram
C0177759|ICD9CM|PT|87.95|Other x-ray of epididymis and vas deferens
C0177759|ICD9CM|AB|87.95|Epididymis/vas x-ray NEC
C0177760|ICD9CM|PT|87.99|Other x-ray of male genital organs
C0177760|ICD9CM|AB|87.99|Male genital x-ray NEC
C0177761|ICD9CM|HT|88.0|Soft tissue x-ray of abdomen
C0177762|ICD9CM|PT|88.02|Other abdomen tomography
C0177762|ICD9CM|AB|88.02|Abdominal tomography NEC
C0177763|ICD9CM|PT|88.09|Other soft tissue x-ray of abdominal wall
C0177763|ICD9CM|AB|88.09|Abdominal wall x-ray NEC
C0177764|ICD9CM|PT|88.11|Pelvic opaque dye contrast radiography
C0177764|ICD9CM|AB|88.11|Pelvic dye contrast xray
C0177766|ICD9CM|PT|88.13|Other peritoneal pneumogram
C0177766|ICD9CM|AB|88.13|Periton pneumogram NEC
C0177767|ICD9CM|PT|88.15|Retroperitoneal pneumogram
C0177767|ICD9CM|AB|88.15|Retroperiton pneumogram
C0177768|ICD9CM|PT|88.16|Other retroperitoneal x-ray
C0177768|ICD9CM|AB|88.16|Retroperitoneal xray NEC
C0177769|ICD9CM|HT|88.2|Skeletal x-ray of extremities and pelvis
C0177770|ICD9CM|PT|88.21|Skeletal x-ray of shoulder and upper arm
C0177770|ICD9CM|AB|88.21|Skl xray-shoulder/up arm
C0177771|ICD9CM|PT|88.26|Other skeletal x-ray of pelvis and hip
C0177771|ICD9CM|AB|88.26|Skel xray-pelvis/hip NEC
C0177772|ICD9CM|PT|88.27|Skeletal x-ray of thigh, knee, and lower leg
C0177772|ICD9CM|AB|88.27|Skel xray-thigh/knee/leg
C0177773|ICD9CM|HT|88.3|Other x-ray
C0177774|ICD9CM|AB|88.33|Other skeletal x-ray
C0177774|ICD9CM|PT|88.33|Other skeletal x-ray
C0177776|ICD9CM|PT|88.35|Other soft tissue x-ray of upper limb
C0177776|ICD9CM|AB|88.35|Up limb sft tis xray NEC
C0177778|ICD9CM|PT|88.37|Other soft tissue x-ray of lower limb
C0177778|ICD9CM|AB|88.37|Lo limb sft tis xray NEC
C0177779|ICD9CM|PT|88.38|Other computerized axial tomography
C0177779|ICD9CM|AB|88.38|Other C.A.T. scan
C0177780|ICD9CM|PT|88.44|Arteriography of other intrathoracic vessels
C0177780|ICD9CM|AB|88.44|Contr thor arteriogr NEC
C0177782|ICD9CM|PT|88.47|Arteriography of other intra-abdominal arteries
C0177782|ICD9CM|AB|88.47|Contr abd arteriogrm NEC
C0177783|ICD9CM|PT|88.48|Arteriography of femoral and other lower extremity arteries
C0177783|ICD9CM|AB|88.48|Contrast arteriogram-leg
C0177784|ICD9CM|PT|88.49|Arteriography of other specified sites
C0177784|ICD9CM|AB|88.49|Contrast arteriogram NEC
C0177785|ICD9CM|HT|88.5|Angiocardiography using contrast material
C0177789|ICD9CM|PT|88.57|Other and unspecified coronary arteriography
C0177789|ICD9CM|AB|88.57|Coronary arteriogram NEC
C0177790|ICD9CM|PT|88.61|Phlebography of veins of head and neck using contrast material
C0177790|ICD9CM|AB|88.61|Contr phlebogram-hd/neck
C0177791|ICD9CM|PT|88.62|Phlebography of pulmonary veins using contrast material
C0177791|ICD9CM|AB|88.62|Contr phlebogram-pulmon
C0177792|ICD9CM|PT|88.63|Phlebography of other intrathoracic veins using contrast material
C0177792|ICD9CM|AB|88.63|Thorac contr phlebog NEC
C0177793|ICD9CM|PT|88.64|Phlebography of the portal venous system using contrast material
C0177793|ICD9CM|AB|88.64|Portal contr phlebogram
C0177794|ICD9CM|PT|88.65|Phlebography of other Intra-Abdominal veins using contrast material
C0177794|ICD9CM|AB|88.65|Abd contr phlebogram NEC
C0177795|ICD9CM|PT|88.66|Phlebography of femoral and other lower extremity veins using contrast material
C0177795|ICD9CM|AB|88.66|Contrast phlebogram-leg
C0177796|ICD9CM|PT|88.67|Phlebography of other specified sites using contrast material
C0177796|ICD9CM|AB|88.67|Contrast phlebogram NEC
C0177800|ICD9CM|PT|88.79|Other diagnostic ultrasound
C0177800|ICD9CM|AB|88.79|Dx ultrasound NEC
C0177801|ICD9CM|HT|88.9|Other diagnostic imaging
C0177804|ICD9CM|AB|88.98|Bone mineral density
C0177804|ICD9CM|PT|88.98|Bone mineral density studies
C0177805|ICD9CM|HT|89.0|Diagnostic interview, consultation, and evaluation
C0177806|ICD9CM|PT|89.01|Interview and evaluation, described as brief
C0177806|ICD9CM|AB|89.01|Brief interview & evalua
C0177807|ICD9CM|PT|89.02|Interview and evaluation, described as limited
C0177807|ICD9CM|AB|89.02|Limited interview/evalua
C0177808|ICD9CM|PT|89.03|Interview and evaluation, described as comprehensive
C0177808|ICD9CM|AB|89.03|Comprehen interview/eval
C0177809|ICD9CM|PT|89.04|Other interview and evaluation
C0177809|ICD9CM|AB|89.04|Interview & evaluat NEC
C0177812|ICD9CM|PT|89.08|Other consultation
C0177812|ICD9CM|AB|89.08|Consultation NEC
C0177813|ICD9CM|HT|89.1|Anatomic and physiologic measurements and manual examinations -- nervous system and sense organs
C0177814|ICD9CM|PT|89.15|Other nonoperative neurologic function tests
C0177814|ICD9CM|AB|89.15|Neurologic func test NEC
C0177815|ICD9CM|PT|89.18|Other sleep disorder function tests
C0177815|ICD9CM|AB|89.18|Oth sleep dis funct test
C0177816|ICD9CM|HT|89.2|Anatomic and physiologic measurements and manual examinations -- genitourinary system
C0177820|ICD9CM|PT|89.29|Other nonoperative genitourinary system measurements
C0177820|ICD9CM|AB|89.29|Other gu system exams
C0177821|ICD9CM|HT|89.3|Other anatomic and physiologic measurements and manual examinations
C0177823|ICD9CM|PT|89.44|Other cardiovascular stress test
C0177823|ICD9CM|AB|89.44|Cardiac stress test NEC
C0177826|ICD9CM|PT|89.48|Artificial pacemaker voltage or amperage threshold check
C0177826|ICD9CM|AB|89.48|Pacemaker volt threshold
C0177828|ICD9CM|HT|89.5|Other nonoperative cardiac and vascular diagnostic procedures
C0177829|ICD9CM|PT|89.50|Ambulatory cardiac monitoring
C0177829|ICD9CM|AB|89.50|Ambu cardiac monitoring
C0177831|ICD9CM|PT|89.54|Electrographic monitoring
C0177831|ICD9CM|AB|89.54|Electrocardiograph monit
C0177834|ICD9CM|PT|89.66|Measurement of mixed venous blood gases
C0177834|ICD9CM|AB|89.66|Mix venous bld gas meas
C0177836|ICD9CM|HT|90.0|Microscopic examination of specimen from nervous system and of spinal fluid
C0177837|ICD9CM|PT|90.01|Microscopic examination of specimen from nervous system and of spinal fluid, bacterial smear
C0177837|ICD9CM|AB|90.01|Bact smear-nervous syst
C0177838|ICD9CM|PT|90.02|Microscopic examination of specimen from nervous system and of spinal fluid, culture
C0177838|ICD9CM|AB|90.02|Culture-nervous syst
C0177839|ICD9CM|PT|90.03|Microscopic examination of specimen from nervous system and of spinal fluid, culture and sensitivity
C0177839|ICD9CM|AB|90.03|C & s-nervous syst
C0177840|ICD9CM|PT|90.04|Microscopic examination of specimen from nervous system and of spinal fluid, parasitology
C0177840|ICD9CM|AB|90.04|Parasitology-nerv syst
C0177841|ICD9CM|PT|90.05|Microscopic examination of specimen from nervous system and of spinal fluid, toxicology
C0177841|ICD9CM|AB|90.05|Toxicology-nervous syst
C0177842|ICD9CM|PT|90.06|Microscopic examination of specimen from nervous system and of spinal fluid, cell block and Papanicolaou smear
C0177842|ICD9CM|AB|90.06|Cell blk/pap-nervous sys
C0177843|ICD9CM|PT|90.09|Microscopic examination of specimen from nervous system and of spinal fluid, other microscopic examination
C0177843|ICD9CM|AB|90.09|Micro exam-nervous NEC
C0177850|ICD9CM|PT|90.16|Microscopic examination of specimen from endocrine gland, not elsewhere classified, cell block and Papanicolaou smear
C0177850|ICD9CM|AB|90.16|Cell block/pap-endocrine
C0177852|ICD9CM|HT|90.2|Microscopic examination of specimen from eye
C0177853|ICD9CM|PT|90.21|Microscopic examination of specimen from eye, bacterial smear
C0177853|ICD9CM|AB|90.21|Bact smear-eye
C0177855|ICD9CM|PT|90.23|Microscopic examination of specimen from eye, culture and sensitivity
C0177855|ICD9CM|AB|90.23|C & s-eye
C0177856|ICD9CM|PT|90.24|Microscopic examination of specimen from eye, parasitology
C0177856|ICD9CM|AB|90.24|Parasitology-eye
C0177857|ICD9CM|PT|90.25|Microscopic examination of specimen from eye, toxicology
C0177857|ICD9CM|AB|90.25|Toxicology-eye
C0177858|ICD9CM|PT|90.26|Microscopic examination of specimen from eye, cell block and Papanicolaou smear
C0177858|ICD9CM|AB|90.26|Cell block/pap-eye
C0177859|ICD9CM|PT|90.29|Microscopic examination of specimen from eye, other microscopic examination
C0177859|ICD9CM|AB|90.29|Micro exam-eye NEC
C0177860|ICD9CM|HT|90.3|Microscopic examination of specimen from ear, nose, throat, and larynx
C0177861|ICD9CM|PT|90.31|Microscopic examination of specimen from ear, nose, throat, and larynx, bacterial smear
C0177861|ICD9CM|AB|90.31|Bact smear-ent/larynx
C0177862|ICD9CM|PT|90.32|Microscopic examination of specimen from ear, nose, throat, and larynx, culture
C0177862|ICD9CM|AB|90.32|Culture-ent/larynx
C0177863|ICD9CM|PT|90.33|Microscopic examination of specimen from ear, nose, throat, and larynx, culture and sensitivity
C0177863|ICD9CM|AB|90.33|C & s-ent/larynx
C0177864|ICD9CM|PT|90.34|Microscopic examination of specimen from ear, nose, throat, and larynx, parasitology
C0177864|ICD9CM|AB|90.34|Parasitology-ent/larynx
C0177865|ICD9CM|PT|90.35|Microscopic examination of specimen from ear, nose, throat, and larynx, toxicology
C0177865|ICD9CM|AB|90.35|Toxicology-ent/larynx
C0177866|ICD9CM|PT|90.36|Microscopic examination of specimen from ear, nose, throat, and larynx, cell block and Papanicolaou smear
C0177866|ICD9CM|AB|90.36|Cell block/pap-ent/laryn
C0177867|ICD9CM|PT|90.39|Microscopic examination of specimen from ear, nose, throat, and larynx, other microscopic examination
C0177867|ICD9CM|AB|90.39|Micro exam-ent/laryn NEC
C0177868|ICD9CM|HT|90.4|Microscopic examination of specimen from trachea, bronchus, pleura, lung, and other thoracic specimen, and of sputum
C0177869|ICD9CM|PT|90.41|Microscopic examination of specimen from trachea, bronchus, pleura, lung, and other thoracic specimen, and of sputum, bacterial smear
C0177869|ICD9CM|AB|90.41|Bact smear-lower resp
C0177870|ICD9CM|PT|90.42|Microscopic examination of specimen from trachea, bronchus, pleura, lung, and other thoracic specimen, and of sputum, culture
C0177870|ICD9CM|AB|90.42|Culture-lower resp
C0177871|ICD9CM|PT|90.43|Microscopic examination of specimen from trachea, bronchus, pleura, lung, and other thoracic specimen, and of sputum, culture and sensitivity
C0177871|ICD9CM|AB|90.43|C & s-lower resp
C0177872|ICD9CM|PT|90.44|Microscopic examination of specimen from trachea, bronchus, pleura, lung, and other thoracic specimen, and of sputum, parasitology
C0177872|ICD9CM|AB|90.44|Parasitology-lower resp
C0177873|ICD9CM|PT|90.45|Microscopic examination of specimen from trachea, bronchus, pleura, lung, and other thoracic specimen, and of sputum, toxicology
C0177873|ICD9CM|AB|90.45|Toxicology-lower resp
C0177874|ICD9CM|PT|90.46|Microscopic examination of specimen from trachea, bronchus, pleura, lung, and other thoracic specimen, and of sputum, cell block and Papanicolaou smear
C0177874|ICD9CM|AB|90.46|Cell block/pap-lowr resp
C0177875|ICD9CM|PT|90.49|Microscopic examination of specimen from trachea, bronchus, pleura, lung, and other thoracic specimen, and of sputum, other microscopic examination
C0177875|ICD9CM|AB|90.49|Micro exam-lowr resp NEC
C0177876|ICD9CM|HT|90.5|Microscopic examination of blood
C0177877|ICD9CM|PT|90.51|Microscopic examination of blood, bacterial smear
C0177877|ICD9CM|AB|90.51|Bact smear-blood
C0177879|ICD9CM|PT|90.53|Microscopic examination of blood, culture and sensitivity
C0177879|ICD9CM|AB|90.53|C & s-blood
C0177880|ICD9CM|PT|90.54|Microscopic examination of blood, parasitology
C0177880|ICD9CM|AB|90.54|Parasitology-blood
C0177881|ICD9CM|AB|90.55|Toxicology-blood
C0177881|ICD9CM|PT|90.55|Microscopic examination of blood, toxicology
C0177882|ICD9CM|PT|90.56|Microscopic examination of blood, cell block and Papanicolaou smear
C0177882|ICD9CM|AB|90.56|Cell block/pap-blood
C0177883|ICD9CM|PT|90.59|Microscopic examination of blood, other microscopic examination
C0177883|ICD9CM|AB|90.59|Micro exam-blood NEC
C0177884|ICD9CM|HT|90.6|Microscopic examination of specimen from spleen and of bone marrow
C0177885|ICD9CM|PT|90.61|Microscopic examination of specimen from spleen and of bone marrow, bacterial smear
C0177885|ICD9CM|AB|90.61|Bact smear-spleen/marrow
C0177886|ICD9CM|PT|90.62|Microscopic examination of specimen from spleen and of bone marrow, culture
C0177886|ICD9CM|AB|90.62|Culture-spleen/marrow
C0177887|ICD9CM|PT|90.63|Microscopic examination of specimen from spleen and of bone marrow, culture and sensitivity
C0177887|ICD9CM|AB|90.63|C & s-spleen/marrow
C0177888|ICD9CM|PT|90.64|Microscopic examination of specimen from spleen and of bone marrow, parasitology
C0177888|ICD9CM|AB|90.64|Parasitol-spleen/marrow
C0177889|ICD9CM|PT|90.65|Microscopic examination of specimen from spleen and of bone marrow, toxicology
C0177889|ICD9CM|AB|90.65|Toxicology-spleen/marrow
C0177890|ICD9CM|PT|90.66|Microscopic examination of specimen from spleen and of bone marrow, cell block and Papanicolaou smear
C0177890|ICD9CM|AB|90.66|Cell blk/pap-spleen/marr
C0177891|ICD9CM|PT|90.69|Microscopic examination of specimen from spleen and of bone marrow, other microscopic examination
C0177891|ICD9CM|AB|90.69|Micro exam-spln/marr NEC
C0177892|ICD9CM|HT|90.7|Microscopic examination of specimen from lymph node and of lymph
C0177893|ICD9CM|PT|90.71|Microscopic examination of specimen from lymph node and of lymph, bacterial smear
C0177893|ICD9CM|AB|90.71|Bact smear-lymph system
C0177894|ICD9CM|PT|90.72|Microscopic examination of specimen from lymph node and of lymph, culture
C0177894|ICD9CM|AB|90.72|Culture-lymph system
C0177895|ICD9CM|PT|90.73|Microscopic examination of specimen from lymph node and of lymph, culture and sensitivity
C0177895|ICD9CM|AB|90.73|C & s-lymph system
C0177896|ICD9CM|PT|90.74|Microscopic examination of specimen from lymph node and of lymph, parasitology
C0177896|ICD9CM|AB|90.74|Parasitology-lymph sys
C0177897|ICD9CM|PT|90.75|Microscopic examination of specimen from lymph node and of lymph, toxicology
C0177897|ICD9CM|AB|90.75|Toxicology-lymph system
C0177898|ICD9CM|PT|90.76|Microscopic examination of specimen from lymph node and of lymph, cell block and Papanicolaou smear
C0177898|ICD9CM|AB|90.76|Cell blk/pap-lymph sys
C0177899|ICD9CM|PT|90.79|Microscopic examination of specimen from lymph node and of lymph, other microscopic examination
C0177899|ICD9CM|AB|90.79|Micro exam-lymph sys NEC
C0177900|ICD9CM|HT|90.8|Microscopic examination of specimen from upper gastrointestinal tract and of vomitus
C0177901|ICD9CM|PT|90.81|Microscopic examination of specimen from upper gastrointestinal tract and of vomitus, bacterial smear
C0177901|ICD9CM|AB|90.81|Bact smear-upper GI
C0177902|ICD9CM|PT|90.82|Microscopic examination of specimen from upper gastrointestinal tract and of vomitus, culture
C0177902|ICD9CM|AB|90.82|Culture-upper GI
C0177903|ICD9CM|PT|90.83|Microscopic examination of specimen from upper gastrointestinal tract and of vomitus, culture and sensitivity
C0177903|ICD9CM|AB|90.83|C & s-upper GI
C0177904|ICD9CM|PT|90.84|Microscopic examination of specimen from upper gastrointestinal tract and of vomitus, parasitology
C0177904|ICD9CM|AB|90.84|Parasitology-upper GI
C0177905|ICD9CM|PT|90.85|Microscopic examination of specimen from upper gastrointestinal tract and of vomitus, toxicology
C0177905|ICD9CM|AB|90.85|Toxicology-upper GI
C0177906|ICD9CM|PT|90.86|Microscopic examination of specimen from upper gastrointestinal tract and of vomitus, cell block and Papanicolaou smear
C0177906|ICD9CM|AB|90.86|Cell blk/pap-upper GI
C0177907|ICD9CM|PT|90.89|Microscopic examination of specimen from upper gastrointestinal tract and of vomitus, other microscopic examination
C0177907|ICD9CM|AB|90.89|Micro exam-upper GI NEC
C0177908|ICD9CM|HT|90.9|Microscopic examination of specimen from lower gastrointestinal tract and of stool
C0177909|ICD9CM|PT|90.91|Microscopic examination of specimen from lower gastrointestinal tract and of stool, bacterial smear
C0177909|ICD9CM|AB|90.91|Bact smear-lower GI
C0177910|ICD9CM|PT|90.92|Microscopic examination of specimen from lower gastrointestinal tract and of stool, culture
C0177910|ICD9CM|AB|90.92|Culture-lower GI
C0177911|ICD9CM|PT|90.93|Microscopic examination of specimen from lower gastrointestinal tract and of stool, culture and sensitivity
C0177911|ICD9CM|AB|90.93|C & s-lower GI
C0177912|ICD9CM|PT|90.94|Microscopic examination of specimen from lower gastrointestinal tract and of stool, parasitology
C0177912|ICD9CM|AB|90.94|Parasitology-lower GI
C0177913|ICD9CM|PT|90.95|Microscopic examination of specimen from lower gastrointestinal tract and of stool, toxicology
C0177913|ICD9CM|AB|90.95|Toxicology-lower GI
C0177914|ICD9CM|PT|90.96|Microscopic examination of specimen from lower gastrointestinal tract and of stool, cell block and Papanicolaou smear
C0177914|ICD9CM|AB|90.96|Cell blk/pap-lower GI
C0177915|ICD9CM|PT|90.99|Microscopic examination of specimen from lower gastrointestinal tract and of stool, other microscopic examination
C0177915|ICD9CM|AB|90.99|Micro exam-lower GI NEC
C0177916|ICD9CM|HT|91.0|Microscopic examination of specimen from liver, biliary tract, and pancreas
C0177917|ICD9CM|PT|91.01|Microscopic examination of specimen from liver, biliary tract, and pancreas, bacterial smear
C0177917|ICD9CM|AB|91.01|Bact smear-bili/pancreas
C0177918|ICD9CM|PT|91.02|Microscopic examination of specimen from liver, biliary tract, and pancreas, culture
C0177918|ICD9CM|AB|91.02|Culture-bili/pancreas
C0177919|ICD9CM|PT|91.03|Microscopic examination of specimen from liver, biliary tract, and pancreas, culture and sensitivity
C0177919|ICD9CM|AB|91.03|C & s-bili/pancreas
C0177920|ICD9CM|PT|91.04|Microscopic examination of specimen from liver, biliary tract, and pancreas, parasitology
C0177920|ICD9CM|AB|91.04|Parasitology-bili/pancr
C0177921|ICD9CM|PT|91.05|Microscopic examination of specimen from liver, biliary tract, and pancreas, toxicology
C0177921|ICD9CM|AB|91.05|Toxicology-bili/pancreas
C0177922|ICD9CM|PT|91.06|Microscopic examination of specimen from liver, biliary tract, and pancreas, cell block and Papanicolaou smear
C0177922|ICD9CM|AB|91.06|Cell blk/pap-bili/pancre
C0177923|ICD9CM|PT|91.09|Microscopic examination of specimen from liver, biliary tract, and pancreas, other microscopic examination
C0177923|ICD9CM|AB|91.09|Micro exam-bili/panc NEC
C0177924|ICD9CM|HT|91.1|Microscopic examination of peritoneal and retroperitoneal specimen
C0177925|ICD9CM|PT|91.11|Microscopic examination of peritoneal and retroperitoneal specimen, bacterial smear
C0177925|ICD9CM|AB|91.11|Bact smear-peritoneum
C0177926|ICD9CM|PT|91.12|Microscopic examination of peritoneal and retroperitoneal specimen, culture
C0177926|ICD9CM|AB|91.12|Culture-peritoneum
C0177927|ICD9CM|PT|91.13|Microscopic examination of peritoneal and retroperitoneal specimen, culture and sensitivity
C0177927|ICD9CM|AB|91.13|C & s-peritoneum
C0177928|ICD9CM|PT|91.14|Microscopic examination of peritoneal and retroperitoneal specimen, parasitology
C0177928|ICD9CM|AB|91.14|Parasitology-peritoneum
C0177929|ICD9CM|PT|91.15|Microscopic examination of peritoneal and retroperitoneal specimen, toxicology
C0177929|ICD9CM|AB|91.15|Toxicology-peritoneum
C0177930|ICD9CM|PT|91.16|Microscopic examination of peritoneal and retroperitoneal specimen, cell block and Papanicolaou smear
C0177930|ICD9CM|AB|91.16|Cell blk/pap-peritoneum
C0177931|ICD9CM|PT|91.19|Microscopic examination of peritoneal and retroperitoneal specimen, other microscopic examination
C0177931|ICD9CM|AB|91.19|Micro exam-periton NEC
C0177932|ICD9CM|HT|91.2|Microscopic examination of specimen from kidney, ureter, perirenal and periureteral tissue
C0177933|ICD9CM|PT|91.21|Microscopic examination of specimen from kidney, ureter, perirenal and periureteral tissue, bacterial smear
C0177933|ICD9CM|AB|91.21|Bact smear-upper urinary
C0177934|ICD9CM|PT|91.22|Microscopic examination of specimen from kidney, ureter, perirenal and periureteral tissue, culture
C0177934|ICD9CM|AB|91.22|Culture-upper urinary
C0177935|ICD9CM|PT|91.23|Microscopic examination of specimen from kidney, ureter, perirenal and periureteral tissue, culture and sensitivity
C0177935|ICD9CM|AB|91.23|C & s-upper urinary
C0177936|ICD9CM|PT|91.24|Microscopic examination of specimen from kidney, ureter, perirenal and periureteral tissue, parasitology
C0177936|ICD9CM|AB|91.24|Parasitology-upper urin
C0177937|ICD9CM|PT|91.25|Microscopic examination of specimen from kidney, ureter, perirenal and periureteral tissue, toxicology
C0177937|ICD9CM|AB|91.25|Toxicology-upper urinary
C0177938|ICD9CM|PT|91.26|Microscopic examination of specimen from kidney, ureter, perirenal and periureteral tissue, cell block and Papanicolaou smear
C0177938|ICD9CM|AB|91.26|Cell blk/pap-upper urin
C0177939|ICD9CM|PT|91.29|Microscopic examination of specimen from kidney, ureter, perirenal and periureteral tissue, other microscopic examination
C0177939|ICD9CM|AB|91.29|Micro exam-uppr urin NEC
C0177940|ICD9CM|HT|91.3|Microscopic examination of specimen from bladder, urethra, prostate, seminal vesicle, perivesical tissue, and of urine and semen
C0177941|ICD9CM|PT|91.31|Microscopic examination of specimen from bladder, urethra, prostate, seminal vesicle, perivesical tissue, and of urine and semen, bacterial smear
C0177941|ICD9CM|AB|91.31|Bact smear-lower urinary
C0177942|ICD9CM|PT|91.32|Microscopic examination of specimen from bladder, urethra, prostate, seminal vesicle, perivesical tissue, and of urine and semen, culture
C0177942|ICD9CM|AB|91.32|Culture-lower urinary
C0177943|ICD9CM|PT|91.33|Microscopic examination of specimen from bladder, urethra, prostate, seminal vesicle, perivesical tissue, and of urine and semen, culture and sensitivity
C0177943|ICD9CM|AB|91.33|C & s-lower urinary
C0177944|ICD9CM|PT|91.34|Microscopic examination of specimen from bladder, urethra, prostate, seminal vesicle, perivesical tissue, and of urine and semen, parasitology
C0177944|ICD9CM|AB|91.34|Parasitlolgy-lower urin
C0177945|ICD9CM|PT|91.35|Microscopic examination of specimen from bladder, urethra, prostate, seminal vesicle, perivesical tissue, and of urine and semen, toxicology
C0177945|ICD9CM|AB|91.35|Toxicology-lower urinary
C0177946|ICD9CM|PT|91.36|Microscopic examination of specimen from bladder, urethra, prostate, seminal vesicle, perivesical tissue, and of urine and semen, cell block and Papanicolaou smear
C0177946|ICD9CM|AB|91.36|Cell blk/pap-lower urin
C0177947|ICD9CM|PT|91.39|Microscopic examination of specimen from bladder, urethra, prostate, seminal vesicle, perivesical tissue, and of urine and semen, other microscopic examination
C0177947|ICD9CM|AB|91.39|Micro exam-low urin NEC
C0177948|ICD9CM|HT|91.4|Microscopic examination of specimen from female genital tract
C0177949|ICD9CM|PT|91.41|Microscopic examination of specimen from female genital tract, bacterial smear
C0177949|ICD9CM|AB|91.41|Bact smear-female genit
C0177950|ICD9CM|PT|91.42|Microscopic examination of specimen from female genital tract, culture
C0177950|ICD9CM|AB|91.42|Culture-female genital
C0177951|ICD9CM|PT|91.43|Microscopic examination of specimen from female genital tract, culture and sensitivity
C0177951|ICD9CM|AB|91.43|C & s-female genital
C0177952|ICD9CM|PT|91.44|Microscopic examination of specimen from female genital tract, parasitology
C0177952|ICD9CM|AB|91.44|Parasitology-female gen
C0177953|ICD9CM|PT|91.45|Microscopic examination of specimen from female genital tract, toxicology
C0177953|ICD9CM|AB|91.45|Toxicology-female genit
C0177954|ICD9CM|PT|91.46|Microscopic examination of specimen from female genital tract, cell block and Papanicolaou smear
C0177954|ICD9CM|AB|91.46|Cell blk/pap-female gen
C0177955|ICD9CM|PT|91.49|Microscopic examination of specimen from female genital tract, other microscopic examination
C0177955|ICD9CM|AB|91.49|Micro exam-femal gen NEC
C0177956|ICD9CM|HT|91.5|Microscopic examination of specimen from musculoskeletal system and of joint fluid
C0177957|ICD9CM|PT|91.51|Microscopic examination of specimen from musculoskeletal system and of joint fluid, bacterial smear
C0177957|ICD9CM|AB|91.51|Bact smear-musculoskel
C0177958|ICD9CM|PT|91.52|Microscopic examination of specimen from musculoskeletal system and of joint fluid, culture
C0177958|ICD9CM|AB|91.52|Culture-musculoskeletal
C0177959|ICD9CM|PT|91.53|Microscopic examination of specimen from musculoskeletal system and of joint fluid, culture and sensitivity
C0177959|ICD9CM|AB|91.53|C & s-musculoskeletal
C0177960|ICD9CM|PT|91.54|Microscopic examination of specimen from musculoskeletal system and of joint fluid, parasitology
C0177960|ICD9CM|AB|91.54|Parasitology-musculoskel
C0177961|ICD9CM|PT|91.55|Microscopic examination of specimen from musculoskeletal system and of joint fluid, toxicology
C0177961|ICD9CM|AB|91.55|Toxicology-musculoskel
C0177962|ICD9CM|PT|91.56|Microscopic examination of specimen from musculoskeletal system and of joint fluid, cell block and Papanicolaou smear
C0177962|ICD9CM|AB|91.56|Cell blk/pap-musculoskel
C0177963|ICD9CM|PT|91.59|Microscopic examination of specimen from musculoskeletal system and of joint fluid, other microscopic examination
C0177963|ICD9CM|AB|91.59|Micro exam-musculosk NEC
C0177964|ICD9CM|HT|91.6|Microscopic examination of specimen from skin and other integument
C0177965|ICD9CM|PT|91.61|Microscopic examination of specimen from skin and other integument, bacterial smear
C0177965|ICD9CM|AB|91.61|Bact smear-integument
C0177966|ICD9CM|PT|91.62|Microscopic examination of specimen from skin and other integument, culture
C0177966|ICD9CM|AB|91.62|Culture-integument
C0177967|ICD9CM|PT|91.63|Microscopic examination of specimen from skin and other integument, culture and sensitivity
C0177967|ICD9CM|AB|91.63|C & s-integument
C0177968|ICD9CM|PT|91.64|Microscopic examination of specimen from skin and other integument, parasitology
C0177968|ICD9CM|AB|91.64|Parasitology-integument
C0177969|ICD9CM|PT|91.65|Microscopic examination of specimen from skin and other integument, toxicology
C0177969|ICD9CM|AB|91.65|Toxicology-integument
C0177970|ICD9CM|PT|91.66|Microscopic examination of specimen from skin and other integument, cell block and Papanicolaou smear
C0177970|ICD9CM|AB|91.66|Cell blk/pap-integument
C0177971|ICD9CM|PT|91.69|Microscopic examination of specimen from skin and other integument, other microscopic examination
C0177971|ICD9CM|AB|91.69|Micro exam-integumen NEC
C0177972|ICD9CM|HT|91.7|Microscopic examination of specimen from operative wound
C0177973|ICD9CM|PT|91.71|Microscopic examination of specimen from operative wound, bacterial smear
C0177973|ICD9CM|AB|91.71|Bact smear-op wound
C0177974|ICD9CM|PT|91.72|Microscopic examination of specimen from operative wound, culture
C0177974|ICD9CM|AB|91.72|Culture-op wound
C0177975|ICD9CM|PT|91.73|Microscopic examination of specimen from operative wound, culture and sensitivity
C0177975|ICD9CM|AB|91.73|C & s-op wound
C0177976|ICD9CM|PT|91.74|Microscopic examination of specimen from operative wound, parasitology
C0177976|ICD9CM|AB|91.74|Parasitology-op wound
C0177977|ICD9CM|PT|91.75|Microscopic examination of specimen from operative wound, toxicology
C0177977|ICD9CM|AB|91.75|Toxicology-op wound
C0177978|ICD9CM|PT|91.76|Microscopic examination of specimen from operative wound, cell block and Papanicolaou smear
C0177978|ICD9CM|AB|91.76|Cell blk/pap-op wound
C0177979|ICD9CM|PT|91.79|Microscopic examination of specimen from operative wound, other microscopic examination
C0177979|ICD9CM|AB|91.79|Micro exam-op wound NEC
C0177980|ICD9CM|HT|91.8|Microscopic examination of specimen from other site
C0177981|ICD9CM|PT|91.81|Microscopic examination of specimen from other site, bacterial smear
C0177981|ICD9CM|AB|91.81|Bact smear NEC
C0177982|ICD9CM|PT|91.82|Microscopic examination of specimen from other site, culture
C0177982|ICD9CM|AB|91.82|Culture NEC
C0177983|ICD9CM|PT|91.83|Microscopic examination of specimen from other site, culture and sensitivity
C0177983|ICD9CM|AB|91.83|C & s NEC
C0177984|ICD9CM|PT|91.84|Microscopic examination of specimen from other site, parasitology
C0177984|ICD9CM|AB|91.84|Parasitology NEC
C0177985|ICD9CM|PT|91.86|Microscopic examination of specimen from other site, cell block and Papanicolaou smear
C0177985|ICD9CM|AB|91.86|Cell blk/pap NEC
C0177986|ICD9CM|PT|91.89|Microscopic examination of specimen from other site, other microscopic examination
C0177986|ICD9CM|AB|91.89|Micro exam NEC
C0177987|ICD9CM|HT|91.9|Microscopic examination of specimen from unspecified site
C0177988|ICD9CM|PT|91.91|Microscopic examination of specimen from unspecified site, bacterial smear
C0177988|ICD9CM|AB|91.91|Bact smear NOS
C0177989|ICD9CM|AB|91.92|Culture NOS
C0177989|ICD9CM|PT|91.92|Microscopic examination of specimen from unspecified site, culture
C0177990|ICD9CM|PT|91.93|Microscopic examination of specimen from unspecified site, culture and sensitivity
C0177990|ICD9CM|AB|91.93|C & s NOS
C0177991|ICD9CM|AB|91.94|Parasitology NOS
C0177991|ICD9CM|PT|91.94|Microscopic examination of specimen from unspecified site, parasitology
C0177992|ICD9CM|PT|91.96|Microscopic examination of specimen from unspecified site, cell block and Papanicolaou smear
C0177992|ICD9CM|AB|91.96|Cell blk/pap NOS
C0177993|ICD9CM|PT|91.99|Microscopic examination of specimen from unspecified site, other microscopic examination
C0177993|ICD9CM|AB|91.99|Micro exam NOS
C0177994|ICD9CM|HT|92.0|Radioisotope scan and function study
C0177996|ICD9CM|PT|92.04|Gastrointestinal scan and radioisotope function study
C0177996|ICD9CM|AB|92.04|GI scan & isotope funct
C0177997|ICD9CM|PT|92.05|Cardiovascular and hematopoietic scan and radioisotope function study
C0177997|ICD9CM|AB|92.05|C-vasc scan/isotop funct
C0177998|ICD9CM|PT|92.09|Other radioisotope function studies
C0177998|ICD9CM|AB|92.09|Other isotope function
C0177999|ICD9CM|HT|92.1|Other radioisotope scan
C0178000|ICD9CM|PT|92.12|Scan of other sites of head
C0178000|ICD9CM|AB|92.12|Head scan NEC
C0178001|ICD9CM|AB|92.19|Scan of other sites
C0178001|ICD9CM|PT|92.19|Scan of other sites
C0178002|ICD9CM|HT|92.2|Therapeutic radiology and nuclear medicine
C0178003|ICD9CM|PT|92.23|Radioisotopic teleradiotherapy
C0178003|ICD9CM|AB|92.23|Radioisot teleradiother
C0178005|ICD9CM|PT|92.26|Teleradiotherapy of other particulate radiation
C0178005|ICD9CM|AB|92.26|Particul teleradioth NEC
C0178006|ICD9CM|PT|92.27|Implantation or insertion of radioactive elements
C0178006|ICD9CM|AB|92.27|Radioactive elem implant
C0178007|ICD9CM|PT|92.29|Other radiotherapeutic procedure
C0178007|ICD9CM|AB|92.29|Radiotherapeut proc NEC
C0178010|ICD9CM|PT|93.09|Other diagnostic physical therapy procedure
C0178010|ICD9CM|AB|93.09|Other dx pt procedure
C0178012|ICD9CM|PT|93.12|Other active musculoskeletal exercise
C0178012|ICD9CM|AB|93.12|Activ musculosk exer NEC
C0178013|ICD9CM|AB|93.15|Mobilization of spine
C0178013|ICD9CM|PT|93.15|Mobilization of spine
C0178014|ICD9CM|PT|93.16|Mobilization of other joints
C0178014|ICD9CM|AB|93.16|Other joint mobilization
C0178015|ICD9CM|PT|93.17|Other passive musculoskeletal exercise
C0178015|ICD9CM|AB|93.17|Pass musculosk exer NEC
C0178016|ICD9CM|HT|93.2|Other physical therapy musculoskeletal manipulation
C0178017|ICD9CM|PT|93.24|Training in use of prosthetic or orthotic device
C0178017|ICD9CM|AB|93.24|Prosthet/orthot training
C0178019|ICD9CM|PT|93.27|Stretching of muscle or tendon
C0178019|ICD9CM|AB|93.27|Musc or tend stretching
C0178020|ICD9CM|AB|93.28|Stretching of fascia
C0178020|ICD9CM|PT|93.28|Stretching of fascia
C0178021|ICD9CM|PT|93.29|Other forcible correction of musculoskeletal deformity
C0178021|ICD9CM|AB|93.29|Forcib correct defor NEC
C0178023|ICD9CM|PT|93.31|Assisted exercise in pool
C0178023|ICD9CM|AB|93.31|Assisted pool exercise
C0178024|ICD9CM|AB|93.37|Prenatal training
C0178024|ICD9CM|PT|93.37|Prenatal training
C0178025|ICD9CM|HT|93.4|Skeletal traction and other traction
C0178026|ICD9CM|PT|93.41|Spinal traction using skull device
C0178026|ICD9CM|AB|93.41|Spine tract w skull dev
C0178027|ICD9CM|AB|93.42|Other spinal traction
C0178027|ICD9CM|PT|93.42|Other spinal traction
C0178028|ICD9CM|PT|93.43|Intermittent skeletal traction
C0178028|ICD9CM|AB|93.43|Intermitt skel traction
C0178029|ICD9CM|AB|93.44|Other skeletal traction
C0178029|ICD9CM|PT|93.44|Other skeletal traction
C0178030|ICD9CM|AB|93.45|Thomas' splint traction
C0178030|ICD9CM|PT|93.45|Thomas' splint traction
C0178031|ICD9CM|PT|93.46|Other skin traction of limbs
C0178031|ICD9CM|AB|93.46|Limb skin traction NEC
C0178032|ICD9CM|HT|93.5|Other immobilization, pressure, and attention to wound
C0178032|ICD9CM|PT|93.59|Other immobilization, pressure, and attention to wound
C0178032|ICD9CM|AB|93.59|Immobiliz/wound attn NEC
C0178033|ICD9CM|PT|93.51|Application of plaster jacket
C0178033|ICD9CM|AB|93.51|Plaster jacket applicat
C0178034|ICD9CM|AB|93.52|Neck support application
C0178034|ICD9CM|PT|93.52|Application of neck support
C0178036|ICD9CM|AB|93.55|Dental wiring
C0178036|ICD9CM|PT|93.55|Dental wiring
C0178037|ICD9CM|PT|93.58|Application of pressure trousers
C0178037|ICD9CM|AB|93.58|Pressure trouser applica
C0178039|ICD9CM|PT|93.61|Osteopathic manipulative treatment for general mobilization
C0178039|ICD9CM|AB|93.61|Omt for gen'l mobilizat
C0178040|ICD9CM|PT|93.63|Osteopathic manipulative treatment using low- velocity, high-amplitude forces
C0178040|ICD9CM|PT|93.62|Osteopathic manipulative treatment using high-velocity, low-amplitude forces
C0178040|ICD9CM|AB|93.62|Omt with hi-vel,lo-ampli
C0178040|ICD9CM|AB|93.63|Omt with lo-vel,hi-ampli
C0178044|ICD9CM|PT|93.67|Other specified osteopathic manipulative treatment
C0178044|ICD9CM|AB|93.67|Osteopath manipulat NEC
C0178045|ICD9CM|HT|93.7|Speech and reading rehabilitation and rehabilitation of the blind
C0178046|ICD9CM|PT|93.78|Other rehabilitation for the blind
C0178046|ICD9CM|AB|93.78|Rehab for the blind NEC
C0178047|ICD9CM|HT|93.8|Other rehabilitation therapy
C0178049|ICD9CM|PT|93.96|Other oxygen enrichment
C0178049|ICD9CM|AB|93.96|Oxygen enrichment NEC
C0178051|ICD9CM|PT|93.98|Other control of atmospheric pressure and composition
C0178051|ICD9CM|AB|93.98|Atmos press/compos contr
C0178052|ICD9CM|HT|94.0|Psychologic evaluation and testing
C0178054|ICD9CM|PT|94.09|Psychologic mental status determination, not otherwise specified
C0178054|ICD9CM|AB|94.09|Psychol mental stat NOS
C0178055|ICD9CM|HT|94.1|Psychiatric interviews, consultations, and evaluations
C0178056|ICD9CM|PT|94.11|Psychiatric mental status determination
C0178056|ICD9CM|AB|94.11|Psychiat mental determin
C0178057|ICD9CM|PT|94.12|Routine psychiatric visit, not otherwise specified
C0178057|ICD9CM|AB|94.12|Routine psychiat visit
C0178058|ICD9CM|PT|94.13|Psychiatric commitment evaluation
C0178058|ICD9CM|AB|94.13|Psychia commitment eval
C0178059|ICD9CM|PT|94.19|Other psychiatric interview and evaluation
C0178059|ICD9CM|AB|94.19|Psychia interv/eval NEC
C0178060|ICD9CM|PT|94.25|Other psychiatric drug therapy
C0178060|ICD9CM|AB|94.25|Psychiat drug therap NEC
C0178061|ICD9CM|PT|94.34|Individual therapy for psychosexual dysfunction
C0178061|ICD9CM|AB|94.34|Ind therap psychsex dysf
C0178062|ICD9CM|HT|94.4|Other psychotherapy and counselling
C0178063|ICD9CM|PT|94.41|Group therapy for psychosexual dysfunction
C0178063|ICD9CM|AB|94.41|Grp therap psychsex dysf
C0178066|ICD9CM|HT|94.5|Referral for psychologic rehabilitation
C0178067|ICD9CM|PT|94.51|Referral for psychotherapy
C0178067|ICD9CM|AB|94.51|Referral for psychother
C0178068|ICD9CM|PT|94.52|Referral for psychiatric aftercare
C0178068|ICD9CM|AB|94.52|Referral psych aftercare
C0178071|ICD9CM|PT|94.55|Referral for vocational rehabilitation
C0178071|ICD9CM|AB|94.55|Referral vocation rehab
C0178072|ICD9CM|PT|94.59|Referral for other psychologic rehabilitation
C0178072|ICD9CM|AB|94.59|Referral psych rehab NEC
C0178073|ICD9CM|HT|94.6|Alcohol and drug rehabilitation and detoxification
C0178074|ICD9CM|HT|95.0|General and subjective eye examination
C0178076|ICD9CM|HT|95.1|Examinations of form and structure of eye
C0178078|ICD9CM|PT|95.12|Fluorescein angiography or angioscopy of eye
C0178078|ICD9CM|AB|95.12|Eye fluorescein angiogra
C0178080|ICD9CM|PT|95.16|P32 and other tracer studies of eye
C0178080|ICD9CM|AB|95.16|P32 & eye tracer NEC
C0178081|ICD9CM|HT|95.2|Objective functional tests of eye
C0178085|ICD9CM|PT|95.26|Tonography, provocative tests, and other glaucoma testing
C0178085|ICD9CM|AB|95.26|Glaucoma testing
C0178086|ICD9CM|HT|95.3|Special vision services
C0178087|ICD9CM|PT|95.33|Dispensing of other low vision aids
C0178087|ICD9CM|AB|95.33|Oth lo vision aid dispen
C0178088|ICD9CM|AB|95.34|Ocular prosthetics
C0178088|ICD9CM|PT|95.34|Ocular prosthetics
C0178089|ICD9CM|HT|95.4|Nonoperative procedures related to hearing
C0178090|ICD9CM|PT|95.44|Clinical vestibular function tests
C0178090|ICD9CM|AB|95.44|Clin vestibul funct test
C0178091|ICD9CM|AB|95.45|Rotation tests
C0178091|ICD9CM|PT|95.45|Rotation tests
C0178092|ICD9CM|HT|96.0|Nonoperative intubation of gastrointestinal and respiratory tracts
C0178093|ICD9CM|PT|96.01|Insertion of nasopharyngeal airway
C0178093|ICD9CM|AB|96.01|Insert nasopharyn airway
C0178094|ICD9CM|PT|96.03|Insertion of esophageal obturator airway
C0178094|ICD9CM|AB|96.03|Insert esoph obtu airway
C0178095|ICD9CM|PT|96.05|Other intubation of respiratory tract
C0178095|ICD9CM|AB|96.05|Resp tract intubat NEC
C0178097|ICD9CM|PT|96.07|Insertion of other (naso-)gastric tube
C0178097|ICD9CM|AB|96.07|Insert gastric tube NEC
C0178098|ICD9CM|PT|96.08|Insertion of (naso-)intestinal tube
C0178098|ICD9CM|AB|96.08|Insert intestinal tube
C0178099|ICD9CM|PT|96.09|Insertion of rectal tube
C0178099|ICD9CM|AB|96.09|Insert rectal tube
C0178100|ICD9CM|HT|96.1|Other nonoperative insertion
C0178102|ICD9CM|AB|96.16|Other vaginal dilation
C0178102|ICD9CM|PT|96.16|Other vaginal dilation
C0178104|ICD9CM|PT|96.18|Insertion of other vaginal pessary
C0178104|ICD9CM|AB|96.18|Oth vagin pessary insert
C0178105|ICD9CM|HT|96.2|Nonoperative dilation and manipulation
C0178106|ICD9CM|PT|96.23|Dilation of anal sphincter
C0178106|ICD9CM|AB|96.23|Dilation anal sphincter
C0178108|ICD9CM|HT|96.3|Nonoperative alimentary tract irrigation, cleaning, and local instillation
C0178109|ICD9CM|PT|96.34|Other irrigation of (naso-)gastric tube
C0178109|ICD9CM|AB|96.34|Gastric tube irrigat NEC
C0178111|ICD9CM|HT|96.4|Nonoperative irrigation, cleaning, and local instillation of other digestive and genitourinary organs
C0178112|ICD9CM|PT|96.41|Irrigation of cholecystostomy and other biliary tube
C0178112|ICD9CM|AB|96.41|Biliary tube irrigation
C0178115|ICD9CM|PT|96.48|Irrigation of other indwelling urinary catheter
C0178115|ICD9CM|AB|96.48|Indwell cath irrig NEC
C0178116|ICD9CM|PT|96.49|Other genitourinary instillation
C0178116|ICD9CM|AB|96.49|Other gu instillation
C0178117|ICD9CM|HT|96.5|Other nonoperative irrigation and cleaning
C0178118|ICD9CM|AB|96.55|Tracheostomy toilette
C0178118|ICD9CM|PT|96.55|Tracheostomy toilette
C0178119|ICD9CM|PT|96.56|Other lavage of bronchus and trachea
C0178119|ICD9CM|AB|96.56|Bronch/trach lavage NEC
C0178121|ICD9CM|PT|96.59|Other irrigation of wound
C0178121|ICD9CM|AB|96.59|Wound irrigation NEC
C0178126|ICD9CM|HT|97.0|Nonoperative replacement of gastrointestinal appliance
C0178127|ICD9CM|PT|97.01|Replacement of (naso-)gastric or esophagostomy tube
C0178127|ICD9CM|AB|97.01|Replace gast/esoph tube
C0178128|ICD9CM|PT|97.05|Replacement of stent (tube) in biliary or pancreatic duct
C0178128|ICD9CM|AB|97.05|Repl stent in bile duct
C0178129|ICD9CM|HT|97.1|Nonoperative replacement of musculoskeletal and integumentary system appliance
C0178130|ICD9CM|PT|97.11|Replacement of cast on upper limb
C0178130|ICD9CM|AB|97.11|Replace upper limb cast
C0178131|ICD9CM|PT|97.12|Replacement of cast on lower limb
C0178131|ICD9CM|AB|97.12|Replace lower limb cast
C0178132|ICD9CM|PT|97.13|Replacement of other cast
C0178132|ICD9CM|AB|97.13|Replace cast NEC
C0178133|ICD9CM|PT|97.14|Replacement of other device for musculoskeletal immobilization
C0178133|ICD9CM|AB|97.14|Replac m/s immob dev NEC
C0178134|ICD9CM|PT|97.15|Replacement of wound catheter
C0178134|ICD9CM|AB|97.15|Replace wound catheter
C0178135|ICD9CM|PT|97.16|Replacement of wound packing or drain
C0178135|ICD9CM|AB|97.16|Replace wound pack/drain
C0178136|ICD9CM|PT|97.29|Other nonoperative replacements
C0178136|ICD9CM|HT|97.2|Other nonoperative replacement
C0178136|ICD9CM|AB|97.29|Non-op replacement NEC
C0178137|ICD9CM|PT|97.22|Replacement of dental packing
C0178137|ICD9CM|AB|97.22|Replace dental packing
C0178139|ICD9CM|PT|97.24|Replacement and refitting of vaginal diaphragm
C0178139|ICD9CM|AB|97.24|Replace vag diaphragm
C0178140|ICD9CM|PT|97.25|Replacement of other vaginal pessary
C0178140|ICD9CM|AB|97.25|Replace vaginal pessary
C0178141|ICD9CM|PT|97.26|Replacement of vaginal or vulvar packing or drain
C0178141|ICD9CM|AB|97.26|Replace vag/vulv packing
C0178143|ICD9CM|HT|97.3|Nonoperative removal of therapeutic device from head and neck
C0178144|ICD9CM|PT|97.33|Removal of dental wiring
C0178144|ICD9CM|AB|97.33|Remove dental wiring
C0178145|ICD9CM|PT|97.34|Removal of dental packing
C0178145|ICD9CM|AB|97.34|Remove dental packing
C0178146|ICD9CM|PT|97.35|Removal of dental prosthesis
C0178146|ICD9CM|AB|97.35|Remove dental prosthesis
C0178147|ICD9CM|PT|97.36|Removal of other external mandibular fixation device
C0178147|ICD9CM|AB|97.36|Remove ext mand fix dev
C0178148|ICD9CM|PT|97.37|Removal of tracheostomy tube
C0178148|ICD9CM|AB|97.37|Remove tracheostomy tube
C0178149|ICD9CM|PT|97.38|Removal of sutures from head and neck
C0178149|ICD9CM|AB|97.38|Remove head/neck sutures
C0178150|ICD9CM|PT|97.39|Removal of other therapeutic device from head and neck
C0178150|ICD9CM|AB|97.39|Remove head/neck dev NEC
C0178151|ICD9CM|HT|97.4|Nonoperative removal of therapeutic device from thorax
C0178152|ICD9CM|PT|97.41|Removal of thoracotomy tube or pleural cavity drain
C0178152|ICD9CM|AB|97.41|Remov thoracotomy tube
C0178153|ICD9CM|PT|97.43|Removal of sutures from thorax
C0178153|ICD9CM|AB|97.43|Remov thorax sutures
C0178154|ICD9CM|PT|97.49|Removal of other device from thorax
C0178154|ICD9CM|AB|97.49|Remov thor ther dev NEC
C0178155|ICD9CM|HT|97.5|Nonoperative removal of therapeutic device from digestive system
C0178156|ICD9CM|PT|97.53|Removal of tube from large intestine or appendix
C0178156|ICD9CM|AB|97.53|Remov large bowel tube
C0178157|ICD9CM|PT|97.55|Removal of T-tube, other bile duct tube, or liver tube
C0178157|ICD9CM|AB|97.55|Remov biliary/liver tube
C0178158|ICD9CM|PT|97.56|Removal of pancreatic tube or drain
C0178158|ICD9CM|AB|97.56|Remov pancreatic tube
C0178159|ICD9CM|PT|97.59|Removal of other device from digestive system
C0178159|ICD9CM|AB|97.59|Remov other GI device
C0178160|ICD9CM|HT|97.6|Nonoperative removal of therapeutic device from urinary system
C0178161|ICD9CM|PT|97.64|Removal of other urinary drainage device
C0178161|ICD9CM|AB|97.64|Remov urin drainage NEC
C0178162|ICD9CM|PT|97.69|Removal of other device from urinary system
C0178162|ICD9CM|AB|97.69|Remov other urin device
C0178163|ICD9CM|HT|97.7|Nonoperative removal of therapeutic device from genital system
C0178165|ICD9CM|PT|97.74|Removal of other vaginal pessary
C0178165|ICD9CM|AB|97.74|Removal oth vag pessary
C0178166|ICD9CM|PT|97.75|Removal of vaginal or vulvar packing
C0178166|ICD9CM|AB|97.75|Remov vag/vulv packing
C0178167|ICD9CM|PT|97.79|Removal of other device from genital tract
C0178167|ICD9CM|AB|97.79|Remov other genit device
C0178168|ICD9CM|HT|97.8|Other nonoperative removal of therapeutic device
C0178169|ICD9CM|PT|97.83|Removal of abdominal wall sutures
C0178169|ICD9CM|AB|97.83|Remov abdom wall suture
C0178172|ICD9CM|PT|97.86|Removal of other device from abdomen
C0178172|ICD9CM|AB|97.86|Remov abdomen device NEC
C0178173|ICD9CM|PT|97.87|Removal of other device from trunk
C0178173|ICD9CM|AB|97.87|Remov trunk device NEC
C0178174|ICD9CM|PT|97.89|Removal of other therapeutic device
C0178174|ICD9CM|AB|97.89|Remov therapeut dev NEC
C0178175|ICD9CM|HT|98.0|Removal of intraluminal foreign body from digestive system without incision
C0178177|ICD9CM|PT|98.03|Removal of intraluminal foreign body from stomach and small intestine without incision
C0178177|ICD9CM|AB|98.03|Remov intralum gastr FB
C0178178|ICD9CM|PT|98.05|Removal of intraluminal foreign body from rectum and anus without incision
C0178178|ICD9CM|AB|98.05|Remov intralum rect FB
C0178179|ICD9CM|HT|98.1|Removal of intraluminal foreign body from other sites without incision
C0178180|ICD9CM|PT|98.14|Removal of intraluminal foreign body from larynx without incision
C0178180|ICD9CM|AB|98.14|Remov intralum laryn FB
C0178181|ICD9CM|PT|98.15|Removal of intraluminal foreign body from trachea and bronchus without incision
C0178181|ICD9CM|AB|98.15|Remov intralum trach FB
C0178182|ICD9CM|PT|98.19|Removal of intraluminal foreign body from urethra without incision
C0178182|ICD9CM|AB|98.19|Remove intralum ureth FB
C0178183|ICD9CM|HT|98.2|Removal of other foreign body without incision
C0178184|ICD9CM|PT|98.22|Removal of other foreign body without incision from head and neck
C0178184|ICD9CM|AB|98.22|Removal head/neck FB
C0178185|ICD9CM|PT|98.23|Removal of foreign body from vulva without incision
C0178185|ICD9CM|AB|98.23|Removal vulvar FB
C0178186|ICD9CM|PT|98.24|Removal of foreign body from scrotum or penis without incision
C0178186|ICD9CM|AB|98.24|Removal scrotal/penis FB
C0178187|ICD9CM|PT|98.25|Removal of other foreign body without incision from trunk except scrotum, penis, or vulva
C0178187|ICD9CM|AB|98.25|Removal trunk FB NEC
C0178189|ICD9CM|PT|98.51|Extracorporeal shockwave lithotripsy [ESWL] of the kidney, ureter and/or bladder
C0178189|ICD9CM|AB|98.51|Eswl kid/ureter/bladder
C0178190|ICD9CM|PT|98.52|Extracorporeal shockwave lithotripsy [ESWL] of the gallbladder and/or bile duct
C0178190|ICD9CM|AB|98.52|Eswl gb/bile duct
C0178192|ICD9CM|PT|99.04|Transfusion of packed cells
C0178192|ICD9CM|AB|99.04|Packed cell transfusion
C0178193|ICD9CM|PT|99.09|Transfusion of other substance
C0178193|ICD9CM|AB|99.09|Transfusion NEC
C0178194|ICD9CM|HT|99.1|Injection or infusion of therapeutic or prophylactic substance
C0178196|ICD9CM|PT|99.18|Injection or infusion of electrolytes
C0178196|ICD9CM|AB|99.18|Inject/infuse electrolyt
C0178197|ICD9CM|HT|99.2|Injection or infusion of other therapeutic or prophylactic substance
C0178197|ICD9CM|PT|99.29|Injection or infusion of other therapeutic or prophylactic substance
C0178197|ICD9CM|AB|99.29|Inject/infuse NEC
C0178198|ICD9CM|PT|99.22|Injection of other anti-infective
C0178198|ICD9CM|AB|99.22|Inject anti-infect NEC
C0178199|ICD9CM|PT|99.24|Injection of other hormone
C0178199|ICD9CM|AB|99.24|Inject hormone NEC
C0178200|ICD9CM|PT|99.25|Injection or infusion of cancer chemotherapeutic substance
C0178200|ICD9CM|AB|99.25|Inject ca chemother NEC
C0178201|ICD9CM|HT|99.3|Prophylactic vaccination and inoculation against certain bacterial diseases
C0178203|ICD9CM|PT|99.32|Vaccination against typhoid and paratyphoid fever
C0178203|ICD9CM|AB|99.32|Typhoid/paratyphoid vacc
C0178209|ICD9CM|HT|99.4|Prophylactic vaccination and inoculation against certain viral diseases
C0178221|ICD9CM|PT|99.54|Prophylactic vaccination against other arthropod-borne viral diseases
C0178221|ICD9CM|AB|99.54|Arbovirus vaccinat NEC
C0178222|ICD9CM|PT|99.58|Administration of other antitoxins
C0178222|ICD9CM|AB|99.58|Antitoxin administra NEC
C0178224|ICD9CM|PT|99.69|Other conversion of cardiac rhythm
C0178224|ICD9CM|AB|99.69|Cardiac rhythm conv NEC
C0178229|ICD9CM|HT|99.8|Miscellaneous physical procedures
C0178230|ICD9CM|PT|99.86|Non-invasive placement of bone growth stimulator
C0178230|ICD9CM|AB|99.86|Non-invasive bone stimul
C0178234|ICD9CM|PT|99.96|Collection of sperm for artificial insemination
C0178234|ICD9CM|AB|99.96|Sperm collection
C0178235|ICD9CM|PT|99.97|Fitting of denture
C0178235|ICD9CM|AB|99.97|Denture fitting
C0178236|ICD9CM|PT|99.98|Extraction of milk from lactating breast
C0178236|ICD9CM|AB|99.98|Milk extraction
C0178237|ICD9CM|HT|001-999.99|DISEASES AND INJURIES
C0178238|ICD9CM|HT|001-009.99|INTESTINAL INFECTIOUS DISEASES
C0178242|ICD9CM|HT|080-088.99|RICKETTSIOSES AND OTHER ARTHROPOD-BORNE DISEASES
C0178243|ICD9CM|HT|090-099.99|SYPHILIS AND OTHER VENEREAL DISEASES
C0178244|ICD9CM|HT|100-104.99|OTHER SPIROCHETAL DISEASES
C0178247|ICD9CM|HT|140-149.99|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY, AND PHARYNX
C0178249|ICD9CM|HT|160-165.99|MALIGNANT NEOPLASM OF RESPIRATORY AND INTRATHORACIC ORGANS
C0178250|ICD9CM|HT|170-176.99|MALIGNANT NEOPLASM OF BONE, CONNECTIVE TISSUE, SKIN, AND BREAST
C0178251|ICD9CM|HT|179-189.99|MALIGNANT NEOPLASM OF GENITOURINARY ORGANS
C0178257|ICD9CM|HT|249-259.99|DISEASES OF OTHER ENDOCRINE GLANDS
C0178259|ICD9CM|HT|270-279.99|OTHER METABOLIC AND IMMUNITY DISORDERS
C0178264|ICD9CM|HT|320-326.99|INFLAMMATORY DISEASES OF THE CENTRAL NERVOUS SYSTEM
C0178266|ICD9CM|HT|340-349.99|OTHER DISORDERS OF THE CENTRAL NERVOUS SYSTEM
C0178269|ICD9CM|HT|380-389.99|DISEASES OF THE EAR AND MASTOID PROCESS
C0178272|ICD9CM|PT|417.9|Unspecified disease of pulmonary circulation
C0178272|ICD9CM|HT|415-417.99|DISEASES OF PULMONARY CIRCULATION
C0178272|ICD9CM|AB|417.9|Pulmon circulat dis NOS
C0178273|ICD9CM|HT|420-429.99|OTHER FORMS OF HEART DISEASE
C0178274|ICD9CM|HT|440-449.99|DISEASES OF ARTERIES, ARTERIOLES, AND CAPILLARIES
C0178278|ICD9CM|HT|490-496.99|CHRONIC OBSTRUCTIVE PULMONARY DISEASE AND ALLIED CONDITIONS
C0178279|ICD9CM|HT|500-508.99|PNEUMOCONIOSES AND OTHER LUNG DISEASES DUE TO EXTERNAL AGENTS
C0178281|ICD9CM|HT|530-539.99|DISEASES OF ESOPHAGUS, STOMACH, AND DUODENUM
C0178282|ICD9CM|HT|550-553.99|HERNIA OF ABDOMINAL CAVITY
C0178283|ICD9CM|HT|555-558.99|NONINFECTIOUS ENTERITIS AND COLITIS
C0178284|ICD9CM|HT|560-569.99|OTHER DISEASES OF INTESTINES AND PERITONEUM
C0178285|ICD9CM|HT|570-579.99|OTHER DISEASES OF DIGESTIVE SYSTEM
C0178287|ICD9CM|HT|580-589.99|NEPHRITIS, NEPHROTIC SYNDROME, AND NEPHROSIS
C0178288|ICD9CM|HT|590-599.99|OTHER DISEASES OF URINARY SYSTEM
C0178291|ICD9CM|HT|617-629.99|OTHER DISORDERS OF FEMALE GENITAL TRACT
C0178292|ICD9CM|HT|630-679.99|COMPLICATIONS OF PREGNANCY, CHILDBIRTH, AND THE PUERPERIUM
C0178293|ICD9CM|HT|630-633.99|ECTOPIC AND MOLAR PREGNANCY
C0178294|ICD9CM|HT|634-639.99|OTHER PREGNANCY WITH ABORTIVE OUTCOME
C0178295|ICD9CM|HT|640-649.99|COMPLICATIONS MAINLY RELATED TO PREGNANCY
C0178296|ICD9CM|HT|650-659.99|NORMAL DELIVERY, AND OTHER INDICATIONS FOR CARE IN PREGNANCY, LABOR, AND DELIVERY
C0178297|ICD9CM|HT|660-669.99|COMPLICATIONS OCCURRING MAINLY IN THE COURSE OF LABOR AND DELIVERY
C0178298|ICD9CM|PT|709.9|Unspecified disorder of skin and subcutaneous tissue
C0178298|ICD9CM|AB|709.9|Skin disorder NOS
C0178298|ICD9CM|HT|680-709.99|DISEASES OF THE SKIN AND SUBCUTANEOUS TISSUE
C0178300|ICD9CM|HT|690-698.99|OTHER INFLAMMATORY CONDITIONS OF SKIN AND SUBCUTANEOUS TISSUE
C0178301|ICD9CM|HT|700-709.99|OTHER DISEASES OF SKIN AND SUBCUTANEOUS TISSUE
C0178301|ICD9CM|HT|709|Other disorders of skin and subcutaneous tissue
C0178303|ICD9CM|HT|710-719.99|ARTHROPATHIES AND RELATED DISORDERS
C0178305|ICD9CM|HT|725-729.99|RHEUMATISM, EXCLUDING THE BACK
C0178306|ICD9CM|HT|730-739.99|OSTEOPATHIES, CHONDROPATHIES, AND ACQUIRED MUSCULOSKELETAL DEFORMITIES
C0178307|ICD9CM|HT|760-779.99|CERTAIN CONDITIONS ORIGINATING IN THE PERINATAL PERIOD
C0178308|ICD9CM|HT|760-763.99|MATERNAL CAUSES OF PERINATAL MORBIDITY AND MORTALITY
C0178309|ICD9CM|HT|764-779.99|OTHER CONDITIONS ORIGINATING IN THE PERINATAL PERIOD
C0178310|ICD9CM|HT|780-799.99|SYMPTOMS, SIGNS, AND ILL-DEFINED CONDITIONS
C0178314|ICD9CM|HT|800-999.99|INJURY AND POISONING
C0178315|ICD9CM|HT|805-809.99|FRACTURE OF NECK AND TRUNK
C0178316|ICD9CM|HT|810-819.99|FRACTURE OF UPPER LIMB
C0178319|ICD9CM|HT|850-854.99|INTRACRANIAL INJURY, EXCLUDING THOSE WITH SKULL FRACTURE
C0178321|ICD9CM|HT|870-879.99|OPEN WOUND OF HEAD, NECK, AND TRUNK
C0178322|ICD9CM|HT|880-887.99|OPEN WOUND OF UPPER LIMB
C0178323|ICD9CM|HT|890-897.99|OPEN WOUND OF LOWER LIMB
C0178324|ICD9CM|PT|904.9|Injury to blood vessels of unspecified site
C0178324|ICD9CM|HT|900-904.99|INJURY TO BLOOD VESSELS
C0178324|ICD9CM|AB|904.9|Blood vessel injury NOS
C0178325|ICD9CM|HT|905-909.99|LATE EFFECTS OF INJURIES, POISONINGS, TOXIC EFFECTS, AND OTHER EXTERNAL CAUSES
C0178327|ICD9CM|HT|920-924.99|CONTUSION WITH INTACT SKIN SURFACE
C0178329|ICD9CM|HT|930-939.99|EFFECTS OF FOREIGN BODY ENTERING THROUGH ORIFICE
C0178330|ICD9CM|HT|950-957.99|INJURY TO NERVES AND SPINAL CORD
C0178331|ICD9CM|HT|958-959.99|CERTAIN TRAUMATIC COMPLICATIONS AND UNSPECIFIED INJURIES
C0178332|ICD9CM|HT|960-979.99|POISONING BY DRUGS, MEDICINAL AND BIOLOGICAL SUBSTANCES
C0178337|ICD9CM|HT|V01-V06.99|PERSONS WITH POTENTIAL HEALTH HAZARDS RELATED TO COMMUNICABLE DISEASES
C0178338|ICD9CM|HT|V10-V19.99|PERSONS WITH POTENTIAL HEALTH HAZARDS RELATED TO PERSONAL AND FAMILY HISTORY
C0178339|ICD9CM|HT|V20-V29.99|PERSONS ENCOUNTERING HEALTH SERVICES IN CIRCUMSTANCES RELATED TO REPRODUCTION AND DEVELOPMENT
C0178340|ICD9CM|HT|V30-V39.99|LIVEBORN INFANTS ACCORDING TO TYPE OF BIRTH
C0178341|ICD9CM|HT|V40-V49.99|PERSONS WITH A CONDITION INFLUENCING THEIR HEALTH STATUS
C0178342|ICD9CM|HT|V50-V59.99|PERSONS ENCOUNTERING HEALTH SERVICES FOR SPECIFIC PROCEDURES AND AFTERCARE
C0178343|ICD9CM|HT|V60-V69.99|PERSONS ENCOUNTERING HEALTH SERVICES IN OTHER CIRCUMSTANCES
C0178348|ICD9CM|HT|E820-E825.9|MOTOR VEHICLE NONTRAFFIC ACCIDENTS
C0178350|ICD9CM|HT|E840-E845.9|AIR AND SPACE TRANSPORT ACCIDENTS
C0178352|ICD9CM|HT|E850-E858.9|ACCIDENTAL POISONING BY DRUGS, MEDICINAL SUBSTANCES, AND BIOLOGICALS
C0178353|ICD9CM|HT|E860-E869.9|ACCIDENTAL POISONING BY OTHER SOLID AND LIQUID SUBSTANCES, GASES, AND VAPORS
C0178355|ICD9CM|HT|E878-E879.9|SURGICAL AND MEDICAL PROCEDURES AS THE CAUSE OF ABNORMAL REACTION OF PATIENT OR LATER COMPLICATION, WITHOUT MENTION OF MISADVENTURE AT THE TIME OF PROCEDURE
C0178356|ICD9CM|HT|E890-E899.9|ACCIDENTS CAUSED BY FIRE AND FLAMES
C0178357|ICD9CM|HT|E900-E909.9|ACCIDENTS DUE TO NATURAL AND ENVIRONMENTAL FACTORS
C0178358|ICD9CM|HT|E910-E915.9|ACCIDENTS CAUSED BY SUBMERSION, SUFFOCATION, AND FOREIGN BODIES
C0178359|ICD9CM|HT|E930-E949.9|DRUGS, MEDICINAL AND BIOLOGICAL SUBSTANCES CAUSING ADVERSE EFFECTS IN THERAPEUTIC USE
C0178360|ICD9CM|HT|E950-E959.9|SUICIDE AND SELF-INFLICTED INJURY
C0178361|ICD9CM|HT|E960-E969.9|HOMICIDE AND INJURY PURPOSELY INFLICTED BY OTHER PERSONS
C0178362|ICD9CM|HT|E970-E978.9|LEGAL INTERVENTION
C0178363|ICD9CM|HT|E980-E989.9|INJURY UNDETERMINED WHETHER ACCIDENTALLY OR PURPOSELY INFLICTED
C0178364|ICD9CM|HT|E990-E999.9|INJURY RESULTING FROM OPERATIONS OF WAR
C0178369|ICD9CM|HT|21-29.99|OPERATIONS ON THE NOSE, MOUTH, AND PHARYNX
C0178372|ICD9CM|HT|40-41.99|OPERATIONS ON THE HEMIC AND LYMPHATIC SYSTEM
C0178380|ICD9CM|HT|87-99.99|MISCELLANEOUS DIAGNOSTIC AND THERAPEUTIC PROCEDURES
C0178415|ICD9CM|PT|790.93|Elevated prostate specific antigen [PSA]
C0178415|ICD9CM|AB|790.93|Elvtd prstate spcf antgn
C0178879|ICD9CM|HT|599.6|Urinary obstruction
C0178879|ICD9CM|AB|599.60|Urinary obstruction NOS
C0178879|ICD9CM|PT|599.60|Urinary obstruction, unspecified
C0184567|ICD9CM|HT|338.1|Acute pain
C0184661|ICD9CM|HT|00-99.99|PROCEDURES
C0184748|ICD9CM|PT|94.53|Referral for alcoholism rehabilitation
C0184748|ICD9CM|AB|94.53|Referral alcohol rehab
C0184749|ICD9CM|PT|94.54|Referral for drug addiction rehabilitation
C0184749|ICD9CM|AB|94.54|Referral for drug rehab
C0184968|ICD9CM|PT|86.93|Insertion of tissue expander
C0184968|ICD9CM|AB|86.93|Insert tissue expander
C0184989|ICD9CM|PT|86.83|Size reduction plastic operation
C0184989|ICD9CM|AB|86.83|Size reduct plastic op
C0185130|ICD9CM|HT|76-84.99|OPERATIONS ON THE MUSCULOSKELETAL SYSTEM
C0185150|ICD9CM|HT|79.9|Unspecified operation on bone injury
C0185153|ICD9CM|HT|77.2|Wedge osteotomy
C0185153|ICD9CM|AB|77.20|Wedge osteotomy NOS
C0185153|ICD9CM|PT|77.20|Wedge osteotomy, unspecified site
C0185171|ICD9CM|PT|83.01|Exploration of tendon sheath
C0185171|ICD9CM|AB|83.01|Tendon sheath explorat
C0185181|ICD9CM|AB|83.02|Myotomy
C0185181|ICD9CM|PT|83.02|Myotomy
C0185188|ICD9CM|AB|83.14|Fasciotomy
C0185188|ICD9CM|PT|83.14|Fasciotomy
C0185195|ICD9CM|AB|83.03|Bursotomy
C0185195|ICD9CM|PT|83.03|Bursotomy
C0185216|ICD9CM|HT|77.0|Sequestrectomy
C0185216|ICD9CM|AB|77.00|Sequestrectomy NOS
C0185216|ICD9CM|PT|77.00|Sequestrectomy, unspecified site
C0185223|ICD9CM|HT|77.7|Excision of bone for graft
C0185234|ICD9CM|HT|77.9|Total ostectomy
C0185249|ICD9CM|HT|80.3|Biopsy of joint structure
C0185259|ICD9CM|PT|83.41|Excision of tendon for graft
C0185259|ICD9CM|AB|83.41|Tendon excision for grft
C0185264|ICD9CM|PT|83.31|Excision of lesion of tendon sheath
C0185264|ICD9CM|AB|83.31|Excis les tendon sheath
C0185287|ICD9CM|PT|83.32|Excision of lesion of muscle
C0185287|ICD9CM|AB|83.32|Excis lesion of muscle
C0185298|ICD9CM|AB|83.5|Bursectomy
C0185298|ICD9CM|PT|83.5|Bursectomy
C0185304|ICD9CM|HT|80.7|Synovectomy
C0185304|ICD9CM|PT|80.70|Synovectomy, unspecified site
C0185304|ICD9CM|AB|80.70|Synovectomy-site NOS
C0185314|ICD9CM|HT|78.6|Removal of implanted device from bone
C0185320|ICD9CM|HT|78.9|Insertion of bone growth stimulator
C0185320|ICD9CM|PT|78.90|Insertion of bone growth stimulator, unspecified site
C0185320|ICD9CM|AB|78.90|Insert bone stimul NOS
C0185333|ICD9CM|PT|83.96|Injection of therapeutic substance into bursa
C0185333|ICD9CM|AB|83.96|Injection into bursa
C0185336|ICD9CM|PT|83.97|Injection of therapeutic substance into tendon
C0185336|ICD9CM|AB|83.97|Injection into tendon
C0185349|ICD9CM|HT|80.0|Arthrotomy for removal of prosthesis
C0185372|ICD9CM|HT|78.5|Internal fixation of bone without fracture reduction
C0185379|ICD9CM|AB|82.83|Repair of macrodactyly
C0185379|ICD9CM|PT|82.83|Repair of macrodactyly
C0185380|ICD9CM|HT|79.5|Open reduction of separated epiphysis
C0185392|ICD9CM|HT|79.8|Open reduction of dislocation
C0185398|ICD9CM|PT|83.73|Reattachment of tendon
C0185398|ICD9CM|AB|83.73|Tendon reattachment
C0185415|ICD9CM|PT|83.74|Reattachment of muscle
C0185415|ICD9CM|AB|83.74|Muscle reattachment
C0185432|ICD9CM|PT|84.3|Revision of amputation stump
C0185432|ICD9CM|AB|84.3|Amputation stump revis
C0185436|ICD9CM|PT|84.93|Separation of unequal conjoined twins
C0185436|ICD9CM|AB|84.93|Separat unequl join twin
C0185439|ICD9CM|PT|83.62|Delayed suture of tendon
C0185439|ICD9CM|AB|83.62|Delayed tendon suture
C0185440|ICD9CM|PT|83.61|Suture of tendon sheath
C0185440|ICD9CM|AB|83.61|Tendon sheath suture
C0185451|ICD9CM|HT|78.7|Osteoclasis
C0185451|ICD9CM|AB|78.70|Osteoclasis NOS
C0185451|ICD9CM|PT|78.70|Osteoclasis, unspecified site
C0185465|ICD9CM|PT|83.71|Advancement of tendon
C0185465|ICD9CM|AB|83.71|Tendon advancement
C0185466|ICD9CM|PT|83.72|Recession of tendon
C0185466|ICD9CM|AB|83.72|Tendon recession
C0185497|ICD9CM|HT|79.0|Closed reduction of fracture without internal fixation
C0185497|ICD9CM|PT|79.00|Closed reduction of fracture without internal fixation, unspecified site
C0185497|ICD9CM|AB|79.00|Closed fx reduction NOS
C0185498|ICD9CM|HT|79.1|Closed reduction of fracture with internal fixation
C0185498|ICD9CM|PT|79.10|Closed reduction of fracture with internal fixation, unspecified site
C0185498|ICD9CM|AB|79.10|Cl fx reduc-int fix NOS
C0185499|ICD9CM|HT|79.4|Closed reduction of separated epiphysis
C0185500|ICD9CM|HT|79.7|Closed reduction of dislocation
C0185505|ICD9CM|HT|84.4|Implantation or fitting of prosthetic limb device
C0185505|ICD9CM|PT|84.40|Implantation or fitting of prosthetic limb device, not otherwise specified
C0185505|ICD9CM|AB|84.40|Implnt/fit pros limb NOS
C0185558|ICD9CM|HT|76.3|Partial ostectomy of facial bone
C0185565|ICD9CM|PT|76.01|Sequestrectomy of facial bone
C0185565|ICD9CM|AB|76.01|Facial bone sequestrect
C0185568|ICD9CM|AB|76.31|Partial mandibulectomy
C0185568|ICD9CM|PT|76.31|Partial mandibulectomy
C0185584|ICD9CM|PT|76.92|Insertion of synthetic implant in facial bone
C0185584|ICD9CM|AB|76.92|Syn implant to face bone
C0185585|ICD9CM|PT|76.97|Removal of internal fixation device from facial bone
C0185585|ICD9CM|AB|76.97|Remove int fix face bone
C0185589|ICD9CM|PT|76.96|Injection of therapeutic substance into temporomandibular joint
C0185589|ICD9CM|AB|76.96|Injec therap sbst tm jnt
C0185594|ICD9CM|HT|76.7|Reduction of facial fracture
C0185594|ICD9CM|PT|76.70|Reduction of facial fracture, not otherwise specified
C0185594|ICD9CM|AB|76.70|Reduction facial fx NOS
C0185605|ICD9CM|PT|86.81|Repair for facial weakness
C0185605|ICD9CM|AB|86.81|Repair facial weakness
C0185649|ICD9CM|PT|76.66|Total osteoplasty [osteotomy] of maxilla
C0185649|ICD9CM|AB|76.66|Tot osteoplasty maxilla
C0185650|ICD9CM|PT|76.65|Segmental osteoplasty [osteotomy] of maxilla
C0185650|ICD9CM|AB|76.65|Seg osteoplasty maxilla
C0185664|ICD9CM|PT|76.74|Open reduction of maxillary fracture
C0185664|ICD9CM|AB|76.74|Open reduct maxillary fx
C0185666|ICD9CM|PT|76.72|Open reduction of malar and zygomatic fracture
C0185666|ICD9CM|AB|76.72|Opn reduct malar/zygo fx
C0185675|ICD9CM|PT|76.41|Total mandibulectomy with synchronous reconstruction
C0185675|ICD9CM|AB|76.41|Tot mandibulec w reconst
C0185680|ICD9CM|PT|76.76|Open reduction of mandibular fracture
C0185680|ICD9CM|AB|76.76|Open reduct mandible fx
C0185688|ICD9CM|PT|76.61|Closed osteoplasty [osteotomy] of mandibular ramus
C0185688|ICD9CM|AB|76.61|Cl osteoplasty mand rami
C0185689|ICD9CM|PT|76.63|Osteoplasty [osteotomy] of body of mandible
C0185689|ICD9CM|AB|76.63|Osteoplasty mandible bdy
C0185690|ICD9CM|PT|76.62|Open osteoplasty [osteotomy] of mandibular ramus
C0185690|ICD9CM|AB|76.62|Open osteoplas mand rami
C0185695|ICD9CM|AB|76.67|Reduction genioplasty
C0185695|ICD9CM|PT|76.67|Reduction genioplasty
C0185696|ICD9CM|AB|76.68|Augmentation genioplasty
C0185696|ICD9CM|PT|76.68|Augmentation genioplasty
C0185702|ICD9CM|PT|76.77|Open reduction of alveolar fracture
C0185702|ICD9CM|AB|76.77|Open reduct alveolar fx
C0185711|ICD9CM|PT|76.94|Open reduction of temporomandibular dislocation
C0185711|ICD9CM|AB|76.94|Open reduct tm dislocat
C0185716|ICD9CM|PT|76.91|Bone graft to facial bone
C0185716|ICD9CM|AB|76.91|Bone graft to face bone
C0185737|ICD9CM|PT|76.93|Closed reduction of temporomandibular dislocation
C0185737|ICD9CM|AB|76.93|Clos reduct tm dislocat
C0185741|ICD9CM|PT|76.75|Closed reduction of mandibular fracture
C0185741|ICD9CM|AB|76.75|Cl reduct mandible fx
C0185760|ICD9CM|PT|76.71|Closed reduction of malar and zygomatic fracture
C0185760|ICD9CM|AB|76.71|Cl reduct malar/zygo fx
C0185762|ICD9CM|PT|76.73|Closed reduction of maxillary fracture
C0185762|ICD9CM|AB|76.73|Cl reduct maxillary fx
C0185824|ICD9CM|AB|84.09|Forequarter amputation
C0185824|ICD9CM|PT|84.09|Interthoracoscapular amputation
C0185912|ICD9CM|PT|03.53|Repair of vertebral fracture
C0185912|ICD9CM|AB|03.53|Vertebral fx repair
C0185990|ICD9CM|HT|81.3|Refusion of spine
C0185990|ICD9CM|PT|81.30|Refusion of spine, not otherwise specified
C0185990|ICD9CM|AB|81.30|Spinal refusion NOS
C0186005|ICD9CM|PT|81.01|Atlas-axis spinal fusion
C0186005|ICD9CM|AB|81.01|Atlas-axis fusion
C0186153|ICD9CM|PT|80.75|Synovectomy, hip
C0186153|ICD9CM|AB|80.75|Hip synovectomy
C0186155|ICD9CM|AB|84.18|Disarticulation of hip
C0186155|ICD9CM|PT|84.18|Disarticulation of hip
C0186190|ICD9CM|PT|80.25|Arthroscopy, hip
C0186190|ICD9CM|AB|80.25|Hip arthroscopy
C0186196|ICD9CM|AB|81.52|Partial hip replacement
C0186196|ICD9CM|PT|81.52|Partial hip replacement
C0186225|ICD9CM|AB|81.21|Arthrodesis of hip
C0186225|ICD9CM|PT|81.21|Arthrodesis of hip
C0186231|ICD9CM|PT|79.85|Open reduction of dislocation of hip
C0186231|ICD9CM|AB|79.85|Open reduc-hip dislocat
C0186325|ICD9CM|PT|78.82|Diagnostic procedures on bone, not elsewhere classified, humerus
C0186325|ICD9CM|AB|78.82|Oth dx proced-humerus
C0186326|ICD9CM|PT|79.91|Unspecified operation on bone injury, humerus
C0186326|ICD9CM|AB|79.91|Humerus injury op NOS
C0186329|ICD9CM|PT|78.83|Diagnostic procedures on bone, not elsewhere classified, radius and ulna
C0186329|ICD9CM|AB|78.83|Oth dx proc-radius/ulna
C0186399|ICD9CM|HT|84.0|Amputation of upper limb
C0186399|ICD9CM|PT|84.00|Upper limb amputation, not otherwise specified
C0186399|ICD9CM|AB|84.00|Upper limb amputat NOS
C0186418|ICD9CM|PT|80.71|Synovectomy, shoulder
C0186418|ICD9CM|AB|80.71|Shoulder synovectomy
C0186423|ICD9CM|PT|80.31|Biopsy of joint structure, shoulder
C0186423|ICD9CM|AB|80.31|Shoulder joint biopsy
C0186428|ICD9CM|PT|84.08|Disarticulation of shoulder
C0186428|ICD9CM|AB|84.08|Shoulder disarticulation
C0186482|ICD9CM|AB|77.22|Humerus wedge osteotomy
C0186482|ICD9CM|PT|77.22|Wedge osteotomy, humerus
C0186483|ICD9CM|AB|77.42|Humerus biopsy
C0186483|ICD9CM|PT|77.42|Biopsy of bone, humerus
C0186485|ICD9CM|PT|77.62|Local excision of lesion or tissue of bone, humerus
C0186485|ICD9CM|AB|77.62|Loc exc bone les humerus
C0186487|ICD9CM|AB|77.92|Total ostectomy-humerus
C0186487|ICD9CM|PT|77.92|Total ostectomy, humerus
C0186488|ICD9CM|PT|77.72|Excision of bone for graft, humerus
C0186488|ICD9CM|AB|77.72|Excise humerus for graft
C0186489|ICD9CM|PT|79.61|Debridement of open fracture site, humerus
C0186489|ICD9CM|AB|79.61|Debrid open fx-humerus
C0186493|ICD9CM|PT|80.32|Biopsy of joint structure, elbow
C0186493|ICD9CM|AB|80.32|Elbow joint biopsy
C0186495|ICD9CM|PT|80.72|Synovectomy, elbow
C0186495|ICD9CM|AB|80.72|Elbow synovectomy
C0186526|ICD9CM|PT|77.23|Wedge osteotomy, radius and ulna
C0186526|ICD9CM|AB|77.23|Radius/ulna wedg osteoto
C0186538|ICD9CM|PT|77.73|Excision of bone for graft, radius and ulna
C0186538|ICD9CM|AB|77.73|Excis radius/ulna-graft
C0186539|ICD9CM|PT|84.05|Amputation through forearm
C0186539|ICD9CM|AB|84.05|Amputation thru forearm
C0186547|ICD9CM|AB|77.43|Radius & ulna biopsy
C0186547|ICD9CM|PT|77.43|Biopsy of bone, radius and ulna
C0186550|ICD9CM|PT|77.63|Local excision of lesion or tissue of bone, radius and ulna
C0186550|ICD9CM|AB|77.63|Loc exc les radius/ulna
C0186554|ICD9CM|PT|77.93|Total ostectomy, radius and ulna
C0186554|ICD9CM|AB|77.93|Tot ostect-radius/ulna
C0186555|ICD9CM|PT|79.62|Debridement of open fracture site, radius and ulna
C0186555|ICD9CM|AB|79.62|Debrid opn fx-radius/uln
C0186562|ICD9CM|PT|84.44|Implantation of prosthetic device of arm
C0186562|ICD9CM|AB|84.44|Implant arm prosthesis
C0186573|ICD9CM|PT|78.92|Insertion of bone growth stimulator, humerus
C0186573|ICD9CM|AB|78.92|Insert bone stim-humerus
C0186581|ICD9CM|PT|78.93|Insertion of bone growth stimulator, radius and ulna
C0186581|ICD9CM|AB|78.93|Inser bone stim-rad/ulna
C0186599|ICD9CM|PT|80.22|Arthroscopy, elbow
C0186599|ICD9CM|AB|80.22|Elbow arthroscopy
C0186643|ICD9CM|PT|79.81|Open reduction of dislocation of shoulder
C0186643|ICD9CM|AB|79.81|Opn reduc disloc-shouldr
C0186650|ICD9CM|AB|81.23|Arthrodesis of shoulder
C0186650|ICD9CM|PT|81.23|Arthrodesis of shoulder
C0186658|ICD9CM|PT|81.81|Partial shoulder replacement
C0186658|ICD9CM|AB|81.81|Partial shoulder replace
C0186659|ICD9CM|PT|81.82|Repair of recurrent dislocation of shoulder
C0186659|ICD9CM|AB|81.82|Rep recur shlder disloc
C0186666|ICD9CM|AB|83.63|Rotator cuff repair
C0186666|ICD9CM|PT|83.63|Rotator cuff repair
C0186771|ICD9CM|PT|78.52|Internal fixation of bone without fracture reduction, humerus
C0186771|ICD9CM|AB|78.52|Int fixation-humerus
C0186772|ICD9CM|PT|79.21|Open reduction of fracture without internal fixation, humerus
C0186772|ICD9CM|AB|79.21|Open reduc-humerus fx
C0186773|ICD9CM|PT|79.31|Open reduction of fracture with internal fixation, humerus
C0186773|ICD9CM|AB|79.31|Open red-int fix humerus
C0186774|ICD9CM|PT|79.51|Open reduction of separated epiphysis, humerus
C0186774|ICD9CM|AB|79.51|Opn red-sep epiphy-humer
C0186781|ICD9CM|AB|81.84|Total elbow replacement
C0186781|ICD9CM|PT|81.84|Total elbow replacement
C0186790|ICD9CM|AB|81.24|Arthrodesis of elbow
C0186790|ICD9CM|PT|81.24|Arthrodesis of elbow
C0186793|ICD9CM|PT|79.82|Open reduction of dislocation of elbow
C0186793|ICD9CM|AB|79.82|Open reduc-elbow disloc
C0186901|ICD9CM|PT|78.53|Internal fixation of bone without fracture reduction, radius and ulna
C0186901|ICD9CM|AB|78.53|Int fixation-radius/ulna
C0186907|ICD9CM|PT|79.52|Open reduction of separated epiphysis, radius and ulna
C0186907|ICD9CM|AB|79.52|Op red-radius/uln epiphy
C0186937|ICD9CM|PT|78.72|Osteoclasis, humerus
C0186937|ICD9CM|AB|78.72|Osteoclasis-humerus
C0186958|ICD9CM|AB|78.03|Bone graft-radius/ulna
C0186958|ICD9CM|PT|78.03|Bone graft, radius and ulna
C0186961|ICD9CM|PT|78.02|Bone graft, humerus
C0186961|ICD9CM|AB|78.02|Bone graft to humerus
C0186986|ICD9CM|PT|79.71|Closed reduction of dislocation of shoulder
C0186986|ICD9CM|AB|79.71|Cl reduc disloc-shoulder
C0187018|ICD9CM|PT|79.11|Closed reduction of fracture with internal fixation, humerus
C0187018|ICD9CM|AB|79.11|Clos red-int fix humerus
C0187019|ICD9CM|PT|79.41|Closed reduction of separated epiphysis, humerus
C0187019|ICD9CM|AB|79.41|Close red-humerus epiphy
C0187023|ICD9CM|PT|79.72|Closed reduction of dislocation of elbow
C0187023|ICD9CM|AB|79.72|Cl reduc disloc-elbow
C0187048|ICD9CM|PT|79.12|Closed reduction of fracture with internal fixation, radius and ulna
C0187048|ICD9CM|AB|79.12|Cl red-int fix rad/ulna
C0187051|ICD9CM|PT|79.42|Closed reduction of separated epiphysis, radius and ulna
C0187051|ICD9CM|AB|79.42|Cls red-radius/ul epiphy
C0187065|ICD9CM|PT|78.84|Diagnostic procedures on bone, not elsewhere classified, carpals and metacarpals
C0187065|ICD9CM|AB|78.84|Oth dx proc-metacar/car
C0187066|ICD9CM|PT|79.93|Unspecified operation on bone injury, carpals and metacarpals
C0187066|ICD9CM|AB|79.93|Metacarp/carp inj op NOS
C0187069|ICD9CM|HT|82|Operations on muscle, tendon, and fascia of hand
C0187075|ICD9CM|PT|79.94|Unspecified operation on bone injury, phalanges of hand
C0187075|ICD9CM|AB|79.94|Finger injury op NOS
C0187106|ICD9CM|PT|82.01|Exploration of tendon sheath of hand
C0187106|ICD9CM|AB|82.01|Explor tend sheath-hand
C0187116|ICD9CM|AB|82.03|Bursotomy of hand
C0187116|ICD9CM|PT|82.03|Bursotomy of hand
C0187120|ICD9CM|AB|82.02|Myotomy of hand
C0187120|ICD9CM|PT|82.02|Myotomy of hand
C0187137|ICD9CM|AB|82.11|Tenotomy of hand
C0187137|ICD9CM|PT|82.11|Tenotomy of hand
C0187138|ICD9CM|AB|82.12|Fasciotomy of hand
C0187138|ICD9CM|PT|82.12|Fasciotomy of hand
C0187144|ICD9CM|PT|82.92|Aspiration of bursa of hand
C0187144|ICD9CM|AB|82.92|Aspiration bursa of hand
C0187194|ICD9CM|PT|80.33|Biopsy of joint structure, wrist
C0187194|ICD9CM|AB|80.33|Wrist joint biopsy
C0187195|ICD9CM|PT|80.73|Synovectomy, wrist
C0187195|ICD9CM|AB|80.73|Wrist synovectomy
C0187205|ICD9CM|PT|77.24|Wedge osteotomy, carpals and metacarpals
C0187205|ICD9CM|AB|77.24|Metacar/car wedg osteoto
C0187209|ICD9CM|PT|77.94|Total ostectomy, carpals and metacarpals
C0187209|ICD9CM|AB|77.94|Tot ostect-metacarp/carp
C0187210|ICD9CM|PT|77.74|Excision of bone for graft, carpals and metacarpals
C0187210|ICD9CM|AB|77.74|Excis metacar/car-graft
C0187239|ICD9CM|PT|80.34|Biopsy of joint structure, hand and finger
C0187239|ICD9CM|AB|80.34|Hand/finger joint biopsy
C0187253|ICD9CM|PT|82.21|Excision of lesion of tendon sheath of hand
C0187253|ICD9CM|AB|82.21|Exc les tend sheath hand
C0187257|ICD9CM|PT|82.22|Excision of lesion of muscle of hand
C0187257|ICD9CM|AB|82.22|Excision hand muscle les
C0187267|ICD9CM|PT|82.32|Excision of tendon of hand for graft
C0187267|ICD9CM|AB|82.32|Excis hand tend for grft
C0187269|ICD9CM|AB|82.31|Bursectomy of hand
C0187269|ICD9CM|PT|82.31|Bursectomy of hand
C0187278|ICD9CM|AB|84.03|Amputation through hand
C0187278|ICD9CM|PT|84.03|Amputation through hand
C0187280|ICD9CM|PT|98.26|Removal of foreign body from hand without incision
C0187280|ICD9CM|AB|98.26|Removal FB from hand
C0187303|ICD9CM|PT|79.64|Debridement of open fracture site, phalanges of hand
C0187303|ICD9CM|AB|79.64|Debrid opn fx-finger
C0187320|ICD9CM|PT|78.94|Insertion of bone growth stimulator, carpals and metacarpals
C0187320|ICD9CM|AB|78.94|Inser bone stim-meta/car
C0187330|ICD9CM|PT|82.94|Injection of therapeutic substance into bursa of hand
C0187330|ICD9CM|AB|82.94|Inject bursa of hand
C0187332|ICD9CM|PT|82.95|Injection of therapeutic substance into tendon of hand
C0187332|ICD9CM|AB|82.95|Inject tendon of hand
C0187394|ICD9CM|AB|81.26|Metacarpocarpal fusion
C0187394|ICD9CM|PT|81.26|Metacarpocarpal fusion
C0187401|ICD9CM|PT|79.83|Open reduction of dislocation of wrist
C0187401|ICD9CM|AB|79.83|Open reduc-wrist disloc
C0187402|ICD9CM|AB|81.25|Carporadial fusion
C0187402|ICD9CM|PT|81.25|Carporadial fusion
C0187442|ICD9CM|PT|78.54|Internal fixation of bone without fracture reduction, carpals and metacarpals
C0187442|ICD9CM|AB|78.54|Int fixation-metacar/car
C0187443|ICD9CM|PT|79.33|Open reduction of fracture with internal fixation, carpals and metacarpals
C0187443|ICD9CM|AB|79.33|Op red-int fix metac/car
C0187489|ICD9CM|PT|82.71|Tendon pulley reconstruction of hand
C0187489|ICD9CM|AB|82.71|Hand tend pulley reconst
C0187495|ICD9CM|AB|82.82|Repair of cleft hand
C0187495|ICD9CM|PT|82.82|Repair of cleft hand
C0187501|ICD9CM|PT|79.34|Open reduction of fracture with internal fixation, phalanges of hand
C0187501|ICD9CM|AB|79.34|Open red-int fix finger
C0187504|ICD9CM|PT|82.53|Reattachment of tendon of hand
C0187504|ICD9CM|AB|82.53|Hand tendon reattachment
C0187505|ICD9CM|PT|82.54|Reattachment of muscle of hand
C0187505|ICD9CM|AB|82.54|Hand muscle reattachment
C0187606|ICD9CM|PT|81.27|Metacarpophalangeal fusion
C0187606|ICD9CM|AB|81.27|Metacarpophalangeal fus
C0187622|ICD9CM|PT|81.71|Arthroplasty of metacarpophalangeal and interphalangeal joint with implant
C0187622|ICD9CM|AB|81.71|Arthroplas metacarp wit
C0187630|ICD9CM|AB|82.84|Repair of mallet finger
C0187630|ICD9CM|PT|82.84|Repair of mallet finger
C0187638|ICD9CM|PT|82.41|Suture of tendon sheath of hand
C0187638|ICD9CM|AB|82.41|Suture tendn sheath hand
C0187643|ICD9CM|PT|82.42|Delayed suture of flexor tendon of hand
C0187643|ICD9CM|AB|82.42|Delay sut flex tend hand
C0187661|ICD9CM|PT|82.91|Lysis of adhesions of hand
C0187661|ICD9CM|AB|82.91|Lysis of hand adhesions
C0187693|ICD9CM|PT|82.51|Advancement of tendon of hand
C0187693|ICD9CM|AB|82.51|Hand tendon advancement
C0187695|ICD9CM|PT|82.52|Recession of tendon of hand
C0187695|ICD9CM|AB|82.52|Hand tendon recession
C0187715|ICD9CM|PT|82.81|Transfer of finger, except thumb
C0187715|ICD9CM|AB|82.81|Transfer of finger
C0187718|ICD9CM|PT|79.73|Closed reduction of dislocation of wrist
C0187718|ICD9CM|AB|79.73|Cl reduc disloc-wrist
C0187732|ICD9CM|PT|79.13|Closed reduction of fracture with internal fixation, carpals and metacarpals
C0187732|ICD9CM|AB|79.13|Cl red-int fix metac/car
C0187747|ICD9CM|PT|79.14|Closed reduction of fracture with internal fixation, phalanges of hand
C0187747|ICD9CM|AB|79.14|Close red-int fix finger
C0187767|ICD9CM|PT|78.85|Diagnostic procedures on bone, not elsewhere classified, femur
C0187767|ICD9CM|AB|78.85|Oth dx proced-femur
C0187768|ICD9CM|PT|79.95|Unspecified operation on bone injury, femur
C0187768|ICD9CM|AB|79.95|Femur injury op NOS
C0187770|ICD9CM|PT|78.86|Diagnostic procedures on bone, not elsewhere classified, patella
C0187770|ICD9CM|AB|78.86|Oth dx proced-patella
C0187772|ICD9CM|PT|78.87|Diagnostic procedures on bone, not elsewhere classified, tibia and fibula
C0187772|ICD9CM|AB|78.87|Oth dx proc-tibia/fibula
C0187775|ICD9CM|PT|79.96|Unspecified operation on bone injury, tibia and fibula
C0187775|ICD9CM|AB|79.96|Tibia/fibula inj op NOS
C0187841|ICD9CM|PT|98.29|Removal of foreign body without incision from lower limb, except foot
C0187841|ICD9CM|AB|98.29|Removal FB from leg
C0187857|ICD9CM|PT|77.65|Local excision of lesion or tissue of bone, femur
C0187857|ICD9CM|AB|77.65|Loc exc bone les femur
C0187858|ICD9CM|PT|77.75|Excision of bone for graft, femur
C0187858|ICD9CM|AB|77.75|Excise femur for graft
C0187861|ICD9CM|PT|77.95|Total ostectomy, femur
C0187861|ICD9CM|AB|77.95|Tot ostectomy-femur
C0187862|ICD9CM|PT|79.65|Debridement of open fracture site, femur
C0187862|ICD9CM|AB|79.65|Debrid opn fx-femur
C0187863|ICD9CM|PT|77.05|Sequestrectomy, femur
C0187863|ICD9CM|AB|77.05|Femoral sequestrectomy
C0187890|ICD9CM|PT|77.26|Wedge osteotomy, patella
C0187890|ICD9CM|AB|77.26|Patellar wedge osteotomy
C0187891|ICD9CM|PT|77.06|Sequestrectomy, patella
C0187891|ICD9CM|AB|77.06|Patellar sequestrectomy
C0187893|ICD9CM|PT|77.66|Local excision of lesion or tissue of bone, patella
C0187893|ICD9CM|AB|77.66|Loc exc bone les patella
C0187897|ICD9CM|PT|79.86|Open reduction of dislocation of knee
C0187897|ICD9CM|AB|79.86|Open reduc-knee dislocat
C0187898|ICD9CM|PT|77.96|Total ostectomy, patella
C0187898|ICD9CM|AB|77.96|Total patellectomy
C0187900|ICD9CM|PT|80.36|Biopsy of joint structure, knee
C0187900|ICD9CM|AB|80.36|Knee joint biopsy
C0187901|ICD9CM|PT|80.6|Excision of semilunar cartilage of knee
C0187901|ICD9CM|AB|80.6|Excis knee semilun cartl
C0187903|ICD9CM|PT|80.76|Synovectomy, knee
C0187903|ICD9CM|AB|80.76|Knee synovectomy
C0187906|ICD9CM|AB|84.16|Disarticulation of knee
C0187906|ICD9CM|PT|84.16|Disarticulation of knee
C0187922|ICD9CM|PT|77.77|Excision of bone for graft, tibia and fibula
C0187922|ICD9CM|AB|77.77|Excise tib/fib for graft
C0187927|ICD9CM|PT|77.07|Sequestrectomy, tibia and fibula
C0187927|ICD9CM|AB|77.07|Tibia/fibula sequestrec
C0187936|ICD9CM|PT|77.67|Local excision of lesion or tissue of bone, tibia and fibula
C0187936|ICD9CM|AB|77.67|Loc exc les tibia/fibula
C0187938|ICD9CM|PT|77.97|Total ostectomy, tibia and fibula
C0187938|ICD9CM|AB|77.97|Tot ostect-tibia/fibula
C0187941|ICD9CM|PT|79.66|Debridement of open fracture site, tibia and fibula
C0187941|ICD9CM|AB|79.66|Debrid opn fx-tibia/fib
C0187948|ICD9CM|PT|84.48|Implantation of prosthetic device of leg
C0187948|ICD9CM|AB|84.48|Implant leg prosthesis
C0187953|ICD9CM|PT|78.95|Insertion of bone growth stimulator, femur
C0187953|ICD9CM|AB|78.95|Insert bone stim-femur
C0187958|ICD9CM|PT|78.96|Insertion of bone growth stimulator, patella
C0187958|ICD9CM|AB|78.96|Insert bone stim-patella
C0187965|ICD9CM|PT|78.97|Insertion of bone growth stimulator, tibia and fibula
C0187965|ICD9CM|AB|78.97|Inser bone stim-tib/fib
C0188093|ICD9CM|AB|78.55|Internal fixation-femur
C0188093|ICD9CM|PT|78.55|Internal fixation of bone without fracture reduction, femur
C0188094|ICD9CM|PT|79.55|Open reduction of separated epiphysis, femur
C0188094|ICD9CM|AB|79.55|Opn red-sep epiphy-femur
C0188107|ICD9CM|AB|83.86|Quadricepsplasty
C0188107|ICD9CM|PT|83.86|Quadricepsplasty
C0188109|ICD9CM|PT|79.35|Open reduction of fracture with internal fixation, femur
C0188109|ICD9CM|AB|79.35|Open reduc-int fix femur
C0188172|ICD9CM|AB|81.22|Arthrodesis of knee
C0188172|ICD9CM|PT|81.22|Arthrodesis of knee
C0188173|ICD9CM|PT|78.56|Internal fixation of bone without fracture reduction, patella
C0188173|ICD9CM|AB|78.56|Internal fix-patella
C0188174|ICD9CM|PT|77.76|Excision of bone for graft, patella
C0188174|ICD9CM|AB|77.76|Excise patella for graft
C0188181|ICD9CM|PT|81.42|Five-in-one repair of knee
C0188181|ICD9CM|AB|81.42|Five-in-one knee repair
C0188182|ICD9CM|AB|81.43|Triad knee repair
C0188182|ICD9CM|PT|81.43|Triad knee repair
C0188210|ICD9CM|PT|79.36|Open reduction of fracture with internal fixation, tibia and fibula
C0188210|ICD9CM|AB|79.36|Op red-int fix tib/fibul
C0188260|ICD9CM|PT|78.57|Internal fixation of bone without fracture reduction, tibia and fibula
C0188260|ICD9CM|AB|78.57|Int fixation-tibia/fibul
C0188273|ICD9CM|PT|79.56|Open reduction of separated epiphysis, tibia and fibula
C0188273|ICD9CM|AB|79.56|Op red-tibia/fib epiphys
C0188292|ICD9CM|PT|78.75|Osteoclasis, femur
C0188292|ICD9CM|AB|78.75|Osteoclasis-femur
C0188293|ICD9CM|PT|78.76|Osteoclasis, patella
C0188293|ICD9CM|AB|78.76|Osteoclasis-patella
C0188299|ICD9CM|AB|78.77|Osteoclasis-tibia/fibula
C0188299|ICD9CM|PT|78.77|Osteoclasis, tibia and fibula
C0188310|ICD9CM|PT|78.05|Bone graft, femur
C0188310|ICD9CM|AB|78.05|Bone graft to femur
C0188313|ICD9CM|AB|78.06|Bone graft to patella
C0188313|ICD9CM|PT|78.06|Bone graft, patella
C0188334|ICD9CM|PT|84.45|Fitting of prosthesis above knee
C0188334|ICD9CM|AB|84.45|Fit above knee prosthes
C0188354|ICD9CM|PT|79.45|Closed reduction of separated epiphysis, femur
C0188354|ICD9CM|AB|79.45|Close reduc-femur epiphy
C0188373|ICD9CM|PT|84.46|Fitting of prosthesis below knee
C0188373|ICD9CM|AB|84.46|Fit below knee prosthes
C0188377|ICD9CM|PT|79.15|Closed reduction of fracture with internal fixation, femur
C0188377|ICD9CM|AB|79.15|Closed red-int fix femur
C0188382|ICD9CM|PT|79.76|Closed reduction of dislocation of knee
C0188382|ICD9CM|AB|79.76|Cl reduc disloc-knee
C0188402|ICD9CM|PT|79.16|Closed reduction of fracture with internal fixation, tibia and fibula
C0188402|ICD9CM|AB|79.16|Cl red-int fix tib/fibu
C0188407|ICD9CM|PT|79.46|Closed reduction of separated epiphysis, tibia and fibula
C0188407|ICD9CM|AB|79.46|Cls red-tibia/fib epiphy
C0188414|ICD9CM|PT|78.88|Diagnostic procedures on bone, not elsewhere classified, tarsals and metatarsals
C0188414|ICD9CM|AB|78.88|Oth dx proc-metatar/tar
C0188415|ICD9CM|PT|79.97|Unspecified operation on bone injury, tarsals and metatarsals
C0188415|ICD9CM|AB|79.97|Metatars/tars inj op NOS
C0188417|ICD9CM|PT|79.98|Unspecified operation on bone injury, phalanges of foot
C0188417|ICD9CM|AB|79.98|Toe injury operation NOS
C0188472|ICD9CM|AB|83.11|Achillotenotomy
C0188472|ICD9CM|PT|83.11|Achillotenotomy
C0188494|ICD9CM|AB|84.13|Disarticulation of ankle
C0188494|ICD9CM|PT|84.13|Disarticulation of ankle
C0188496|ICD9CM|PT|80.37|Biopsy of joint structure, ankle
C0188496|ICD9CM|AB|80.37|Ankle joint biopsy
C0188497|ICD9CM|PT|80.77|Synovectomy, ankle
C0188497|ICD9CM|AB|80.77|Ankle synovectomy
C0188570|ICD9CM|PT|79.67|Debridement of open fracture site, tarsals and metatarsals
C0188570|ICD9CM|AB|79.67|Debrid opn fx-metat/tar
C0188571|ICD9CM|PT|79.68|Debridement of open fracture site, phalanges of foot
C0188571|ICD9CM|AB|79.68|Debrid opn fx-toe
C0188579|ICD9CM|AB|77.48|Metatarsal/tarsal biopsy
C0188579|ICD9CM|PT|77.48|Biopsy of bone, tarsals and metatarsals
C0188582|ICD9CM|PT|77.78|Excision of bone for graft, tarsals and metatarsals
C0188582|ICD9CM|AB|77.78|Excis metatar/tar-graft
C0188585|ICD9CM|PT|77.51|Bunionectomy with soft tissue correction and osteotomy of the first metatarsal
C0188585|ICD9CM|AB|77.51|Bunionect/sft/osteotomy
C0188591|ICD9CM|PT|80.38|Biopsy of joint structure, foot and toe
C0188591|ICD9CM|AB|80.38|Foot & toe joint biopsy
C0188596|ICD9CM|PT|77.98|Total ostectomy, tarsals and metatarsals
C0188596|ICD9CM|AB|77.98|Tot ostect-metatars/tars
C0188601|ICD9CM|PT|77.28|Wedge osteotomy, tarsals and metatarsals
C0188601|ICD9CM|AB|77.28|Metatar/tar wedg osteot
C0188602|ICD9CM|PT|84.11|Amputation of toe
C0188602|ICD9CM|AB|84.11|Toe amputation
C0188617|ICD9CM|PT|78.98|Insertion of bone growth stimulator, tarsals and metatarsals
C0188617|ICD9CM|AB|78.98|Inser bone stim-meta/tar
C0188624|ICD9CM|PT|80.27|Arthroscopy, ankle
C0188624|ICD9CM|AB|80.27|Ankle arthroscopy
C0188661|ICD9CM|AB|81.11|Ankle fusion
C0188661|ICD9CM|PT|81.11|Ankle fusion
C0188664|ICD9CM|AB|81.56|Total ankle replacement
C0188664|ICD9CM|PT|81.56|Total ankle replacement
C0188665|ICD9CM|PT|79.87|Open reduction of dislocation of ankle
C0188665|ICD9CM|AB|79.87|Open reduc-ankle disloc
C0188673|ICD9CM|AB|81.13|Subtalar fusion
C0188673|ICD9CM|PT|81.13|Subtalar fusion
C0188725|ICD9CM|AB|77.56|Repair of hammer toe
C0188725|ICD9CM|PT|77.56|Repair of hammer toe
C0188740|ICD9CM|PT|77.52|Bunionectomy with soft tissue correction and arthrodesis
C0188740|ICD9CM|AB|77.52|Bunionect/sft/arthrodes
C0188743|ICD9CM|PT|77.53|Other bunionectomy with soft tissue correction
C0188743|ICD9CM|AB|77.53|Oth bunionect w sft corr
C0188822|ICD9CM|AB|81.15|Tarsometatarsal fusion
C0188822|ICD9CM|PT|81.15|Tarsometatarsal fusion
C0188827|ICD9CM|AB|81.14|Midtarsal fusion
C0188827|ICD9CM|PT|81.14|Midtarsal fusion
C0188832|ICD9CM|PT|81.16|Metatarsophalangeal fusion
C0188832|ICD9CM|AB|81.16|Metatarsophalangeal fus
C0188844|ICD9CM|PT|78.58|Internal fixation of bone without fracture reduction, tarsals and metatarsals
C0188844|ICD9CM|AB|78.58|Int fixation-metatar/tar
C0188847|ICD9CM|PT|79.37|Open reduction of fracture with internal fixation, tarsals and metatarsals
C0188847|ICD9CM|AB|79.37|Op red-int fix metat/tar
C0188849|ICD9CM|PT|79.38|Open reduction of fracture with internal fixation, phalanges of foot
C0188849|ICD9CM|AB|79.38|Open reduct-int fix toe
C0188850|ICD9CM|PT|79.88|Open reduction of dislocation of foot and toe
C0188850|ICD9CM|AB|79.88|Opn reduc disloc-ft/toe
C0188866|ICD9CM|PT|81.57|Replacement of joint of foot and toe
C0188866|ICD9CM|AB|81.57|Repl joint of foot, toe
C0188918|ICD9CM|PT|79.77|Closed reduction of dislocation of ankle
C0188918|ICD9CM|AB|79.77|Cl reduc disloc-ankle
C0188954|ICD9CM|PT|79.17|Closed reduction of fracture with internal fixation, tarsals and metatarsals
C0188954|ICD9CM|AB|79.17|Cl red-int fix metat/tar
C0188955|ICD9CM|PT|79.18|Closed reduction of fracture with internal fixation, phalanges of foot
C0188955|ICD9CM|AB|79.18|Close red-int fix toe fx
C0188958|ICD9CM|PT|79.78|Closed reduction of dislocation of foot and toe
C0188958|ICD9CM|AB|79.78|Cl reduc disloc-foot/toe
C0188970|ICD9CM|HT|21|Operations on nose
C0188972|ICD9CM|HT|21.0|Control of epistaxis
C0188972|ICD9CM|AB|21.00|Control of epistaxis NOS
C0188972|ICD9CM|PT|21.00|Control of epistaxis, not otherwise specified
C0188974|ICD9CM|AB|21.1|Incision of nose
C0188974|ICD9CM|PT|21.1|Incision of nose
C0188990|ICD9CM|PT|98.12|Removal of intraluminal foreign body from nose without incision
C0188990|ICD9CM|AB|98.12|Remov intralum nose FB
C0188993|ICD9CM|PT|21.5|Submucous resection of nasal septum
C0188993|ICD9CM|AB|21.5|Submuc nasal sept resect
C0189015|ICD9CM|PT|21.02|Control of epistaxis by posterior (and anterior) packing
C0189015|ICD9CM|AB|21.02|Post nasal pac for epist
C0189016|ICD9CM|PT|97.21|Replacement of nasal packing
C0189016|ICD9CM|AB|97.21|Replace nasal packing
C0189024|ICD9CM|AB|21.21|Rhinoscopy
C0189024|ICD9CM|PT|21.21|Rhinoscopy
C0189030|ICD9CM|PT|21.81|Suture of laceration of nose
C0189030|ICD9CM|AB|21.81|Nasal laceration suture
C0189037|ICD9CM|PT|21.72|Open reduction of nasal fracture
C0189037|ICD9CM|AB|21.72|Open reduction nasal fx
C0189040|ICD9CM|PT|21.04|Control of epistaxis by ligation of ethmoidal arteries
C0189040|ICD9CM|AB|21.04|Ethmoid art ligat-epist
C0189041|ICD9CM|PT|21.05|Control of epistaxis by (transantral) ligation of the maxillary artery
C0189041|ICD9CM|AB|21.05|Max art lig for epistax
C0189042|ICD9CM|AB|21.86|Limited rhinoplasty
C0189042|ICD9CM|PT|21.86|Limited rhinoplasty
C0189047|ICD9CM|PT|21.83|Total nasal reconstruction
C0189047|ICD9CM|AB|21.83|Tot nasal reconstruction
C0189051|ICD9CM|AB|21.84|Revision rhinoplasty
C0189051|ICD9CM|PT|21.84|Revision rhinoplasty
C0189064|ICD9CM|PT|21.03|Control of epistaxis by cauterization (and packing)
C0189064|ICD9CM|AB|21.03|Cautery to stop epistax
C0189071|ICD9CM|PT|21.91|Lysis of adhesions of nose
C0189071|ICD9CM|AB|21.91|Lysis of nasal adhesions
C0189090|ICD9CM|PT|21.71|Closed reduction of nasal fracture
C0189090|ICD9CM|AB|21.71|Clos reduction nasal fx
C0189094|ICD9CM|PT|96.21|Dilation of frontonasal duct
C0189094|ICD9CM|AB|96.21|Dilat frontonasal duct
C0189111|ICD9CM|PT|22.31|Radical maxillary antrotomy
C0189111|ICD9CM|AB|22.31|Radical maxillary antrot
C0189113|ICD9CM|AB|22.41|Frontal sinusotomy
C0189113|ICD9CM|PT|22.41|Frontal sinusotomy
C0189123|ICD9CM|AB|22.51|Ethmoidotomy
C0189123|ICD9CM|PT|22.51|Ethmoidotomy
C0189124|ICD9CM|AB|22.52|Sphenoidotomy
C0189124|ICD9CM|PT|22.52|Sphenoidotomy
C0189137|ICD9CM|PT|22.61|Excision of lesion of maxillary sinus with Caldwell-Luc approach
C0189137|ICD9CM|AB|22.61|C-luc exc max sinus les
C0189146|ICD9CM|AB|22.42|Frontal sinusectomy
C0189146|ICD9CM|PT|22.42|Frontal sinusectomy
C0189149|ICD9CM|AB|22.63|Ethmoidectomy
C0189149|ICD9CM|PT|22.63|Ethmoidectomy
C0189156|ICD9CM|AB|22.64|Sphenoidectomy
C0189156|ICD9CM|PT|22.64|Sphenoidectomy
C0189160|ICD9CM|HT|22.0|Aspiration and lavage of nasal sinus
C0189160|ICD9CM|PT|22.00|Aspiration and lavage of nasal sinus, not otherwise specified
C0189160|ICD9CM|AB|22.00|Sinus aspirat/lavage NOS
C0189186|ICD9CM|HT|22.7|Repair of nasal sinus
C0189193|ICD9CM|PT|22.71|Closure of nasal sinus fistula
C0189193|ICD9CM|AB|22.71|Nasal sinus fistula clos
C0189222|ICD9CM|AB|30.22|Vocal cordectomy
C0189222|ICD9CM|PT|30.22|Vocal cordectomy
C0189224|ICD9CM|AB|30.21|Epiglottidectomy
C0189224|ICD9CM|PT|30.21|Epiglottidectomy
C0189231|ICD9CM|AB|30.3|Complete laryngectomy
C0189231|ICD9CM|PT|30.3|Complete laryngectomy
C0189233|ICD9CM|AB|30.1|Hemilaryngectomy
C0189233|ICD9CM|PT|30.1|Hemilaryngectomy
C0189253|ICD9CM|AB|31.0|Injection of larynx
C0189253|ICD9CM|PT|31.0|Injection of larynx
C0189261|ICD9CM|PT|96.02|Insertion of oropharyngeal airway
C0189261|ICD9CM|AB|96.02|Insert oropharyn airway
C0189299|ICD9CM|HT|31.6|Repair of larynx
C0189300|ICD9CM|AB|31.63|Laryngostomy revision
C0189300|ICD9CM|PT|31.63|Revision of laryngostomy
C0189305|ICD9CM|PT|30.01|Marsupialization of laryngeal cyst
C0189305|ICD9CM|AB|30.01|Larynx cyst marsupializ
C0189346|ICD9CM|AB|31.21|Mediastinal tracheostomy
C0189346|ICD9CM|PT|31.21|Mediastinal tracheostomy
C0189347|ICD9CM|AB|33.0|Incision of bronchus
C0189347|ICD9CM|PT|33.0|Incision of bronchus
C0189361|ICD9CM|PT|33.25|Open biopsy of bronchus
C0189361|ICD9CM|AB|33.25|Open bronchial biopsy
C0189388|ICD9CM|PT|31.44|Closed [endoscopic] biopsy of trachea
C0189388|ICD9CM|AB|31.44|Closed biopsy trachea
C0189391|ICD9CM|AB|33.22|Fiber-optic bronchoscopy
C0189391|ICD9CM|PT|33.22|Fiber-optic bronchoscopy
C0189426|ICD9CM|AB|31.72|Closure of tracheostomy
C0189426|ICD9CM|PT|31.72|Closure of external fistula of trachea
C0189427|ICD9CM|AB|31.74|Revision of tracheostomy
C0189427|ICD9CM|PT|31.74|Revision of tracheostomy
C0189456|ICD9CM|PT|33.92|Ligation of bronchus
C0189456|ICD9CM|AB|33.92|Bronchial ligation
C0189463|ICD9CM|AB|33.91|Bronchial dilation
C0189463|ICD9CM|PT|33.91|Bronchial dilation
C0189471|ICD9CM|AB|33.1|Incision of lung
C0189471|ICD9CM|PT|33.1|Incision of lung
C0189477|ICD9CM|AB|34.91|Thoracentesis
C0189477|ICD9CM|PT|34.91|Thoracentesis
C0189488|ICD9CM|HT|32.3|Segmental resection of lung
C0189497|ICD9CM|HT|32.4|Lobectomy of lung
C0189507|ICD9CM|PT|32.21|Plication of emphysematous bleb
C0189507|ICD9CM|AB|32.21|Emphysema bleb plication
C0189551|ICD9CM|HT|33.3|Surgical collapse of lung
C0189557|ICD9CM|AB|34.6|Scarification of pleura
C0189557|ICD9CM|PT|34.6|Scarification of pleura
C0189575|ICD9CM|HT|38.2|Diagnostic procedures on blood vessels
C0189577|ICD9CM|PT|39.41|Control of hemorrhage following vascular surgery
C0189577|ICD9CM|AB|39.41|Postop vasc op hem contr
C0189579|ICD9CM|HT|38.0|Incision of vessel
C0189579|ICD9CM|AB|38.00|Incision of vessel NOS
C0189579|ICD9CM|PT|38.00|Incision of vessel, unspecified site
C0189594|ICD9CM|PT|38.21|Biopsy of blood vessel
C0189594|ICD9CM|AB|38.21|Blood vessel biopsy
C0189606|ICD9CM|HT|38.3|Resection of vessel with anastomosis
C0189606|ICD9CM|PT|38.30|Resection of vessel with anastomosis, unspecified site
C0189606|ICD9CM|AB|38.30|Vessel resect/anast NOS
C0189617|ICD9CM|HT|38.4|Resection of vessel with replacement
C0189622|ICD9CM|PT|39.93|Insertion of vessel-to-vessel cannula
C0189622|ICD9CM|AB|39.93|Insert ves-to-ves cannul
C0189634|ICD9CM|PT|96.57|Irrigation of vascular catheter
C0189634|ICD9CM|AB|96.57|Vascular cath irrigation
C0189635|ICD9CM|AB|39.96|Total body perfusion
C0189635|ICD9CM|PT|39.96|Total body perfusion
C0189649|ICD9CM|PT|39.43|Removal of arteriovenous shunt for renal dialysis
C0189649|ICD9CM|AB|39.43|Remov ren dialysis shunt
C0189662|ICD9CM|PT|39.53|Repair of arteriovenous fistula
C0189662|ICD9CM|AB|39.53|Arterioven fistula rep
C0189693|ICD9CM|PT|39.27|Arteriovenostomy for renal dialysis
C0189693|ICD9CM|AB|39.27|Dialysis arteriovenostom
C0189700|ICD9CM|HT|39.4|Revision of vascular procedure
C0189711|ICD9CM|AB|39.51|Clipping of aneurysm
C0189711|ICD9CM|PT|39.51|Clipping of aneurysm
C0189746|ICD9CM|PT|39.62|Hypothermia (systemic) incidental to open heart surgery
C0189746|ICD9CM|AB|39.62|Hypothermia w open heart
C0189750|ICD9CM|PT|35.95|Revision of corrective procedure on heart
C0189750|ICD9CM|AB|35.95|Heart repair revision
C0189752|ICD9CM|PT|35.32|Operations on chordae tendineae
C0189752|ICD9CM|AB|35.32|Chordae tendineae ops
C0189753|ICD9CM|PT|35.35|Operations on trabeculae carneae cordis
C0189753|ICD9CM|AB|35.35|Trabecul carneae cord op
C0189758|ICD9CM|AB|37.10|Incision of heart NOS
C0189758|ICD9CM|AB|37.11|Cardiotomy
C0189758|ICD9CM|PT|37.11|Cardiotomy
C0189758|ICD9CM|PT|37.10|Incision of heart, not otherwise specified
C0189784|ICD9CM|PT|37.25|Biopsy of heart
C0189784|ICD9CM|AB|37.25|Cardiac biopsy
C0189786|ICD9CM|PT|37.32|Excision of aneurysm of heart
C0189786|ICD9CM|AB|37.32|Heart aneurysm excision
C0189815|ICD9CM|PT|37.92|Injection of therapeutic substance into heart
C0189815|ICD9CM|AB|37.92|Injection into heart
C0189824|ICD9CM|PT|37.72|Initial insertion of transvenous leads [electrodes] into atrium and ventricle
C0189824|ICD9CM|AB|37.72|Int inser lead atri-vent
C0189826|ICD9CM|PT|37.73|Initial insertion of transvenous lead [electrode] into atrium
C0189826|ICD9CM|AB|37.73|Int inser lead in atrium
C0189831|ICD9CM|PT|37.75|Revision of lead [electrode]
C0189831|ICD9CM|AB|37.75|Revision of lead
C0189846|ICD9CM|PT|37.81|Initial insertion of single-chamber device, not specified as rate responsive
C0189846|ICD9CM|AB|37.81|Int insert 1-cham, non
C0189847|ICD9CM|PT|37.82|Initial insertion of single-chamber device, rate responsive
C0189847|ICD9CM|AB|37.82|Int insert 1-cham, rate
C0189848|ICD9CM|PT|37.83|Initial insertion of dual-chamber device
C0189848|ICD9CM|AB|37.83|Int insert dual-cham dev
C0189856|ICD9CM|PT|37.86|Replacement of any type of pacemaker device with single-chamber device, rate responsive
C0189856|ICD9CM|AB|37.86|Repl pacem 1-cham, rate
C0189857|ICD9CM|PT|37.87|Replacement of any type pacemaker device with dual-chamber device
C0189857|ICD9CM|AB|37.87|Repl pacem w dual-cham
C0189868|ICD9CM|PT|37.96|Implantation of automatic cardioverter/defibrillator pulse generator only
C0189868|ICD9CM|AB|37.96|Implt cardiodefib genatr
C0189870|ICD9CM|PT|37.98|Replacement of automatic cardioverter/defibrillator pulse generator only
C0189870|ICD9CM|AB|37.98|Repl cardiodefib genratr
C0189883|ICD9CM|PT|37.63|Repair of heart assist system
C0189883|ICD9CM|AB|37.63|Repair heart assist sys
C0189887|ICD9CM|PT|37.77|Removal of lead(s) [electrode] without replacement
C0189887|ICD9CM|AB|37.77|Removal of lead w/o repl
C0189896|ICD9CM|PT|37.21|Right heart cardiac catheterization
C0189896|ICD9CM|AB|37.21|Rt heart cardiac cath
C0189897|ICD9CM|PT|37.22|Left heart cardiac catheterization
C0189897|ICD9CM|AB|37.22|Left heart cardiac cath
C0189898|ICD9CM|PT|37.23|Combined right and left heart cardiac catheterization
C0189898|ICD9CM|AB|37.23|Rt/left heart card cath
C0189920|ICD9CM|HT|37.4|Repair of heart and pericardium
C0189944|ICD9CM|PT|35.51|Repair of atrial septal defect with prosthesis, open technique
C0189944|ICD9CM|AB|35.51|Pros rep atrial def-opn
C0189954|ICD9CM|PT|35.60|Repair of unspecified septal defect of heart with tissue graft
C0189954|ICD9CM|AB|35.60|Grft repair hrt sept NOS
C0189959|ICD9CM|PT|35.62|Repair of ventricular septal defect with tissue graft
C0189959|ICD9CM|AB|35.62|Graft repair ventric def
C0189962|ICD9CM|PT|35.63|Repair of endocardial cushion defect with tissue graft
C0189962|ICD9CM|AB|35.63|Grft rep endocar cushion
C0189974|ICD9CM|PT|35.54|Repair of endocardial cushion defect with prosthesis
C0189974|ICD9CM|AB|35.54|Pros rep endocar cushion
C0189976|ICD9CM|PT|36.2|Heart revascularization by arterial implant
C0189976|ICD9CM|AB|36.2|Arterial implant revasc
C0189982|ICD9CM|PT|35.81|Total repair of tetralogy of fallot
C0189982|ICD9CM|AB|35.81|Tot repair tetral fallot
C0189998|ICD9CM|PT|35.83|Total repair of truncus arteriosus
C0189998|ICD9CM|AB|35.83|Tot rep truncus arterios
C0190009|ICD9CM|PT|35.93|Creation of conduit between left ventricle and aorta
C0190009|ICD9CM|AB|35.93|Conduit left ventr-aorta
C0190043|ICD9CM|PT|37.91|Open chest cardiac massage
C0190043|ICD9CM|AB|37.91|Opn chest cardiac massag
C0190066|ICD9CM|HT|35.3|Operations on structures adjacent to heart valves
C0190074|ICD9CM|PT|35.03|Closed heart valvotomy, pulmonary valve
C0190074|ICD9CM|AB|35.03|Closed pulmon valvotomy
C0190084|ICD9CM|PT|35.02|Closed heart valvotomy, mitral valve
C0190084|ICD9CM|AB|35.02|Closed mitral valvotomy
C0190086|ICD9CM|PT|35.01|Closed heart valvotomy, aortic valve
C0190086|ICD9CM|AB|35.01|Closed aortic valvotomy
C0190117|ICD9CM|PT|35.14|Open heart valvuloplasty of tricuspid valve without replacement
C0190117|ICD9CM|AB|35.14|Opn tricus valvuloplasty
C0190130|ICD9CM|PT|35.13|Open heart valvuloplasty of pulmonary valve without replacement
C0190130|ICD9CM|AB|35.13|Opn pulmon valvuloplasty
C0190150|ICD9CM|PT|35.12|Open heart valvuloplasty of mitral valve without replacement
C0190150|ICD9CM|AB|35.12|Opn mitral valvuloplasty
C0190155|ICD9CM|PT|35.11|Open heart valvuloplasty of aortic valve without replacement
C0190155|ICD9CM|AB|35.11|Opn aortic valvuloplasty
C0190165|ICD9CM|AB|35.33|Annuloplasty
C0190165|ICD9CM|PT|35.33|Annuloplasty
C0190175|ICD9CM|HT|35.1|Open heart valvuloplasty without replacement
C0190176|ICD9CM|PT|35.96|Percutaneous balloon valvuloplasty
C0190176|ICD9CM|AB|35.96|Perc balloon valvuplasty
C0190189|ICD9CM|HT|36|Operations on vessels of heart
C0190205|ICD9CM|PT|36.04|Intracoronary artery thrombolytic infusion
C0190205|ICD9CM|AB|36.04|Intrcoronry thromb infus
C0190214|ICD9CM|PT|36.91|Repair of aneurysm of coronary vessel
C0190214|ICD9CM|AB|36.91|Coron vess aneurysm rep
C0190224|ICD9CM|PT|36.11|(Aorto)coronary bypass of one coronary artery
C0190224|ICD9CM|AB|36.11|Aortocor bypas-1 cor art
C0190228|ICD9CM|PT|36.12|(Aorto)coronary bypass of two coronary arteries
C0190228|ICD9CM|AB|36.12|Aortocor bypas-2 cor art
C0190232|ICD9CM|PT|36.13|(Aorto)coronary bypass of three coronary arteries
C0190232|ICD9CM|AB|36.13|Aortocor bypas-3 cor art
C0190236|ICD9CM|PT|36.14|(Aorto)coronary bypass of four or more coronary arteries
C0190236|ICD9CM|AB|36.14|Aortcor bypas-4+ cor art
C0190242|ICD9CM|PT|36.16|Double internal mammary-coronary artery bypass
C0190242|ICD9CM|AB|36.16|2 int mam-cor art bypass
C0190267|ICD9CM|AB|38.04|Incision of aorta
C0190267|ICD9CM|PT|38.04|Incision of vessel, aorta
C0190280|ICD9CM|PT|38.34|Resection of vessel with anastomosis, aorta
C0190280|ICD9CM|AB|38.34|Aorta resection & anast
C0190305|ICD9CM|AB|38.14|Endarterectomy of aorta
C0190305|ICD9CM|PT|38.14|Endarterectomy, aorta
C0190338|ICD9CM|PT|38.44|Resection of vessel with replacement, aorta, abdominal
C0190338|ICD9CM|AB|38.44|Resect abdm aorta w repl
C0190368|ICD9CM|PT|39.54|Re-entry operation (aorta)
C0190368|ICD9CM|AB|39.54|Re-entry operation
C0190388|ICD9CM|PT|39.0|Systemic to pulmonary artery shunt
C0190388|ICD9CM|AB|39.0|Systemic-pulm art shunt
C0190431|ICD9CM|PT|39.25|Aorta-iliac-femoral bypass
C0190431|ICD9CM|AB|39.25|Aorta-iliac-femor bypass
C0190485|ICD9CM|PT|38.11|Endarterectomy, intracranial vessels
C0190485|ICD9CM|AB|38.11|Intracran endarterectomy
C0190568|ICD9CM|PT|99.64|Carotid sinus stimulation
C0190568|ICD9CM|AB|99.64|Carotid sinus stiumlat
C0190578|ICD9CM|PT|38.06|Incision of vessel, abdominal arteries
C0190578|ICD9CM|AB|38.06|Abdomen artery incision
C0190618|ICD9CM|PT|38.36|Resection of vessel with anastomosis, abdominal arteries
C0190618|ICD9CM|AB|38.36|Abd vessel resect/anast
C0190646|ICD9CM|PT|38.16|Endarterectomy, abdominal arteries
C0190646|ICD9CM|AB|38.16|Abdominal endarterectomy
C0190653|ICD9CM|PT|38.46|Resection of vessel with replacement, abdominal arteries
C0190653|ICD9CM|AB|38.46|Abd artery resec w repla
C0190763|ICD9CM|PT|39.21|Caval-pulmonary artery anastomosis
C0190763|ICD9CM|AB|39.21|Caval-pulmon art anastom
C0190809|ICD9CM|PT|38.08|Incision of vessel, lower limb arteries
C0190809|ICD9CM|AB|38.08|Lower limb artery incis
C0190822|ICD9CM|PT|38.13|Endarterectomy, upper limb vessels
C0190822|ICD9CM|AB|38.13|Upper limb endarterectom
C0190858|ICD9CM|PT|38.38|Resection of vessel with anastomosis, lower limb arteries
C0190858|ICD9CM|AB|38.38|Leg artery resect/anast
C0190863|ICD9CM|PT|38.18|Endarterectomy, lower limb arteries
C0190863|ICD9CM|AB|38.18|Lower limb endarterect
C0190998|ICD9CM|AB|38.07|Abdominal vein incision
C0190998|ICD9CM|PT|38.07|Incision of vessel, abdominal veins
C0191002|ICD9CM|AB|38.09|Lower limb vein incision
C0191002|ICD9CM|PT|38.09|Incision of vessel, lower limb veins
C0191018|ICD9CM|HT|38.5|Ligation and stripping of varicose veins
C0191072|ICD9CM|PT|38.37|Resection of vessel with anastomosis, abdominal veins
C0191072|ICD9CM|AB|38.37|Abd vein resect & anast
C0191095|ICD9CM|PT|38.39|Resection of vessel with anastomosis, lower limb veins
C0191095|ICD9CM|AB|38.39|Leg vein resect/anastom
C0191118|ICD9CM|PT|38.92|Umbilical vein catheterization
C0191118|ICD9CM|AB|38.92|Umbilical vein cath
C0191126|ICD9CM|PT|38.95|Venous catheterization for renal dialysis
C0191126|ICD9CM|AB|38.95|Ven cath renal dialysis
C0191172|ICD9CM|PT|38.7|Interruption of the vena cava
C0191172|ICD9CM|AB|38.7|Interruption vena cava
C0191234|ICD9CM|AB|37.0|Pericardiocentesis
C0191234|ICD9CM|PT|37.0|Pericardiocentesis
C0191244|ICD9CM|PT|37.24|Biopsy of pericardium
C0191244|ICD9CM|AB|37.24|Pericardial biopsy
C0191257|ICD9CM|PT|37.93|Injection of therapeutic substance into pericardium
C0191257|ICD9CM|AB|37.93|Injection into pericard
C0191274|ICD9CM|HT|85-86.99|OPERATIONS ON THE INTEGUMENTARY SYSTEM
C0191326|ICD9CM|PT|86.4|Radical excision of skin lesion
C0191326|ICD9CM|AB|86.4|Radical excis skin les
C0191402|ICD9CM|PT|98.18|Removal of intraluminal foreign body from artificial stoma without incision
C0191402|ICD9CM|AB|98.18|Remov intralum stoma FB
C0191427|ICD9CM|PT|86.85|Correction of syndactyly
C0191427|ICD9CM|AB|86.85|Syndactyly correction
C0191472|ICD9CM|PT|86.91|Excision of skin for graft
C0191472|ICD9CM|AB|86.91|Skin excision for graft
C0191483|ICD9CM|PT|86.72|Advancement of pedicle graft
C0191483|ICD9CM|AB|86.72|Pedicle graft advancemen
C0191498|ICD9CM|AB|86.66|Homograft to skin
C0191498|ICD9CM|PT|86.66|Homograft to skin
C0191625|ICD9CM|AB|86.51|Replantation of scalp
C0191625|ICD9CM|PT|86.51|Replantation of scalp
C0191626|ICD9CM|AB|86.64|Hair transplant
C0191626|ICD9CM|PT|86.64|Hair transplant
C0191654|ICD9CM|PT|86.21|Excision of pilonidal cyst or sinus
C0191654|ICD9CM|AB|86.21|Excision of pilonid cyst
C0191729|ICD9CM|PT|86.27|Debridement of nail, nail bed, or nail fold
C0191729|ICD9CM|AB|86.27|Debridement of nail
C0191796|ICD9CM|AB|86.86|Onychoplasty
C0191796|ICD9CM|PT|86.86|Onychoplasty
C0191835|ICD9CM|HT|85.1|Diagnostic procedures on breast
C0191840|ICD9CM|AB|85.0|Mastotomy
C0191840|ICD9CM|PT|85.0|Mastotomy
C0191846|ICD9CM|AB|85.91|Aspiration of breast
C0191846|ICD9CM|PT|85.91|Aspiration of breast
C0191864|ICD9CM|AB|85.25|Excision of nipple
C0191864|ICD9CM|PT|85.25|Excision of nipple
C0191879|ICD9CM|PT|85.42|Bilateral simple mastectomy
C0191879|ICD9CM|AB|85.42|Bilat simple mastectomy
C0191880|ICD9CM|PT|85.43|Unilateral extended simple mastectomy
C0191880|ICD9CM|AB|85.43|Unilat exten simp mastec
C0191881|ICD9CM|PT|85.44|Bilateral extended simple mastectomy
C0191881|ICD9CM|AB|85.44|Bilat extend simp mastec
C0191883|ICD9CM|PT|85.46|Bilateral radical mastectomy
C0191883|ICD9CM|AB|85.46|Bilat radical mastectomy
C0191895|ICD9CM|PT|85.33|Unilateral subcutaneous mammectomy with synchronous implant
C0191895|ICD9CM|AB|85.33|Unil subq mammect-implnt
C0191896|ICD9CM|PT|85.35|Bilateral subcutaneous mammectomy with synchronous implant
C0191896|ICD9CM|AB|85.35|Bil subq mammect-implant
C0191902|ICD9CM|PT|85.53|Unilateral breast implant
C0191902|ICD9CM|AB|85.53|Unilat breast implant
C0191909|ICD9CM|PT|85.94|Removal of implant of breast
C0191909|ICD9CM|AB|85.94|Breast implant removal
C0191912|ICD9CM|AB|85.92|Breast injection
C0191912|ICD9CM|PT|85.92|Injection of therapeutic agent into breast
C0191917|ICD9CM|PT|85.81|Suture of laceration of breast
C0191917|ICD9CM|AB|85.81|Suture breast laceration
C0191918|ICD9CM|AB|85.6|Mastopexy
C0191918|ICD9CM|PT|85.6|Mastopexy
C0191920|ICD9CM|PT|85.93|Revision of implant of breast
C0191920|ICD9CM|AB|85.93|Breast implant revision
C0191923|ICD9CM|PT|85.31|Unilateral reduction mammoplasty
C0191923|ICD9CM|AB|85.31|Unilat reduct mammoplast
C0191924|ICD9CM|PT|85.32|Bilateral reduction mammoplasty
C0191924|ICD9CM|AB|85.32|Bilat reduct mammoplasty
C0191925|ICD9CM|HT|85.5|Augmentation mammoplasty
C0191925|ICD9CM|PT|85.50|Augmentation mammoplasty, not otherwise specified
C0191925|ICD9CM|AB|85.50|Augment mammoplasty NOS
C0191937|ICD9CM|PT|85.84|Pedicle graft to breast
C0191937|ICD9CM|AB|85.84|Breast pedicle graft
C0191938|ICD9CM|PT|85.82|Split-thickness graft to breast
C0191938|ICD9CM|AB|85.82|Breast split-thick graft
C0191939|ICD9CM|PT|85.83|Full-thickness graft to breast
C0191939|ICD9CM|AB|85.83|Breast full-thick graft
C0191941|ICD9CM|PT|85.85|Muscle flap graft to breast
C0191941|ICD9CM|AB|85.85|Breast muscle flap graft
C0191943|ICD9CM|AB|85.86|Transposition of nipple
C0191943|ICD9CM|PT|85.86|Transposition of nipple
C0191960|ICD9CM|HT|27.7|Operations on uvula
C0191966|ICD9CM|AB|27.91|Labial frenotomy
C0191966|ICD9CM|PT|27.91|Labial frenotomy
C0191982|ICD9CM|AB|27.1|Incision of palate
C0191982|ICD9CM|PT|27.1|Incision of palate
C0191984|ICD9CM|AB|27.71|Incision of uvula
C0191984|ICD9CM|PT|27.71|Incision of uvula
C0191987|ICD9CM|PT|27.23|Biopsy of lip
C0191987|ICD9CM|AB|27.23|Lip biopsy
C0191994|ICD9CM|PT|27.41|Labial frenectomy
C0191994|ICD9CM|AB|27.41|Labial frenumectomy
C0192024|ICD9CM|AB|27.72|Excision of uvula
C0192024|ICD9CM|PT|27.72|Excision of uvula
C0192029|ICD9CM|PT|27.22|Biopsy of uvula and soft palate
C0192029|ICD9CM|AB|27.22|Uvula and soft palate bx
C0192061|ICD9CM|PT|27.53|Closure of fistula of mouth
C0192061|ICD9CM|AB|27.53|Closure of mouth fistula
C0192065|ICD9CM|PT|27.61|Suture of laceration of palate
C0192065|ICD9CM|AB|27.61|Suture of palate lacerat
C0192068|ICD9CM|AB|27.73|Repair of uvula
C0192068|ICD9CM|PT|27.73|Repair of uvula
C0192070|ICD9CM|AB|27.54|Repair of cleft lip
C0192070|ICD9CM|PT|27.54|Repair of cleft lip
C0192086|ICD9CM|PT|27.62|Correction of cleft palate
C0192086|ICD9CM|AB|27.62|Cleft palate correction
C0192100|ICD9CM|PT|27.63|Revision of cleft palate repair
C0192100|ICD9CM|AB|27.63|Revis cleft palat repair
C0192121|ICD9CM|PT|27.57|Attachment of pedicle or flap graft to lip and mouth
C0192121|ICD9CM|AB|27.57|Pedicle attach to mouth
C0192131|ICD9CM|PT|98.01|Removal of intraluminal foreign body from mouth without incision
C0192131|ICD9CM|AB|98.01|Remov intralum mouth FB
C0192135|ICD9CM|HT|25|Operations on tongue
C0192139|ICD9CM|AB|25.91|Lingual frenotomy
C0192139|ICD9CM|PT|25.91|Lingual frenotomy
C0192146|ICD9CM|AB|25.92|Lingual frenectomy
C0192146|ICD9CM|PT|25.92|Lingual frenectomy
C0192153|ICD9CM|AB|25.2|Partial glossectomy
C0192153|ICD9CM|PT|25.2|Partial glossectomy
C0192181|ICD9CM|PT|25.93|Lysis of adhesions of tongue
C0192181|ICD9CM|AB|25.93|Lysis of tongue adhesion
C0192189|ICD9CM|HT|29|Operations on pharynx
C0192198|ICD9CM|AB|29.0|Pharyngotomy
C0192198|ICD9CM|PT|29.0|Pharyngotomy
C0192207|ICD9CM|AB|29.31|Cricopharyngeal myotomy
C0192207|ICD9CM|PT|29.31|Cricopharyngeal myotomy
C0192210|ICD9CM|AB|29.12|Pharyngeal biopsy
C0192210|ICD9CM|PT|29.12|Pharyngeal biopsy
C0192217|ICD9CM|PT|98.13|Removal of intraluminal foreign body from pharynx without incision
C0192217|ICD9CM|AB|98.13|Remov intralum pharyn FB
C0192220|ICD9CM|PT|29.33|Pharyngectomy (partial)
C0192220|ICD9CM|AB|29.33|Pharyngectomy
C0192232|ICD9CM|AB|29.11|Pharyngoscopy
C0192232|ICD9CM|PT|29.11|Pharyngoscopy
C0192243|ICD9CM|PT|29.51|Suture of laceration of pharynx
C0192243|ICD9CM|AB|29.51|Suture of pharyngeal lac
C0192249|ICD9CM|PT|29.54|Lysis of pharyngeal adhesions
C0192249|ICD9CM|AB|29.54|Lysis pharyngeal adhes
C0192256|ICD9CM|PT|29.91|Dilation of pharynx
C0192256|ICD9CM|AB|29.91|Pharyngeal dilation
C0192259|ICD9CM|HT|42|Operations on esophagus
C0192265|ICD9CM|AB|42.7|Esophagomyotomy
C0192265|ICD9CM|PT|42.7|Esophagomyotomy
C0192288|ICD9CM|AB|42.42|Total esophagectomy
C0192288|ICD9CM|PT|42.42|Total esophagectomy
C0192289|ICD9CM|AB|42.41|Partial esophagectomy
C0192289|ICD9CM|PT|42.41|Partial esophagectomy
C0192307|ICD9CM|PT|42.22|Esophagoscopy through artificial stoma
C0192307|ICD9CM|AB|42.22|Esophagoscopy thru stoma
C0192308|ICD9CM|PT|42.24|Closed [endoscopic] biopsy of esophagus
C0192308|ICD9CM|AB|42.24|Closed bx of esophagus
C0192312|ICD9CM|PT|98.02|Removal of intraluminal foreign body from esophagus without incision
C0192312|ICD9CM|AB|98.02|Remov intralum esoph FB
C0192324|ICD9CM|PT|42.85|Repair of esophageal stricture
C0192324|ICD9CM|AB|42.85|Esophag stricture repair
C0192331|ICD9CM|PT|42.91|Ligation of esophageal varices
C0192331|ICD9CM|AB|42.91|Ligation esoph varix
C0192332|ICD9CM|PT|42.55|Intrathoracic esophageal anastomosis with interposition of colon
C0192332|ICD9CM|AB|42.55|Thorac lg bowel interpos
C0192333|ICD9CM|PT|42.58|Intrathoracic esophageal anastomosis with other interposition
C0192333|ICD9CM|AB|42.58|Thorac interposition NEC
C0192336|ICD9CM|PT|42.12|Exteriorization of esophageal pouch
C0192336|ICD9CM|AB|42.12|Esoph pouch exteriorizat
C0192347|ICD9CM|PT|42.83|Closure of esophagostomy
C0192347|ICD9CM|AB|42.83|Esophagostomy closure
C0192353|ICD9CM|PT|42.52|Intrathoracic esophagogastrostomy
C0192353|ICD9CM|AB|42.52|Thorac esophagogastrost
C0192359|ICD9CM|PT|42.53|Intrathoracic esophageal anastomosis with interposition of small bowel
C0192359|ICD9CM|AB|42.53|Thorac sm bowel interpos
C0192401|ICD9CM|AB|43.0|Gastrotomy
C0192401|ICD9CM|PT|43.0|Gastrotomy
C0192421|ICD9CM|PT|44.15|Open biopsy of stomach
C0192421|ICD9CM|AB|44.15|Open gastric biopsy
C0192444|ICD9CM|PT|43.7|Partial gastrectomy with anastomosis to jejunum
C0192444|ICD9CM|AB|43.7|Part gastrec w jej anast
C0192447|ICD9CM|PT|43.91|Total gastrectomy with intestinal interposition
C0192447|ICD9CM|AB|43.91|Tot gast w intes interpo
C0192448|ICD9CM|PT|43.81|Partial gastrectomy with jejunal transposition
C0192448|ICD9CM|AB|43.81|Part gast w jej transpos
C0192456|ICD9CM|AB|96.35|Gastric gavage
C0192456|ICD9CM|PT|96.35|Gastric gavage
C0192457|ICD9CM|PT|44.93|Insertion of gastric bubble (balloon)
C0192457|ICD9CM|AB|44.93|Insert gastric bubble
C0192458|ICD9CM|PT|44.94|Removal of gastric bubble (balloon)
C0192458|ICD9CM|AB|44.94|Remove gastric bubble
C0192461|ICD9CM|PT|97.02|Replacement of gastrostomy tube
C0192461|ICD9CM|AB|97.02|Replace gastrostomy tube
C0192462|ICD9CM|PT|97.51|Removal of gastrostomy tube
C0192462|ICD9CM|AB|97.51|Remov gastrostomy tube
C0192468|ICD9CM|PT|44.11|Transabdominal gastroscopy
C0192468|ICD9CM|AB|44.11|Transabdomin gastroscopy
C0192469|ICD9CM|PT|44.12|Gastroscopy through artificial stoma
C0192469|ICD9CM|AB|44.12|Gastroscopy thru stoma
C0192472|ICD9CM|PT|44.14|Closed [endoscopic] biopsy of stomach
C0192472|ICD9CM|AB|44.14|Closed gastric biopsy
C0192475|ICD9CM|PT|44.22|Endoscopic dilation of pylorus
C0192475|ICD9CM|AB|44.22|Endoscop dilate pylorus
C0192486|ICD9CM|AB|44.65|Esophagogastroplasty
C0192486|ICD9CM|PT|44.65|Esophagogastroplasty
C0192489|ICD9CM|HT|44.2|Pyloroplasty
C0192504|ICD9CM|AB|44.64|Gastropexy
C0192504|ICD9CM|PT|44.64|Gastropexy
C0192543|ICD9CM|PT|44.62|Closure of gastrostomy
C0192543|ICD9CM|AB|44.62|Gastrostomy closure
C0192552|ICD9CM|PT|44.61|Suture of laceration of stomach
C0192552|ICD9CM|AB|44.61|Suture gastric lacerat
C0192557|ICD9CM|PT|44.91|Ligation of gastric varices
C0192557|ICD9CM|AB|44.91|Ligate gastric varices
C0192579|ICD9CM|HT|45.0|Enterotomy
C0192579|ICD9CM|PT|45.00|Incision of intestine, not otherwise specified
C0192579|ICD9CM|AB|45.00|Intestinal incision NOS
C0192584|ICD9CM|PT|45.01|Incision of duodenum
C0192584|ICD9CM|AB|45.01|Duodenal incision
C0192611|ICD9CM|PT|45.15|Open biopsy of small intestine
C0192611|ICD9CM|AB|45.15|Open small bowel biopsy
C0192617|ICD9CM|PT|45.61|Multiple segmental resection of small intestine
C0192617|ICD9CM|AB|45.61|Mult seg sm bowel excis
C0192618|ICD9CM|PT|45.63|Total removal of small intestine
C0192618|ICD9CM|AB|45.63|Total removal sm bowel
C0192620|ICD9CM|PT|46.02|Resection of exteriorized segment of small intestine
C0192620|ICD9CM|AB|46.02|Resect ext seg sm bowel
C0192647|ICD9CM|PT|97.52|Removal of tube from small intestine
C0192647|ICD9CM|AB|97.52|Remov small bowel tube
C0192649|ICD9CM|PT|97.03|Replacement of tube or enterostomy device of small intestine
C0192649|ICD9CM|AB|97.03|Replace small bowel tube
C0192675|ICD9CM|PT|45.14|Closed [endoscopic] biopsy of small intestine
C0192675|ICD9CM|AB|45.14|Clos small bowel biopsy
C0192683|ICD9CM|PT|45.12|Endoscopy of small intestine through artificial stoma
C0192683|ICD9CM|AB|45.12|Endosc sm bowel thru st
C0192708|ICD9CM|HT|46.6|Fixation of intestine
C0192708|ICD9CM|PT|46.60|Fixation of intestine, not otherwise specified
C0192708|ICD9CM|AB|46.60|Intestinal fixation NOS
C0192710|ICD9CM|HT|46.0|Exteriorization of intestine
C0192711|ICD9CM|HT|45.9|Intestinal anastomosis
C0192711|ICD9CM|PT|45.90|Intestinal anastomosis, not otherwise specified
C0192711|ICD9CM|AB|45.90|Intestinal anastom NOS
C0192716|ICD9CM|HT|46.4|Revision of intestinal stoma
C0192716|ICD9CM|PT|46.40|Revision of intestinal stoma, not otherwise specified
C0192716|ICD9CM|AB|46.40|Intest stoma revis NOS
C0192718|ICD9CM|PT|46.24|Delayed opening of ileostomy
C0192718|ICD9CM|AB|46.24|Delay opening ileostomy
C0192719|ICD9CM|HT|46.5|Closure of intestinal stoma
C0192719|ICD9CM|PT|46.50|Closure of intestinal stoma, not otherwise specified
C0192719|ICD9CM|AB|46.50|Intest stoma closure NOS
C0192737|ICD9CM|PT|46.61|Fixation of small intestine to abdominal wall
C0192737|ICD9CM|AB|46.61|Sm bowel-abd wall fixat
C0192741|ICD9CM|PT|45.91|Small-to-small intestinal anastomosis
C0192741|ICD9CM|AB|45.91|Sm-to-sm bowel anastom
C0192745|ICD9CM|PT|45.92|Anastomosis of small intestine to rectal stump
C0192745|ICD9CM|AB|45.92|Sm bowel-rect stump anas
C0192747|ICD9CM|PT|46.93|Revision of anastomosis of small intestine
C0192747|ICD9CM|AB|46.93|Revise sm bowel anastom
C0192757|ICD9CM|PT|46.51|Closure of stoma of small intestine
C0192757|ICD9CM|AB|46.51|Sm bowel stoma closure
C0192758|ICD9CM|AB|46.72|Duodenal fistula closure
C0192758|ICD9CM|PT|46.72|Closure of fistula of duodenum
C0192764|ICD9CM|PT|44.42|Suture of duodenal ulcer site
C0192764|ICD9CM|AB|44.42|Suture duoden ulcer site
C0192770|ICD9CM|PT|46.41|Revision of stoma of small intestine
C0192770|ICD9CM|AB|46.41|Sm bowel stoma revision
C0192800|ICD9CM|PT|46.80|Intra-abdominal manipulation of intestine, not otherwise specified
C0192800|ICD9CM|AB|46.80|Intra-ab bowel manip NOS
C0192801|ICD9CM|PT|46.81|Intra-abdominal manipulation of small intestine
C0192801|ICD9CM|AB|46.81|Intra-abd sm bowel manip
C0192810|ICD9CM|PT|96.24|Dilation and manipulation of enterostomy stoma
C0192810|ICD9CM|AB|96.24|Dilat enterostomy stoma
C0192819|ICD9CM|HT|47|Operations on appendix
C0192822|ICD9CM|PT|45.03|Incision of large intestine
C0192822|ICD9CM|AB|45.03|Large bowel incision
C0192837|ICD9CM|PT|46.04|Resection of exteriorized segment of large intestine
C0192837|ICD9CM|AB|46.04|Resect ext seg lg bowel
C0192840|ICD9CM|PT|45.26|Open biopsy of large intestine
C0192840|ICD9CM|AB|45.26|Open large bowel biopsy
C0192882|ICD9CM|HT|47.1|Incidental appendectomy
C0192888|ICD9CM|PT|97.04|Replacement of tube or enterostomy device of large intestine
C0192888|ICD9CM|AB|97.04|Replace large bowel tube
C0192891|ICD9CM|PT|45.25|Closed [endoscopic] biopsy of large intestine
C0192891|ICD9CM|AB|45.25|Clos large bowel biopsy
C0192894|ICD9CM|PT|45.42|Endoscopic polypectomy of large intestine
C0192894|ICD9CM|AB|45.42|Endo polpectomy lrge int
C0192896|ICD9CM|PT|98.04|Removal of intraluminal foreign body from large intestine without incision
C0192896|ICD9CM|AB|98.04|Remov intralum colon FB
C0192897|ICD9CM|PT|45.22|Endoscopy of large intestine through artificial stoma
C0192897|ICD9CM|AB|45.22|Endosc lg bowel thru st
C0192928|ICD9CM|PT|48.22|Proctosigmoidoscopy through artificial stoma
C0192928|ICD9CM|AB|48.22|Proctosigmoidosc thru st
C0192943|ICD9CM|PT|46.63|Fixation of large intestine to abdominal wall
C0192943|ICD9CM|AB|46.63|Lg bowel-abd wall fixat
C0192952|ICD9CM|PT|46.03|Exteriorization of large intestine
C0192952|ICD9CM|AB|46.03|Lg bowel exteriorization
C0192953|ICD9CM|AB|47.91|Appendicostomy
C0192953|ICD9CM|PT|47.91|Appendicostomy
C0192955|ICD9CM|PT|45.94|Large-to-large intestinal anastomosis
C0192955|ICD9CM|AB|45.94|Lg-to-lg bowel anastom
C0192960|ICD9CM|PT|46.94|Revision of anastomosis of large intestine
C0192960|ICD9CM|AB|46.94|Revise lg bowel anastom
C0192971|ICD9CM|AB|46.11|Temporary colostomy
C0192971|ICD9CM|PT|46.11|Temporary colostomy
C0192973|ICD9CM|AB|46.13|Permanent colostomy
C0192973|ICD9CM|PT|46.13|Permanent colostomy
C0192976|ICD9CM|PT|46.76|Closure of fistula of large intestine
C0192976|ICD9CM|AB|46.76|Close lg bowel fistula
C0192980|ICD9CM|PT|46.52|Closure of stoma of large intestine
C0192980|ICD9CM|AB|46.52|Lg bowel stoma closure
C0192983|ICD9CM|PT|47.92|Closure of appendiceal fistula
C0192983|ICD9CM|AB|47.92|Close appendiceal fistul
C0192991|ICD9CM|PT|46.14|Delayed opening of colostomy
C0192991|ICD9CM|AB|46.14|Delay opening colostomy
C0192992|ICD9CM|PT|46.42|Repair of pericolostomy hernia
C0192992|ICD9CM|AB|46.42|Pericolost hernia repair
C0193004|ICD9CM|PT|46.82|Intra-abdominal manipulation of large intestine
C0193004|ICD9CM|AB|46.82|Intra-abd lg bowel manip
C0193014|ICD9CM|HT|49|Operations on anus
C0193017|ICD9CM|AB|48.0|Proctotomy
C0193017|ICD9CM|PT|48.0|Proctotomy
C0193019|ICD9CM|PT|48.91|Incision of rectal stricture
C0193019|ICD9CM|AB|48.91|Incis rectal stricture
C0193020|ICD9CM|PT|48.81|Incision of perirectal tissue
C0193020|ICD9CM|AB|48.81|Perirectal incision
C0193037|ICD9CM|PT|49.51|Left lateral anal sphincterotomy
C0193037|ICD9CM|AB|49.51|Left lat sphincterotomy
C0193042|ICD9CM|AB|49.11|Anal fistulotomy
C0193042|ICD9CM|PT|49.11|Anal fistulotomy
C0193047|ICD9CM|PT|49.47|Evacuation of thrombosed hemorrhoids
C0193047|ICD9CM|AB|49.47|Hemorrhoid evacuation
C0193056|ICD9CM|PT|48.92|Anorectal myectomy
C0193056|ICD9CM|AB|48.92|Anorectal myomectomy
C0193082|ICD9CM|PT|48.61|Transsacral rectosigmoidectomy
C0193082|ICD9CM|AB|48.61|Transsac rectosigmoidect
C0193085|ICD9CM|PT|48.64|Posterior resection of rectum
C0193085|ICD9CM|AB|48.64|Posterior rect resection
C0193101|ICD9CM|PT|49.45|Ligation of hemorrhoids
C0193101|ICD9CM|AB|49.45|Hemorrhoid ligation
C0193114|ICD9CM|PT|49.23|Biopsy of anus
C0193114|ICD9CM|AB|49.23|Anal biopsy
C0193115|ICD9CM|PT|49.22|Biopsy of perianal tissue
C0193115|ICD9CM|AB|49.22|Perianal biopsy
C0193125|ICD9CM|AB|49.12|Anal fistulectomy
C0193125|ICD9CM|PT|49.12|Anal fistulectomy
C0193134|ICD9CM|PT|49.03|Excision of perianal skin tags
C0193134|ICD9CM|AB|49.03|Excis perianal skin tag
C0193144|ICD9CM|AB|96.37|Proctoclysis
C0193144|ICD9CM|PT|96.37|Proctoclysis
C0193147|ICD9CM|AB|96.19|Rectal packing
C0193147|ICD9CM|PT|96.19|Rectal packing
C0193149|ICD9CM|PT|49.92|Insertion of subcutaneous electrical anal stimulator
C0193149|ICD9CM|AB|49.92|Insert subq anal stimul
C0193156|ICD9CM|PT|48.24|Closed [endoscopic] biopsy of rectum
C0193156|ICD9CM|AB|48.24|Closed rectal biopsy
C0193158|ICD9CM|AB|49.21|Anoscopy
C0193158|ICD9CM|PT|49.21|Anoscopy
C0193171|ICD9CM|AB|48.74|Rectorectostomy
C0193171|ICD9CM|PT|48.74|Rectorectostomy
C0193184|ICD9CM|AB|48.1|Proctostomy
C0193184|ICD9CM|PT|48.1|Proctostomy
C0193186|ICD9CM|AB|48.72|Closure of proctostomy
C0193186|ICD9CM|PT|48.72|Closure of proctostomy
C0193187|ICD9CM|PT|48.71|Suture of laceration of rectum
C0193187|ICD9CM|AB|48.71|Suture of rectal lacer
C0193189|ICD9CM|PT|48.93|Repair of perirectal fistula
C0193189|ICD9CM|AB|48.93|Repair perirect fistula
C0193192|ICD9CM|AB|49.73|Closure of anal fistula
C0193192|ICD9CM|PT|49.73|Closure of anal fistula
C0193200|ICD9CM|HT|49.7|Repair of anus
C0193206|ICD9CM|PT|49.71|Suture of laceration of anus
C0193206|ICD9CM|AB|49.71|Suture anal laceration
C0193210|ICD9CM|AB|49.72|Anal cerclage
C0193210|ICD9CM|PT|49.72|Anal cerclage
C0193219|ICD9CM|PT|49.74|Gracilis muscle transplant for anal incontinence
C0193219|ICD9CM|AB|49.74|Gracilis musc transplan
C0193247|ICD9CM|PT|49.44|Destruction of hemorrhoids by cryotherapy
C0193247|ICD9CM|AB|49.44|Hemorrhoid cryotherapy
C0193248|ICD9CM|PT|49.43|Cauterization of hemorrhoids
C0193248|ICD9CM|AB|49.43|Hemorrhoid cauterizat
C0193249|ICD9CM|PT|49.42|Injection of hemorrhoids
C0193249|ICD9CM|AB|49.42|Hemorrhoid injection
C0193264|ICD9CM|AB|96.22|Dilation of rectum
C0193264|ICD9CM|PT|96.22|Dilation of rectum
C0193268|ICD9CM|PT|99.93|Rectal massage (for levator spasm)
C0193268|ICD9CM|AB|99.93|Rectal massage
C0193270|ICD9CM|PT|96.26|Manual reduction of rectal prolapse
C0193270|ICD9CM|AB|96.26|Manual reduc rect prolap
C0193305|ICD9CM|HT|26.2|Excision of lesion of salivary gland
C0193311|ICD9CM|HT|26.3|Sialoadenectomy
C0193311|ICD9CM|AB|26.30|Sialoadenectomy NOS
C0193311|ICD9CM|PT|26.30|Sialoadenectomy, not otherwise specified
C0193312|ICD9CM|AB|26.31|Partial sialoadenectomy
C0193312|ICD9CM|PT|26.31|Partial sialoadenectomy
C0193313|ICD9CM|AB|26.32|Complete sialoadenectomy
C0193313|ICD9CM|PT|26.32|Complete sialoadenectomy
C0193344|ICD9CM|PT|26.21|Marsupialization of salivary gland cyst
C0193344|ICD9CM|AB|26.21|Salivary cyst marsupial
C0193348|ICD9CM|PT|26.41|Suture of laceration of salivary gland
C0193348|ICD9CM|AB|26.41|Suture of saliv glnd lac
C0193349|ICD9CM|PT|26.42|Closure of salivary fistula
C0193349|ICD9CM|AB|26.42|Salivary fistula closure
C0193369|ICD9CM|PT|26.91|Probing of salivary duct
C0193369|ICD9CM|AB|26.91|Salivary duct probing
C0193373|ICD9CM|HT|50|Operations on liver
C0193374|ICD9CM|HT|50.1|Diagnostic procedures on liver
C0193377|ICD9CM|AB|50.0|Hepatotomy
C0193377|ICD9CM|PT|50.0|Hepatotomy
C0193384|ICD9CM|PT|50.91|Percutaneous aspiration of liver
C0193384|ICD9CM|AB|50.91|Percutan liver aspirat
C0193389|ICD9CM|PT|50.12|Open biopsy of liver
C0193389|ICD9CM|AB|50.12|Open liver biopsy
C0193398|ICD9CM|AB|50.22|Partial hepatectomy
C0193398|ICD9CM|PT|50.22|Partial hepatectomy
C0193399|ICD9CM|PT|50.3|Lobectomy of liver
C0193399|ICD9CM|AB|50.3|Hepatic lobectomy
C0193436|ICD9CM|HT|51|Operations on gallbladder and biliary tract
C0193444|ICD9CM|PT|51.01|Percutaneous aspiration of gallbladder
C0193444|ICD9CM|AB|51.01|Percutan aspiration gb
C0193470|ICD9CM|PT|51.96|Percutaneous extraction of common duct stones
C0193470|ICD9CM|AB|51.96|Perc extrac com duc calc
C0193480|ICD9CM|PT|51.61|Excision of cystic duct remnant
C0193480|ICD9CM|AB|51.61|Excis cyst duct remnant
C0193483|ICD9CM|PT|51.62|Excision of ampulla of Vater (with reimplantation of common duct)
C0193483|ICD9CM|AB|51.62|Excis ampulla of vater
C0193491|ICD9CM|PT|51.43|Insertion of choledochohepatic tube for decompression
C0193491|ICD9CM|AB|51.43|Choledochohepat intubat
C0193496|ICD9CM|PT|51.95|Removal of prosthetic device from bile duct
C0193496|ICD9CM|AB|51.95|Remove bile duct prosth
C0193498|ICD9CM|PT|97.54|Removal of cholecystostomy tube
C0193498|ICD9CM|AB|97.54|Remov cholecystost tube
C0193504|ICD9CM|PT|51.11|Endoscopic retrograde cholangiography [ERC]
C0193504|ICD9CM|AB|51.11|Endosc retro cholangio
C0193530|ICD9CM|PT|51.31|Anastomosis of gallbladder to hepatic ducts
C0193530|ICD9CM|AB|51.31|Gb-to-hepat duct anast
C0193531|ICD9CM|PT|51.37|Anastomosis of hepatic duct to gastrointestinal tract
C0193531|ICD9CM|AB|51.37|Hepatic duct-gi anastom
C0193543|ICD9CM|PT|51.94|Revision of anastomosis of biliary tract
C0193543|ICD9CM|AB|51.94|Revis bile tract anastom
C0193544|ICD9CM|PT|51.32|Anastomosis of gallbladder to intestine
C0193544|ICD9CM|AB|51.32|Gb-to-intestine anastom
C0193546|ICD9CM|PT|51.34|Anastomosis of gallbladder to stomach
C0193546|ICD9CM|AB|51.34|Gb-to-stomach anastomos
C0193547|ICD9CM|PT|51.33|Anastomosis of gallbladder to pancreas
C0193547|ICD9CM|AB|51.33|Gb-to-pancreas anastom
C0193558|ICD9CM|AB|51.36|Choledochoenterostomy
C0193558|ICD9CM|PT|51.36|Choledochoenterostomy
C0193561|ICD9CM|PT|51.92|Closure of cholecystostomy
C0193561|ICD9CM|AB|51.92|Closure cholecystostomy
C0193566|ICD9CM|HT|51.7|Repair of bile ducts
C0193591|ICD9CM|PT|51.81|Dilation of sphincter of Oddi
C0193591|ICD9CM|AB|51.81|Sphincter of oddi dilat
C0193594|ICD9CM|HT|52|Operations on pancreas
C0193596|ICD9CM|HT|52.0|Pancreatotomy
C0193599|ICD9CM|PT|52.4|Internal drainage of pancreatic cyst
C0193599|ICD9CM|AB|52.4|Int drain pancreat cyst
C0193607|ICD9CM|PT|52.12|Open biopsy of pancreas
C0193607|ICD9CM|AB|52.12|Open pancreatic biopsy
C0193612|ICD9CM|PT|52.7|Radical pancreaticoduodenectomy
C0193612|ICD9CM|AB|52.7|Rad pancreaticoduodenect
C0193625|ICD9CM|PT|96.42|Irrigation of pancreatic tube
C0193625|ICD9CM|AB|96.42|Pancreatic tube irrigat
C0193634|ICD9CM|PT|52.98|Endoscopic dilation of pancreatic duct
C0193634|ICD9CM|AB|52.98|Endosc dil pancreat duct
C0193635|ICD9CM|PT|52.97|Endoscopic insertion of nasopancreatic drainage tube
C0193635|ICD9CM|AB|52.97|Endosc inser nasopan tub
C0193637|ICD9CM|PT|52.94|Endoscopic removal of stone(s) from pancreatic duct
C0193637|ICD9CM|AB|52.94|Endosc remove panc stone
C0193648|ICD9CM|PT|52.3|Marsupialization of pancreatic cyst
C0193648|ICD9CM|AB|52.3|Pancreat cyst marsupiali
C0193657|ICD9CM|PT|52.82|Homotransplant of pancreas
C0193657|ICD9CM|AB|52.82|Pancreatic homotransplan
C0193658|ICD9CM|PT|52.83|Heterotransplant of pancreas
C0193658|ICD9CM|AB|52.83|Pancreatic heterotranspl
C0193669|ICD9CM|HT|07.5|Operations on pineal gland
C0193676|ICD9CM|PT|07.41|Incision of adrenal gland
C0193676|ICD9CM|AB|07.41|Adrenal incision
C0193679|ICD9CM|PT|07.02|Bilateral exploration of adrenal field
C0193679|ICD9CM|AB|07.02|Bilat adrenal explorat
C0193682|ICD9CM|PT|07.72|Incision of pituitary gland
C0193682|ICD9CM|AB|07.72|Pituitary gland incision
C0193689|ICD9CM|PT|07.52|Incision of pineal gland
C0193689|ICD9CM|AB|07.52|Pineal gland incision
C0193694|ICD9CM|PT|06.13|Biopsy of parathyroid gland
C0193694|ICD9CM|AB|06.13|Parathyroid biopsy
C0193696|ICD9CM|PT|06.81|Complete parathyroidectomy
C0193696|ICD9CM|AB|06.81|Total parathyroidectomy
C0193702|ICD9CM|PT|07.21|Excision of lesion of adrenal gland
C0193702|ICD9CM|AB|07.21|Adrenal lesion excision
C0193704|ICD9CM|AB|07.3|Bilateral adrenalectomy
C0193704|ICD9CM|PT|07.3|Bilateral adrenalectomy
C0193725|ICD9CM|PT|07.61|Partial excision of pituitary gland, transfrontal approach
C0193725|ICD9CM|AB|07.61|Exc pituit les-transfron
C0193726|ICD9CM|PT|07.62|Partial excision of pituitary gland, transsphenoidal approach
C0193726|ICD9CM|AB|07.62|Exc pituit les-transphen
C0193727|ICD9CM|PT|07.63|Partial excision of pituitary gland, unspecified approach
C0193727|ICD9CM|AB|07.63|Part excis pituitary NOS
C0193728|ICD9CM|PT|07.64|Total excision of pituitary gland, transfrontal approach
C0193728|ICD9CM|AB|07.64|Tot exc pituit-transfron
C0193729|ICD9CM|PT|07.65|Total excision of pituitary gland, transsphenoidal approach
C0193729|ICD9CM|AB|07.65|Tot exc pituit-transphen
C0193734|ICD9CM|PT|07.53|Partial excision of pineal gland
C0193734|ICD9CM|AB|07.53|Partial pinealectomy
C0193735|ICD9CM|PT|07.54|Total excision of pineal gland
C0193735|ICD9CM|AB|07.54|Total pinealectomy
C0193745|ICD9CM|PT|07.44|Repair of adrenal gland
C0193745|ICD9CM|AB|07.44|Adrenal repair
C0193774|ICD9CM|PT|06.02|Reopening of wound of thyroid field
C0193774|ICD9CM|AB|06.02|Reopen thyroid field wnd
C0193775|ICD9CM|PT|06.01|Aspiration of thyroid field
C0193775|ICD9CM|AB|06.01|Thyroid field aspiration
C0193777|ICD9CM|PT|06.91|Division of thyroid isthmus
C0193777|ICD9CM|AB|06.91|Thyroid isthmus division
C0193782|ICD9CM|PT|06.31|Excision of lesion of thyroid
C0193782|ICD9CM|AB|06.31|Excision thyroid lesion
C0193788|ICD9CM|AB|06.4|Complete thyroidectomy
C0193788|ICD9CM|PT|06.4|Complete thyroidectomy
C0193794|ICD9CM|PT|06.52|Complete substernal thyroidectomy
C0193794|ICD9CM|AB|06.52|Tot substern thyroidect
C0193795|ICD9CM|PT|06.51|Partial substernal thyroidectomy
C0193795|ICD9CM|AB|06.51|Part substern thyroidect
C0193805|ICD9CM|PT|06.6|Excision of lingual thyroid
C0193805|ICD9CM|AB|06.6|Lingual thyroid excision
C0193818|ICD9CM|PT|06.93|Suture of thyroid gland
C0193818|ICD9CM|AB|06.93|Thyroid suture
C0193823|ICD9CM|PT|06.94|Thyroid tissue reimplantation
C0193823|ICD9CM|AB|06.94|Thyroid reimplantation
C0193831|ICD9CM|HT|40.6|Operations on thoracic duct
C0193843|ICD9CM|PT|40.11|Biopsy of lymphatic structure
C0193843|ICD9CM|AB|40.11|Lymphatic struct biopsy
C0193854|ICD9CM|PT|40.50|Radical excision of lymph nodes, not otherwise specified
C0193854|ICD9CM|AB|40.50|Rad node dissection NOS
C0193857|ICD9CM|PT|40.21|Excision of deep cervical lymph node
C0193857|ICD9CM|AB|40.21|Excis deep cervical node
C0193862|ICD9CM|PT|40.41|Radical neck dissection, unilateral
C0193862|ICD9CM|AB|40.41|Unilat rad neck dissect
C0193863|ICD9CM|PT|40.42|Radical neck dissection, bilateral
C0193863|ICD9CM|AB|40.42|Bilat rad neck dissect
C0193867|ICD9CM|PT|40.23|Excision of axillary lymph node
C0193867|ICD9CM|AB|40.23|Excise axillary node
C0193871|ICD9CM|PT|40.22|Excision of internal mammary lymph node
C0193871|ICD9CM|AB|40.22|Excise int mammary node
C0193880|ICD9CM|PT|40.53|Radical excision of iliac lymph nodes
C0193880|ICD9CM|AB|40.53|Rad dissect iliac nodes
C0193884|ICD9CM|PT|40.24|Excision of inguinal lymph node
C0193884|ICD9CM|AB|40.24|Excise inguinal node
C0193888|ICD9CM|AB|40.54|Radical groin dissection
C0193888|ICD9CM|PT|40.54|Radical groin dissection
C0193891|ICD9CM|PT|40.61|Cannulation of thoracic duct
C0193891|ICD9CM|AB|40.61|Thorac duct cannulation
C0193902|ICD9CM|PT|40.62|Fistulization of thoracic duct
C0193902|ICD9CM|AB|40.62|Thoracic duct fistulizat
C0193903|ICD9CM|PT|40.63|Closure of fistula of thoracic duct
C0193903|ICD9CM|AB|40.63|Close thoracic duct fist
C0193907|ICD9CM|PT|40.64|Ligation of thoracic duct
C0193907|ICD9CM|AB|40.64|Ligate thoracic duct
C0193926|ICD9CM|PT|28.7|Control of hemorrhage after tonsillectomy and adenoidectomy
C0193926|ICD9CM|AB|28.7|Hemorr contrl post T & A
C0193940|ICD9CM|AB|28.4|Excision of tonsil tag
C0193940|ICD9CM|PT|28.4|Excision of tonsil tag
C0193941|ICD9CM|PT|28.5|Excision of lingual tonsil
C0193941|ICD9CM|AB|28.5|Excision lingual tonsil
C0193959|ICD9CM|PT|28.3|Tonsillectomy with adenoidectomy
C0193959|ICD9CM|AB|28.3|Tonsillectomy/adenoidec
C0193987|ICD9CM|AB|41.2|Splenotomy
C0193987|ICD9CM|PT|41.2|Splenotomy
C0193995|ICD9CM|PT|41.42|Excision of lesion or tissue of spleen
C0193995|ICD9CM|AB|41.42|Exc splenic lesion/tiss
C0193997|ICD9CM|AB|41.43|Partial splenectomy
C0193997|ICD9CM|PT|41.43|Partial splenectomy
C0193998|ICD9CM|PT|41.93|Excision of accessory spleen
C0193998|ICD9CM|AB|41.93|Exc of accessory spleen
C0194001|ICD9CM|PT|07.16|Biopsy of thymus
C0194001|ICD9CM|AB|07.16|Thymus biopsy
C0194015|ICD9CM|PT|41.91|Aspiration of bone marrow from donor for transplant
C0194015|ICD9CM|AB|41.91|Donor marrow aspiration
C0194018|ICD9CM|PT|41.92|Injection into bone marrow
C0194018|ICD9CM|AB|41.92|Injection into marrow
C0194026|ICD9CM|PT|41.41|Marsupialization of splenic cyst
C0194026|ICD9CM|AB|41.41|Splenic cyst marsupial
C0194028|ICD9CM|AB|07.93|Repair of thymus
C0194028|ICD9CM|PT|07.93|Repair of thymus
C0194034|ICD9CM|PT|41.94|Transplantation of spleen
C0194034|ICD9CM|AB|41.94|Spleen transplantation
C0194035|ICD9CM|AB|07.94|Thymus transplantation
C0194035|ICD9CM|PT|07.94|Transplantation of thymus
C0194039|ICD9CM|PT|41.01|Autologous bone marrow transplant without purging
C0194039|ICD9CM|AB|41.01|Auto bone mt w/o purg
C0194053|ICD9CM|HT|55|Operations on kidney
C0194056|ICD9CM|AB|55.01|Nephrotomy
C0194056|ICD9CM|PT|55.01|Nephrotomy
C0194061|ICD9CM|PT|55.92|Percutaneous aspiration of kidney (pelvis)
C0194061|ICD9CM|AB|55.92|Percutan renal aspirat
C0194063|ICD9CM|AB|55.11|Pyelotomy
C0194063|ICD9CM|PT|55.11|Pyelotomy
C0194074|ICD9CM|PT|55.24|Open biopsy of kidney
C0194074|ICD9CM|AB|55.24|Open renal biopsy
C0194084|ICD9CM|AB|55.54|Bilateral nephrectomy
C0194084|ICD9CM|PT|55.54|Bilateral nephrectomy
C0194085|ICD9CM|PT|55.52|Nephrectomy of remaining kidney
C0194085|ICD9CM|AB|55.52|Solitary kidney nephrect
C0194086|ICD9CM|AB|55.4|Partial nephrectomy
C0194086|ICD9CM|PT|55.4|Partial nephrectomy
C0194089|ICD9CM|PT|55.91|Decapsulation of kidney
C0194089|ICD9CM|AB|55.91|Renal decapsulation
C0194121|ICD9CM|AB|55.12|Pyelostomy
C0194121|ICD9CM|PT|55.12|Pyelostomy
C0194127|ICD9CM|PT|55.93|Replacement of nephrostomy tube
C0194127|ICD9CM|AB|55.93|Replace nephrostomy tube
C0194129|ICD9CM|PT|55.94|Replacement of pyelostomy tube
C0194129|ICD9CM|AB|55.94|Replace pyelostomy tube
C0194130|ICD9CM|PT|97.61|Removal of pyelostomy and nephrostomy tube
C0194130|ICD9CM|AB|97.61|Remov pyelos/nephros tub
C0194133|ICD9CM|PT|55.95|Local perfusion of kidney
C0194133|ICD9CM|AB|55.95|Local renal perfusion
C0194135|ICD9CM|AB|55.21|Nephroscopy
C0194135|ICD9CM|PT|55.21|Nephroscopy
C0194159|ICD9CM|AB|55.7|Nephropexy
C0194159|ICD9CM|PT|55.7|Nephropexy
C0194194|ICD9CM|PT|55.61|Renal autotransplantation
C0194194|ICD9CM|AB|55.61|Renal autotransplant
C0194203|ICD9CM|PT|55.98|Removal of mechanical kidney
C0194203|ICD9CM|AB|55.98|Remov mechanical kidney
C0194204|ICD9CM|PT|39.55|Reimplantation of aberrant renal vessel
C0194204|ICD9CM|AB|39.55|Reimplan aberr renal ves
C0194206|ICD9CM|PT|55.84|Reduction of torsion of renal pedicle
C0194206|ICD9CM|AB|55.84|Reduce renal pedicl tors
C0194209|ICD9CM|HT|56|Operations on ureter
C0194211|ICD9CM|AB|56.2|Ureterotomy
C0194211|ICD9CM|PT|56.2|Ureterotomy
C0194224|ICD9CM|HT|56.4|Ureterectomy
C0194224|ICD9CM|AB|56.40|Ureterectomy NOS
C0194224|ICD9CM|PT|56.40|Ureterectomy, not otherwise specified
C0194225|ICD9CM|AB|56.42|Total ureterectomy
C0194225|ICD9CM|PT|56.42|Total ureterectomy
C0194239|ICD9CM|PT|96.46|Irrigation of ureterostomy and ureteral catheter
C0194239|ICD9CM|AB|96.46|Urterost/urete cth irrig
C0194251|ICD9CM|PT|59.93|Replacement of ureterostomy tube
C0194251|ICD9CM|AB|59.93|Replace ureterost tube
C0194252|ICD9CM|PT|56.92|Implantation of electronic ureteral stimulator
C0194252|ICD9CM|AB|56.92|Implant ureteral stimul
C0194253|ICD9CM|PT|56.94|Removal of electronic ureteral stimulator
C0194253|ICD9CM|AB|56.94|Remove ureteral stimulat
C0194254|ICD9CM|PT|56.93|Replacement of electronic ureteral stimulator
C0194254|ICD9CM|AB|56.93|Replace ureteral stimul
C0194258|ICD9CM|PT|97.62|Removal of ureterostomy tube and ureteral catheter
C0194258|ICD9CM|AB|97.62|Remov ureteral drain
C0194261|ICD9CM|AB|56.31|Ureteroscopy
C0194261|ICD9CM|PT|56.31|Ureteroscopy
C0194271|ICD9CM|PT|56.0|Transurethral removal of obstruction from ureter and renal pelvis
C0194271|ICD9CM|AB|56.0|Tu remov ureter obstruct
C0194298|ICD9CM|PT|56.35|Endoscopy (cystoscopy) (looposcopy) of ileal conduit
C0194298|ICD9CM|AB|56.35|Endoscopic ileal conduit
C0194300|ICD9CM|AB|56.95|Ligation of ureter
C0194300|ICD9CM|PT|56.95|Ligation of ureter
C0194303|ICD9CM|AB|56.85|Ureteropexy
C0194303|ICD9CM|PT|56.85|Ureteropexy
C0194306|ICD9CM|AB|56.75|Transureteroureterostomy
C0194306|ICD9CM|PT|56.75|Transureteroureterostomy
C0194307|ICD9CM|AB|56.74|Ureteroneocystostomy
C0194307|ICD9CM|PT|56.74|Ureteroneocystostomy
C0194316|ICD9CM|PT|56.83|Closure of ureterostomy
C0194316|ICD9CM|AB|56.83|Ureterostomy closure
C0194328|ICD9CM|PT|56.71|Urinary diversion to intestine
C0194328|ICD9CM|AB|56.71|Urin diversion to bowel
C0194331|ICD9CM|PT|56.52|Revision of cutaneous uretero-ileostomy
C0194331|ICD9CM|AB|56.52|Revis cutan ileoureteros
C0194336|ICD9CM|PT|56.72|Revision of ureterointestinal anastomosis
C0194336|ICD9CM|AB|56.72|Revis ureteroenterostomy
C0194346|ICD9CM|PT|56.81|Lysis of intraluminal adhesions of ureter
C0194346|ICD9CM|AB|56.81|Intralum urete adhesioly
C0194355|ICD9CM|PT|56.91|Dilation of ureteral meatus
C0194355|ICD9CM|AB|56.91|Ureteral meatus dilation
C0194364|ICD9CM|PT|57.93|Control of (postoperative) hemorrhage of bladder
C0194364|ICD9CM|AB|57.93|Control bladd hemorrhage
C0194373|ICD9CM|HT|59.1|Incision of perivesical tissue
C0194396|ICD9CM|AB|57.6|Partial cystectomy
C0194396|ICD9CM|PT|57.6|Partial cystectomy
C0194401|ICD9CM|HT|57.7|Total cystectomy
C0194401|ICD9CM|AB|57.71|Radical cystectomy
C0194401|ICD9CM|PT|57.71|Radical cystectomy
C0194419|ICD9CM|PT|59.94|Replacement of cystostomy tube
C0194419|ICD9CM|AB|59.94|Replace cystostomy tube
C0194424|ICD9CM|PT|96.47|Irrigation of cystostomy
C0194424|ICD9CM|AB|96.47|Cystostomy irrigation
C0194429|ICD9CM|PT|58.93|Implantation of artificial urinary sphincter [AUS]
C0194429|ICD9CM|AB|58.93|Implt artf urin sphinct
C0194432|ICD9CM|PT|57.98|Removal of electronic bladder stimulator
C0194432|ICD9CM|AB|57.98|Remove bladder stimulat
C0194479|ICD9CM|AB|57.85|Cystourethroplasty
C0194479|ICD9CM|PT|57.85|Cystourethroplasty and plastic repair of bladder neck
C0194483|ICD9CM|PT|57.83|Repair of fistula involving bladder and intestine
C0194483|ICD9CM|AB|57.83|Enterovesico fist repair
C0194503|ICD9CM|PT|59.4|Suprapubic sling operation
C0194503|ICD9CM|AB|59.4|Suprapubic sling op
C0194512|ICD9CM|PT|59.71|Levator muscle operation for urethrovesical suspension
C0194512|ICD9CM|AB|59.71|Levator musc suspension
C0194520|ICD9CM|PT|57.87|Reconstruction of urinary bladder
C0194520|ICD9CM|AB|57.87|Bladder reconstruction
C0194522|ICD9CM|PT|57.82|Closure of cystostomy
C0194522|ICD9CM|AB|57.82|Cystostomy closure
C0194523|ICD9CM|PT|57.86|Repair of bladder exstrophy
C0194523|ICD9CM|AB|57.86|Bladder exstrophy repair
C0194542|ICD9CM|PT|57.92|Dilation of bladder neck
C0194542|ICD9CM|AB|57.92|Bladder neck dilation
C0194546|ICD9CM|HT|58|Operations on urethra
C0194550|ICD9CM|AB|58.0|Urethrotomy
C0194550|ICD9CM|PT|58.0|Urethrotomy
C0194552|ICD9CM|PT|58.5|Release of urethral stricture
C0194552|ICD9CM|AB|58.5|Ureth stricture release
C0194553|ICD9CM|PT|58.91|Incision of periurethral tissue
C0194553|ICD9CM|AB|58.91|Periurethral incision
C0194558|ICD9CM|AB|58.1|Urethral meatotomy
C0194558|ICD9CM|PT|58.1|Urethral meatotomy
C0194564|ICD9CM|PT|58.23|Biopsy of urethra
C0194564|ICD9CM|AB|58.23|Urethral biopsy
C0194574|ICD9CM|PT|58.24|Biopsy of periurethral tissue
C0194574|ICD9CM|AB|58.24|Periurethral biopsy
C0194592|ICD9CM|PT|97.65|Removal of urethral stent
C0194592|ICD9CM|AB|97.65|Remov urethral stent
C0194603|ICD9CM|AB|58.21|Perineal urethroscopy
C0194603|ICD9CM|PT|58.21|Perineal urethroscopy
C0194611|ICD9CM|AB|58.42|Urethrostomy closure
C0194611|ICD9CM|PT|58.42|Closure of urethrostomy
C0194633|ICD9CM|AB|58.47|Urethral meatoplasty
C0194633|ICD9CM|PT|58.47|Urethral meatoplasty
C0194639|ICD9CM|PT|59.3|Plication of urethrovesical junction
C0194639|ICD9CM|AB|59.3|Urethroves junct plicat
C0194643|ICD9CM|PT|58.44|Reanastomosis of urethra
C0194643|ICD9CM|AB|58.44|Urethral reanastomosis
C0194648|ICD9CM|AB|59.6|Paraurethral suspension
C0194648|ICD9CM|PT|59.6|Paraurethral suspension
C0194664|ICD9CM|PT|58.6|Dilation of urethra
C0194664|ICD9CM|AB|58.6|Urethral dilation
C0194675|ICD9CM|HT|60-64.99|OPERATIONS ON THE MALE GENITAL ORGANS
C0194682|ICD9CM|HT|64|Operations on penis
C0194684|ICD9CM|AB|64.92|Incision of penis
C0194684|ICD9CM|PT|64.92|Incision of penis
C0194708|ICD9CM|AB|64.3|Amputation of penis
C0194708|ICD9CM|PT|64.3|Amputation of penis
C0194718|ICD9CM|PT|64.94|Fitting of external prosthesis of penis
C0194718|ICD9CM|AB|64.94|Fit ext penile prosthes
C0194742|ICD9CM|PT|64.41|Suture of laceration of penis
C0194742|ICD9CM|AB|64.41|Suture penile laceration
C0194750|ICD9CM|AB|64.45|Replantation of penis
C0194750|ICD9CM|PT|64.45|Replantation of penis
C0194792|ICD9CM|AB|60.0|Incision of prostate
C0194792|ICD9CM|PT|60.0|Incision of prostate
C0194801|ICD9CM|PT|60.81|Incision of periprostatic tissue
C0194801|ICD9CM|AB|60.81|Periprostatic incision
C0194810|ICD9CM|AB|60.5|Radical prostatectomy
C0194810|ICD9CM|PT|60.5|Radical prostatectomy
C0194818|ICD9CM|AB|60.62|Perineal prostatectomy
C0194818|ICD9CM|PT|60.62|Perineal prostatectomy
C0194823|ICD9CM|AB|60.4|Retropubic prostatectomy
C0194823|ICD9CM|PT|60.4|Retropubic prostatectomy
C0194828|ICD9CM|AB|60.3|Suprapubic prostatectomy
C0194828|ICD9CM|PT|60.3|Suprapubic prostatectomy
C0194835|ICD9CM|AB|60.92|Injection into prostate
C0194835|ICD9CM|PT|60.92|Injection into prostate
C0194842|ICD9CM|AB|60.93|Repair of prostate
C0194842|ICD9CM|PT|60.93|Repair of prostate
C0194852|ICD9CM|AB|99.94|Prostatic massage
C0194852|ICD9CM|PT|99.94|Prostatic massage
C0194855|ICD9CM|HT|62|Operations on testes
C0194858|ICD9CM|PT|62.0|Incision of testis
C0194858|ICD9CM|AB|62.0|Incision of testes
C0194863|ICD9CM|AB|63.92|Epididymotomy
C0194863|ICD9CM|PT|63.92|Epididymotomy
C0194866|ICD9CM|PT|63.91|Aspiration of spermatocele
C0194866|ICD9CM|AB|63.91|Spermatocele aspiration
C0194873|ICD9CM|AB|62.3|Unilateral orchiectomy
C0194873|ICD9CM|PT|62.3|Unilateral orchiectomy
C0194876|ICD9CM|PT|62.42|Removal of remaining testis
C0194876|ICD9CM|AB|62.42|Remove solitary testis
C0194890|ICD9CM|AB|63.4|Epididymectomy
C0194890|ICD9CM|PT|63.4|Epididymectomy
C0194898|ICD9CM|PT|62.92|Injection of therapeutic substance into testis
C0194898|ICD9CM|AB|62.92|Injection into testes
C0194899|ICD9CM|PT|62.7|Insertion of testicular prosthesis
C0194899|ICD9CM|AB|62.7|Insert testicular prosth
C0194906|ICD9CM|HT|62.6|Repair of testes
C0194907|ICD9CM|AB|62.5|Orchiopexy
C0194907|ICD9CM|PT|62.5|Orchiopexy
C0194919|ICD9CM|HT|63.5|Repair of spermatic cord and epididymis
C0194920|ICD9CM|AB|63.83|Epididymovasostomy
C0194920|ICD9CM|PT|63.83|Epididymovasostomy
C0194924|ICD9CM|PT|63.51|Suture of laceration of spermatic cord and epididymis
C0194924|ICD9CM|AB|63.51|Suture cord & epid lacer
C0194939|ICD9CM|HT|60.7|Operations on seminal vesicles
C0194950|ICD9CM|PT|63.93|Incision of spermatic cord
C0194950|ICD9CM|AB|63.93|Spermatic cord incision
C0194957|ICD9CM|PT|60.72|Incision of seminal vesicle
C0194957|ICD9CM|AB|60.72|Seminal vesicle incision
C0194959|ICD9CM|PT|60.71|Percutaneous aspiration of seminal vesicle
C0194959|ICD9CM|AB|60.71|Percut semin ves aspirat
C0194971|ICD9CM|PT|63.84|Removal of ligature from vas deferens
C0194971|ICD9CM|AB|63.84|Removal vas ligature
C0194972|ICD9CM|PT|63.85|Removal of valve from vas deferens
C0194972|ICD9CM|AB|63.85|Remov vas deferens valve
C0194977|ICD9CM|PT|61.2|Excision of hydrocele (of tunica vaginalis)
C0194977|ICD9CM|AB|61.2|Excision of hydrocele
C0194992|ICD9CM|PT|60.73|Excision of seminal vesicle
C0194992|ICD9CM|AB|60.73|Seminal vesicle excision
C0194996|ICD9CM|PT|63.95|Insertion of valve in vas deferens
C0194996|ICD9CM|AB|63.95|Insert valve in vas def
C0195004|ICD9CM|PT|61.42|Repair of scrotal fistula
C0195004|ICD9CM|AB|61.42|Scrotal fistula repair
C0195021|ICD9CM|PT|63.72|Ligation of spermatic cord
C0195021|ICD9CM|AB|63.72|Spermatic cord ligation
C0195022|ICD9CM|PT|63.94|Lysis of adhesions of spermatic cord
C0195022|ICD9CM|AB|63.94|Sperm cord adhesiolysis
C0195047|ICD9CM|AB|71.4|Operations on clitoris
C0195047|ICD9CM|PT|71.4|Operations on clitoris
C0195048|ICD9CM|HT|71.2|Operations on Bartholin's gland
C0195067|ICD9CM|AB|71.61|Unilateral vulvectomy
C0195067|ICD9CM|PT|71.61|Unilateral vulvectomy
C0195098|ICD9CM|PT|71.01|Lysis of vulvar adhesions
C0195098|ICD9CM|AB|71.01|Vulvar adhesiolysis
C0195107|ICD9CM|PT|71.23|Marsupialization of Bartholin's gland (cyst)
C0195107|ICD9CM|AB|71.23|Bartholin gland marsup
C0195127|ICD9CM|AB|70.0|Culdocentesis
C0195127|ICD9CM|PT|70.0|Culdocentesis
C0195131|ICD9CM|AB|70.11|Hymenotomy
C0195131|ICD9CM|PT|70.11|Hymenotomy
C0195133|ICD9CM|AB|70.24|Vaginal biopsy
C0195133|ICD9CM|PT|70.24|Vaginal biopsy
C0195135|ICD9CM|PT|70.33|Excision or destruction of lesion of vagina
C0195135|ICD9CM|AB|70.33|Excision vaginal lesion
C0195147|ICD9CM|AB|70.31|Hymenectomy
C0195147|ICD9CM|PT|70.31|Hymenectomy
C0195150|ICD9CM|PT|70.23|Biopsy of cul-de-sac
C0195150|ICD9CM|AB|70.23|Cul-de-sac biopsy
C0195155|ICD9CM|PT|96.17|Insertion of vaginal diaphragm
C0195155|ICD9CM|AB|96.17|Vag diaphragm insertion
C0195157|ICD9CM|PT|97.73|Removal of vaginal diaphragm
C0195157|ICD9CM|AB|97.73|Remov vaginal diaphragm
C0195169|ICD9CM|PT|98.17|Removal of intraluminal foreign body from vagina without incision
C0195169|ICD9CM|AB|98.17|Remov intralum vag FB
C0195170|ICD9CM|PT|96.15|Insertion of vaginal mold
C0195170|ICD9CM|AB|96.15|Vaginal mold insertion
C0195191|ICD9CM|PT|70.8|Obliteration of vaginal vault
C0195191|ICD9CM|AB|70.8|Vaginal vault obliterat
C0195196|ICD9CM|AB|70.62|Vaginal reconstruction
C0195196|ICD9CM|PT|70.62|Vaginal reconstruction
C0195211|ICD9CM|PT|70.72|Repair of colovaginal fistula
C0195211|ICD9CM|AB|70.72|Repair colovagin fistula
C0195213|ICD9CM|PT|70.73|Repair of rectovaginal fistula
C0195213|ICD9CM|AB|70.73|Repair rectovag fistula
C0195230|ICD9CM|PT|70.52|Repair of rectocele
C0195230|ICD9CM|AB|70.52|Rectocele repair
C0195232|ICD9CM|HT|70.5|Repair of cystocele and rectocele
C0195232|ICD9CM|PT|70.50|Repair of cystocele and rectocele
C0195232|ICD9CM|AB|70.50|Cystocel/rectocel repair
C0195257|ICD9CM|HT|67|Operations on cervix
C0195270|ICD9CM|AB|69.95|Incision of cervix
C0195270|ICD9CM|PT|69.95|Incision of cervix
C0195277|ICD9CM|PT|98.16|Removal of intraluminal foreign body from uterus without incision
C0195277|ICD9CM|AB|98.16|Remov intralum uter FB
C0195289|ICD9CM|HT|68.3|Subtotal abdominal hysterectomy
C0195299|ICD9CM|HT|68.7|Radical vaginal hysterectomy
C0195324|ICD9CM|AB|67.2|Conization of cervix
C0195324|ICD9CM|PT|67.2|Conization of cervix
C0195331|ICD9CM|AB|67.4|Amputation of cervix
C0195331|ICD9CM|PT|67.4|Amputation of cervix
C0195341|ICD9CM|PT|69.96|Removal of cerclage material from cervix
C0195341|ICD9CM|AB|69.96|Remove cervical cerclage
C0195343|ICD9CM|AB|67.11|Endocervical biopsy
C0195343|ICD9CM|PT|67.11|Endocervical biopsy
C0195363|ICD9CM|PT|69.91|Insertion of therapeutic device into uterus
C0195363|ICD9CM|AB|69.91|Insert uterine device
C0195365|ICD9CM|PT|97.72|Removal of intrauterine pack
C0195365|ICD9CM|AB|97.72|Remov intrauterine pack
C0195379|ICD9CM|HT|69.4|Uterine repair
C0195404|ICD9CM|PT|69.42|Closure of fistula of uterus
C0195404|ICD9CM|AB|69.42|Closure uterine fistula
C0195410|ICD9CM|HT|67.5|Repair of internal cervical os
C0195412|ICD9CM|PT|67.62|Repair of fistula of cervix
C0195412|ICD9CM|AB|67.62|Cervical fistula repair
C0195436|ICD9CM|PT|68.21|Division of endometrial synechiae
C0195436|ICD9CM|AB|68.21|Endomet synechiae divis
C0195462|ICD9CM|HT|65.1|Diagnostic procedures on ovaries
C0195463|ICD9CM|HT|66|Operations on fallopian tubes
C0195465|ICD9CM|HT|65.0|Oophorotomy
C0195474|ICD9CM|AB|65.91|Aspiration of ovary
C0195474|ICD9CM|PT|65.91|Aspiration of ovary
C0195475|ICD9CM|AB|66.01|Salpingotomy
C0195475|ICD9CM|PT|66.01|Salpingotomy
C0195477|ICD9CM|PT|66.91|Aspiration of fallopian tube
C0195477|ICD9CM|AB|66.91|Fallopian tube aspirat
C0195495|ICD9CM|HT|65.6|Bilateral salpingo-oophorectomy
C0195504|ICD9CM|PT|66.11|Biopsy of fallopian tube
C0195504|ICD9CM|AB|66.11|Fallopian tube biopsy
C0195505|ICD9CM|PT|66.61|Excision or destruction of lesion of fallopian tube
C0195505|ICD9CM|AB|66.61|Destroy fallop tube les
C0195509|ICD9CM|HT|66.5|Total bilateral salpingectomy
C0195543|ICD9CM|PT|66.21|Bilateral endoscopic ligation and crushing of fallopian tubes
C0195543|ICD9CM|AB|66.21|Bilat endosc crush tube
C0195544|ICD9CM|PT|66.22|Bilateral endoscopic ligation and division of fallopian tubes
C0195544|ICD9CM|AB|66.22|Bilat endosc divis tube
C0195549|ICD9CM|HT|65.7|Repair of ovary
C0195551|ICD9CM|AB|66.72|Salpingo-oophorostomy
C0195551|ICD9CM|PT|66.72|Salpingo-oophorostomy
C0195553|ICD9CM|PT|65.95|Release of torsion of ovary
C0195553|ICD9CM|AB|65.95|Ovarian torsion release
C0195554|ICD9CM|PT|65.21|Marsupialization of ovarian cyst
C0195554|ICD9CM|AB|65.21|Ovarian cyst marsupializ
C0195561|ICD9CM|PT|66.97|Burying of fimbriae in uterine wall
C0195561|ICD9CM|AB|66.97|Bury fimbriae in uterus
C0195580|ICD9CM|HT|65.8|Lysis of adhesions of ovary and fallopian tube
C0195583|ICD9CM|AB|65.94|Ovarian denervation
C0195583|ICD9CM|PT|65.94|Ovarian denervation
C0195600|ICD9CM|PT|65.93|Manual rupture of ovarian cyst
C0195600|ICD9CM|AB|65.93|Manual rupt ovarian cyst
C0195601|ICD9CM|PT|66.96|Dilation of fallopian tube
C0195601|ICD9CM|AB|66.96|Fallopian tube dilation
C0195612|ICD9CM|PT|73.93|Incision of cervix to assist delivery
C0195612|ICD9CM|AB|73.93|Incis cx to assist deliv
C0195613|ICD9CM|PT|73.94|Pubiotomy to assist delivery
C0195613|ICD9CM|AB|73.94|Pubiotomy to assist del
C0195619|ICD9CM|PT|74.0|Classical cesarean section
C0195619|ICD9CM|AB|74.0|Classical c-section
C0195620|ICD9CM|PT|74.1|Low cervical cesarean section
C0195620|ICD9CM|AB|74.1|Low cervical c-section
C0195621|ICD9CM|PT|74.2|Extraperitoneal cesarean section
C0195621|ICD9CM|AB|74.2|Extraperitoneal c-sect
C0195641|ICD9CM|PT|69.01|Dilation and curettage for termination of pregnancy
C0195641|ICD9CM|AB|69.01|D & C for preg terminat
C0195643|ICD9CM|PT|74.91|Hysterotomy to terminate pregnancy
C0195643|ICD9CM|AB|74.91|Hysterotomy to termin pg
C0195679|ICD9CM|HT|75.5|Repair of current obstetric laceration of uterus
C0195679|ICD9CM|PT|75.52|Repair of current obstetric laceration of corpus uteri
C0195679|ICD9CM|PT|75.50|Repair of current obstetric laceration of uterus, not otherwise specified
C0195679|ICD9CM|AB|75.52|Repair ob lac corp uteri
C0195679|ICD9CM|AB|75.50|Repair ob lac uterus NOS
C0195704|ICD9CM|PT|73.51|Manual rotation of fetal head
C0195704|ICD9CM|AB|73.51|Manual rotat fetal head
C0195711|ICD9CM|PT|72.51|Partial breech extraction with forceps to aftercoming head
C0195711|ICD9CM|AB|72.51|Part brch extrac w forcp
C0195712|ICD9CM|PT|72.53|Total breech extraction with forceps to aftercoming head
C0195712|ICD9CM|AB|72.53|Tot brch extrac w forcep
C0195720|ICD9CM|AB|73.3|Failed forceps
C0195720|ICD9CM|PT|73.3|Failed forceps
C0195724|ICD9CM|AB|72.0|Low forceps operation
C0195724|ICD9CM|PT|72.0|Low forceps operation
C0195728|ICD9CM|HT|72.3|High forceps operation
C0195732|ICD9CM|PT|73.91|External version assisting delivery
C0195732|ICD9CM|AB|73.91|Ext version-assist deliv
C0195743|ICD9CM|PT|73.21|Internal and combined version without extraction
C0195743|ICD9CM|AB|73.21|Int/comb version no extr
C0195744|ICD9CM|PT|73.22|Internal and combined version with extraction
C0195744|ICD9CM|HT|73.2|Internal and combined version and extraction
C0195744|ICD9CM|AB|73.22|Int/comb version w extr
C0195755|ICD9CM|PT|75.4|Manual removal of retained placenta
C0195755|ICD9CM|AB|75.4|Manual removal-placenta
C0195756|ICD9CM|PT|75.7|Manual exploration of uterine cavity, postpartum
C0195756|ICD9CM|AB|75.7|Manual explor uterus p/p
C0195758|ICD9CM|PT|73.92|Replacement of prolapsed umbilical cord
C0195758|ICD9CM|AB|73.92|Replace prolapsed cord
C0195781|ICD9CM|PT|01.42|Operations on globus pallidus
C0195781|ICD9CM|AB|01.42|Globus pallidus ops
C0195791|ICD9CM|PT|01.23|Reopening of craniotomy site
C0195791|ICD9CM|AB|01.23|Reopen craniotomy site
C0195806|ICD9CM|PT|01.32|Lobotomy and tractotomy
C0195806|ICD9CM|AB|01.32|Lobotomy & tractotomy
C0195838|ICD9CM|HT|01.0|Cranial puncture
C0195842|ICD9CM|PT|01.31|Incision of cerebral meninges
C0195842|ICD9CM|AB|01.31|Incise cerebral meninges
C0195877|ICD9CM|AB|01.01|Cisternal puncture
C0195877|ICD9CM|PT|01.01|Cisternal puncture
C0195889|ICD9CM|PT|01.21|Incision and drainage of cranial sinus
C0195889|ICD9CM|AB|01.21|Cranial sinus i & d
C0195898|ICD9CM|PT|01.15|Biopsy of skull
C0195898|ICD9CM|AB|01.15|Skull biopsy
C0195899|ICD9CM|PT|01.6|Excision of lesion of skull
C0195899|ICD9CM|AB|01.6|Excise skull lesion
C0195916|ICD9CM|PT|01.13|Closed [percutaneous] [needle] biopsy of brain
C0195916|ICD9CM|AB|01.13|Closed brain biopsy
C0195961|ICD9CM|PT|01.53|Lobectomy of brain
C0195961|ICD9CM|AB|01.53|Brain lobectomy
C0195984|ICD9CM|PT|01.11|Closed [percutaneous] [needle] biopsy of cerebral meninges
C0195984|ICD9CM|AB|01.11|Clos cereb meninges bx
C0195997|ICD9CM|AB|02.14|Choroid plexectomy
C0195997|ICD9CM|PT|02.14|Choroid plexectomy
C0196024|ICD9CM|PT|02.05|Insertion of skull plate
C0196024|ICD9CM|AB|02.05|Skull plate insertion
C0196050|ICD9CM|PT|02.41|Irrigation and exploration of ventricular shunt
C0196050|ICD9CM|AB|02.41|Irrigate/expl vent shunt
C0196087|ICD9CM|PT|02.07|Removal of skull plate
C0196087|ICD9CM|AB|02.07|Skull plate removal
C0196103|ICD9CM|PT|02.43|Removal of ventricular shunt
C0196103|ICD9CM|AB|02.43|Remove ventricle shunt
C0196112|ICD9CM|HT|02.0|Cranioplasty
C0196118|ICD9CM|PT|02.02|Elevation of skull fracture fragments
C0196118|ICD9CM|AB|02.02|Elevate skull fx fragmnt
C0196162|ICD9CM|PT|02.11|Simple suture of dura mater of brain
C0196162|ICD9CM|AB|02.11|Simple suture of dura
C0196173|ICD9CM|PT|02.32|Ventricular shunt to circulatory system
C0196173|ICD9CM|AB|02.32|Ventri shunt-circula sys
C0196190|ICD9CM|PT|02.35|Ventricular shunt to urinary system
C0196190|ICD9CM|AB|02.35|Ventri shunt-uninary sys
C0196194|ICD9CM|HT|02.3|Extracranial ventricular shunt
C0196224|ICD9CM|AB|02.04|Bone graft to skull
C0196224|ICD9CM|PT|02.04|Bone graft to skull
C0196243|ICD9CM|AB|03.21|Percutaneous chordotomy
C0196243|ICD9CM|PT|03.21|Percutaneous chordotomy
C0196383|ICD9CM|PT|03.01|Removal of foreign body from spinal canal
C0196383|ICD9CM|AB|03.01|Removal FB spinal canal
C0196458|ICD9CM|PT|03.98|Removal of spinal thecal shunt
C0196458|ICD9CM|AB|03.98|Remove spine theca shunt
C0196469|ICD9CM|PT|03.51|Repair of spinal meningocele
C0196469|ICD9CM|AB|03.51|Spine meningocele repair
C0196477|ICD9CM|PT|03.52|Repair of spinal myelomeningocele
C0196477|ICD9CM|AB|03.52|Myelomeningocel repair
C0196487|ICD9CM|PT|03.71|Spinal subarachnoid-peritoneal shunt
C0196487|ICD9CM|AB|03.71|Subarach-periton shunt
C0196489|ICD9CM|PT|03.72|Spinal subarachnoid-ureteral shunt
C0196489|ICD9CM|AB|03.72|Subarach-ureteral shunt
C0196492|ICD9CM|PT|03.97|Revision of spinal thecal shunt
C0196492|ICD9CM|AB|03.97|Revise spine theca shunt
C0196504|ICD9CM|PT|03.8|Injection of destructive agent into spinal canal
C0196504|ICD9CM|AB|03.8|Destr inject-spine canal
C0196521|ICD9CM|PT|03.6|Lysis of adhesions of spinal cord and nerve roots
C0196521|ICD9CM|AB|03.6|Spinal cord adhesiolysis
C0196526|ICD9CM|PT|03.96|Percutaneous denervation of facet
C0196526|ICD9CM|AB|03.96|Percutan facet denervat
C0196576|ICD9CM|AB|04.43|Carpal tunnel release
C0196576|ICD9CM|PT|04.43|Release of carpal tunnel
C0196577|ICD9CM|AB|04.44|Tarsal tunnel release
C0196577|ICD9CM|PT|04.44|Release of tarsal tunnel
C0196589|ICD9CM|PT|04.41|Decompression of trigeminal nerve root
C0196589|ICD9CM|AB|04.41|Decompress trigem root
C0196608|ICD9CM|PT|29.92|Division of glossopharyngeal nerve
C0196608|ICD9CM|AB|29.92|Divis glossopharyng nerv
C0196609|ICD9CM|PT|31.91|Division of laryngeal nerve
C0196609|ICD9CM|AB|31.91|Laryngeal nerv division
C0196617|ICD9CM|PT|07.42|Division of nerves to adrenal glands
C0196617|ICD9CM|AB|07.42|Adrenal nerve division
C0196664|ICD9CM|AB|05.22|Cervical sympathectomy
C0196664|ICD9CM|PT|05.22|Cervical sympathectomy
C0196667|ICD9CM|AB|05.23|Lumbar sympathectomy
C0196667|ICD9CM|PT|05.23|Lumbar sympathectomy
C0196669|ICD9CM|AB|05.24|Presacral sympathectomy
C0196669|ICD9CM|PT|05.24|Presacral sympathectomy
C0196674|ICD9CM|PT|05.25|Periarterial sympathectomy
C0196674|ICD9CM|AB|05.25|Periart sympathectomy
C0196686|ICD9CM|AB|04.05|Gasserian ganglionectomy
C0196686|ICD9CM|PT|04.05|Gasserian ganglionectomy
C0196687|ICD9CM|PT|05.21|Sphenopalatine ganglionectomy
C0196687|ICD9CM|AB|05.21|Sphenopalatin ganglionec
C0196696|ICD9CM|PT|04.80|Peripheral nerve injection, not otherwise specified
C0196696|ICD9CM|AB|04.80|Periph nerve inject NOS
C0196806|ICD9CM|PT|04.72|Accessory-facial anastomosis
C0196806|ICD9CM|AB|04.72|Accessory-facial anastom
C0196807|ICD9CM|PT|04.73|Accessory-hypoglossal anastomosis
C0196807|ICD9CM|AB|04.73|Access-hypogloss anastom
C0196809|ICD9CM|PT|69.3|Paracervical uterine denervation
C0196809|ICD9CM|AB|69.3|Paracerv uterine denerv
C0196940|ICD9CM|AB|04.91|Neurectasis
C0196940|ICD9CM|PT|04.91|Neurectasis
C0196947|ICD9CM|HT|16|Operations on orbit and eyeball
C0196952|ICD9CM|HT|16.6|Secondary procedures after removal of eyeball
C0196955|ICD9CM|PT|16.01|Orbitotomy with bone flap
C0196955|ICD9CM|AB|16.01|Orbitotomy w bone flap
C0196969|ICD9CM|PT|16.23|Biopsy of eyeball and orbit
C0196969|ICD9CM|AB|16.23|Eyeball & orbit biopsy
C0196972|ICD9CM|PT|16.22|Diagnostic aspiration of orbit
C0196972|ICD9CM|AB|16.22|Diagnostic asp of orbit
C0196973|ICD9CM|PT|16.92|Excision of lesion of orbit
C0196973|ICD9CM|AB|16.92|Excision orbital lesion
C0196984|ICD9CM|PT|16.52|Exenteration of orbit with therapeutic removal of orbital bone
C0196984|ICD9CM|AB|16.52|Orbit exent w bone remov
C0196985|ICD9CM|PT|16.51|Exenteration of orbit with removal of adjacent structures
C0196985|ICD9CM|AB|16.51|Radical orbitomaxillect
C0196988|ICD9CM|PT|16.41|Enucleation of eyeball with synchronous implant into Tenon's capsule with attachment of muscles
C0196988|ICD9CM|AB|16.41|Eye enuc/implan/musc att
C0196990|ICD9CM|PT|98.21|Removal of superficial foreign body from eye without incision
C0196990|ICD9CM|AB|98.21|Removal superfic FB eye
C0196991|ICD9CM|PT|16.1|Removal of penetrating foreign body from eye, not otherwise specified
C0196991|ICD9CM|AB|16.1|Remove penetrat FB eye
C0196999|ICD9CM|PT|16.91|Retrobulbar injection of therapeutic agent
C0196999|ICD9CM|AB|16.91|Retrobulbar injection
C0197003|ICD9CM|PT|16.61|Secondary insertion of ocular implant
C0197003|ICD9CM|AB|16.61|2ndry ocular imp insert
C0197017|ICD9CM|PT|16.71|Removal of ocular implant
C0197017|ICD9CM|AB|16.71|Remove ocular implant
C0197019|ICD9CM|PT|16.72|Removal of orbital implant
C0197019|ICD9CM|AB|16.72|Remove orbital implant
C0197022|ICD9CM|PT|16.62|Revision and reinsertion of ocular implant
C0197022|ICD9CM|AB|16.62|Revis/reinsert ocul imp
C0197030|ICD9CM|PT|16.81|Repair of wound of orbit
C0197030|ICD9CM|AB|16.81|Repair of orbital wound
C0197034|ICD9CM|PT|16.63|Revision of enucleation socket with graft
C0197034|ICD9CM|AB|16.63|Revis enuc socket w grft
C0197050|ICD9CM|HT|08|Operations on eyelids
C0197051|ICD9CM|HT|08.1|Diagnostic procedures on eyelid
C0197056|ICD9CM|HT|09|Operations on lacrimal system
C0197057|ICD9CM|HT|09.1|Diagnostic procedures on lacrimal system
C0197059|ICD9CM|HT|10|Operations on conjunctiva
C0197060|ICD9CM|HT|10.2|Diagnostic procedures on conjunctiva
C0197063|ICD9CM|HT|08.0|Incision of eyelid
C0197064|ICD9CM|AB|08.01|Incision of lid margin
C0197064|ICD9CM|PT|08.01|Incision of lid margin
C0197075|ICD9CM|AB|08.51|Canthotomy
C0197075|ICD9CM|PT|08.51|Canthotomy
C0197083|ICD9CM|PT|09.0|Incision of lacrimal gland
C0197083|ICD9CM|AB|09.0|Lacrimal gland incision
C0197086|ICD9CM|PT|09.52|Incision of lacrimal canaliculi
C0197086|ICD9CM|AB|09.52|Lac canaliculi incision
C0197088|ICD9CM|PT|09.51|Incision of lacrimal punctum
C0197088|ICD9CM|AB|09.51|Lac punctum incision
C0197105|ICD9CM|PT|08.23|Excision of major lesion of eyelid, partial-thickness
C0197105|ICD9CM|AB|08.23|Exc maj les lid prt-thic
C0197124|ICD9CM|PT|08.86|Lower eyelid rhytidectomy
C0197124|ICD9CM|AB|08.86|Lower lid rhytidectomy
C0197125|ICD9CM|PT|08.87|Upper eyelid rhytidectomy
C0197125|ICD9CM|AB|08.87|Upper lid rhytidectomy
C0197128|ICD9CM|AB|10.21|Conjunctival biopsy
C0197128|ICD9CM|PT|10.21|Biopsy of conjunctiva
C0197133|ICD9CM|HT|11.3|Excision of pterygium
C0197139|ICD9CM|PT|09.11|Biopsy of lacrimal gland
C0197139|ICD9CM|AB|09.11|Lacrimal gland biopsy
C0197140|ICD9CM|PT|09.12|Biopsy of lacrimal sac
C0197140|ICD9CM|AB|09.12|Lacrimal sac biopsy
C0197145|ICD9CM|PT|09.20|Excision of lacrimal gland, not otherwise specified
C0197145|ICD9CM|AB|09.20|Exc lacrimal gland NOS
C0197147|ICD9CM|AB|09.23|Total dacryoadenectomy
C0197147|ICD9CM|PT|09.23|Total dacryoadenectomy
C0197180|ICD9CM|PT|10.91|Subconjunctival injection
C0197180|ICD9CM|AB|10.91|Subconjunctival inject
C0197182|ICD9CM|PT|09.41|Probing of lacrimal punctum
C0197182|ICD9CM|AB|09.41|Lacrimal punctum probe
C0197185|ICD9CM|PT|09.42|Probing of lacrimal canaliculi
C0197185|ICD9CM|AB|09.42|Lac canaliculi probe
C0197194|ICD9CM|PT|09.44|Intubation of nasolacrimal duct
C0197194|ICD9CM|AB|09.44|Nasolac duct intubat
C0197223|ICD9CM|PT|08.82|Repair of laceration involving lid margin, partial-thickness
C0197223|ICD9CM|AB|08.82|Lid marg lac rx-part th
C0197225|ICD9CM|PT|08.84|Repair of laceration involving lid margin, full-thickness
C0197225|ICD9CM|AB|08.84|Lid marg lac rx-ful thic
C0197226|ICD9CM|PT|08.38|Correction of lid retraction
C0197226|ICD9CM|AB|08.38|Correct lid retraction
C0197254|ICD9CM|HT|10.4|Conjunctivoplasty
C0197255|ICD9CM|PT|10.6|Repair of laceration of conjunctiva
C0197255|ICD9CM|AB|10.6|Repair conjunct lacerat
C0197270|ICD9CM|PT|11.31|Transposition of pterygium
C0197270|ICD9CM|AB|11.31|Pterygium transposition
C0197283|ICD9CM|PT|08.31|Repair of blepharoptosis by frontalis muscle technique with suture
C0197283|ICD9CM|AB|08.31|Ptosis rep-front mus sut
C0197284|ICD9CM|PT|08.32|Repair of blepharoptosis by frontalis muscle technique with fascial sling
C0197284|ICD9CM|AB|08.32|Ptosis rep-fron mus slng
C0197286|ICD9CM|PT|08.34|Repair of blepharoptosis by other levator muscle techniques
C0197286|ICD9CM|AB|08.34|Ptosis rep-levat mus NEC
C0197292|ICD9CM|PT|08.35|Repair of blepharoptosis by tarsal technique
C0197292|ICD9CM|AB|08.35|Ptos rep-tarsal techniq
C0197300|ICD9CM|PT|08.37|Reduction of overcorrection of ptosis
C0197300|ICD9CM|AB|08.37|Reduc overcorrect ptosis
C0197313|ICD9CM|PT|08.70|Reconstruction of eyelid, not otherwise specified
C0197313|ICD9CM|AB|08.70|Lid reconstruction NOS
C0197316|ICD9CM|PT|08.71|Reconstruction of eyelid involving lid margin, partial-thickness
C0197316|ICD9CM|AB|08.71|Lid marg recon-part thic
C0197318|ICD9CM|PT|08.73|Reconstruction of eyelid involving lid margin, full-thickness
C0197318|ICD9CM|AB|08.73|Lid marg recons ful thic
C0197323|ICD9CM|PT|08.63|Reconstruction of eyelid with hair follicle graft
C0197323|ICD9CM|AB|08.63|Lid reconst w hair graft
C0197324|ICD9CM|PT|08.64|Reconstruction of eyelid with tarsoconjunctival flap
C0197324|ICD9CM|AB|08.64|Lid recon-tarsoconj flap
C0197334|ICD9CM|PT|10.41|Repair of symblepharon with free graft
C0197334|ICD9CM|AB|10.41|Symbleph rep w free grft
C0197346|ICD9CM|PT|09.91|Obliteration of lacrimal punctum
C0197346|ICD9CM|AB|09.91|Lac punctum obliteration
C0197353|ICD9CM|PT|08.25|Destruction of lesion of eyelid
C0197353|ICD9CM|AB|08.25|Destruction lid lesion
C0197363|ICD9CM|PT|08.92|Cryosurgical epilation of eyelid
C0197363|ICD9CM|AB|08.92|Cryosurg lid epilation
C0197372|ICD9CM|PT|10.32|Destruction of lesion of conjunctiva
C0197372|ICD9CM|AB|10.32|Destruct conjunc les NEC
C0197393|ICD9CM|HT|09.4|Manipulation of lacrimal passage
C0197397|ICD9CM|PT|09.43|Probing of nasolacrimal duct
C0197397|ICD9CM|AB|09.43|Nasolacrimal duct probe
C0197402|ICD9CM|HT|11|Operations on cornea
C0197403|ICD9CM|HT|11.2|Diagnostic procedures on cornea
C0197405|ICD9CM|PT|11.1|Incision of cornea
C0197405|ICD9CM|AB|11.1|Corneal incision
C0197411|ICD9CM|PT|11.41|Mechanical removal of corneal epithelium
C0197411|ICD9CM|AB|11.41|Mech remov cornea epith
C0197417|ICD9CM|AB|11.22|Corneal biopsy
C0197417|ICD9CM|PT|11.22|Biopsy of cornea
C0197424|ICD9CM|PT|11.92|Removal of artificial implant from cornea
C0197424|ICD9CM|AB|11.92|Remove corneal implant
C0197431|ICD9CM|PT|11.91|Tattooing of cornea
C0197431|ICD9CM|AB|11.91|Corneal tattooing
C0197440|ICD9CM|PT|11.61|Lamellar keratoplasty with autograft
C0197440|ICD9CM|AB|11.61|Lam keratplast w autgrft
C0197444|ICD9CM|PT|11.63|Penetrating keratoplasty with autograft
C0197444|ICD9CM|AB|11.63|Perf keratopl w autogrft
C0197448|ICD9CM|AB|11.72|Keratophakia
C0197448|ICD9CM|PT|11.72|Keratophakia
C0197453|ICD9CM|PT|11.52|Repair of postoperative wound dehiscence of cornea
C0197453|ICD9CM|AB|11.52|Rep cornea postop dehisc
C0197455|ICD9CM|PT|11.51|Suture of corneal laceration
C0197455|ICD9CM|AB|11.51|Suture cornea laceration
C0197459|ICD9CM|AB|11.74|Thermokeratoplasty
C0197459|ICD9CM|PT|11.74|Thermokeratoplasty
C0197472|ICD9CM|PT|11.43|Cryotherapy of corneal lesion
C0197472|ICD9CM|AB|11.43|Cryotherap cornea lesion
C0197494|ICD9CM|HT|12.8|Operations on sclera
C0197499|ICD9CM|PT|12.11|Iridotomy with transfixion
C0197499|ICD9CM|AB|12.11|Iridotomy w transfixion
C0197511|ICD9CM|PT|12.91|Therapeutic evacuation of anterior chamber
C0197511|ICD9CM|AB|12.91|Therapeut evac ant chamb
C0197512|ICD9CM|PT|12.21|Diagnostic aspiration of anterior chamber of eye
C0197512|ICD9CM|AB|12.21|Dx aspirat-ant chamber
C0197526|ICD9CM|AB|12.55|Cyclodialysis
C0197526|ICD9CM|PT|12.55|Cyclodialysis
C0197527|ICD9CM|PT|12.53|Goniotomy with goniopuncture
C0197527|ICD9CM|AB|12.53|Goniotomy w goniopunctur
C0197534|ICD9CM|AB|12.54|Trabeculotomy ab externo
C0197534|ICD9CM|PT|12.54|Trabeculotomy ab externo
C0197538|ICD9CM|HT|12.6|Scleral fistulization
C0197540|ICD9CM|HT|12.5|Facilitation of intraocular circulation
C0197542|ICD9CM|PT|12.40|Removal of lesion of anterior segment of eye, not otherwise specified
C0197542|ICD9CM|AB|12.40|Remov ant segmnt les NOS
C0197545|ICD9CM|PT|12.22|Biopsy of iris
C0197545|ICD9CM|AB|12.22|Iris biopsy
C0197546|ICD9CM|PT|12.42|Excision of lesion of iris
C0197546|ICD9CM|AB|12.42|Excision of iris lesion
C0197547|ICD9CM|PT|12.13|Excision of prolapsed iris
C0197547|ICD9CM|AB|12.13|Prolapsed iris excision
C0197549|ICD9CM|PT|12.44|Excision of lesion of ciliary body
C0197549|ICD9CM|AB|12.44|Excise ciliary body les
C0197562|ICD9CM|PT|12.61|Trephination of sclera with iridectomy
C0197562|ICD9CM|AB|12.61|Trephin sclera w iridect
C0197582|ICD9CM|HT|12.0|Removal of intraocular foreign body from anterior segment of eye
C0197582|ICD9CM|PT|12.00|Removal of intraocular foreign body from anterior segment of eye, not otherwise specified
C0197582|ICD9CM|AB|12.00|Remov ant segmnt FB NOS
C0197593|ICD9CM|PT|12.01|Removal of intraocular foreign body from anterior segment of eye with use of magnet
C0197593|ICD9CM|AB|12.01|Magnet remov ant seg FB
C0197613|ICD9CM|AB|12.35|Coreoplasty
C0197613|ICD9CM|PT|12.35|Coreoplasty
C0197621|ICD9CM|PT|12.63|Iridencleisis and iridotasis
C0197621|ICD9CM|AB|12.63|Iridencleisis/iridotasis
C0197622|ICD9CM|PT|12.82|Repair of scleral fistula
C0197622|ICD9CM|AB|12.82|Scleral fistula repair
C0197624|ICD9CM|PT|12.85|Repair of scleral staphyloma with graft
C0197624|ICD9CM|AB|12.85|Repair staphylom w graft
C0197625|ICD9CM|PT|12.81|Suture of laceration of sclera
C0197625|ICD9CM|AB|12.81|Suture scleral lacer
C0197630|ICD9CM|PT|12.66|Postoperative revision of scleral fistulization procedure
C0197630|ICD9CM|AB|12.66|Postop revis scl fistul
C0197641|ICD9CM|PT|12.74|Diminution of ciliary body, not otherwise specified
C0197641|ICD9CM|AB|12.74|Cil body diminution NOS
C0197646|ICD9CM|PT|12.41|Destruction of lesion of iris, nonexcisional
C0197646|ICD9CM|AB|12.41|Nonexc destruc iris les
C0197648|ICD9CM|PT|12.31|Lysis of goniosynechiae
C0197648|ICD9CM|AB|12.31|Goniosynechiae lysis
C0197652|ICD9CM|PT|12.33|Lysis of posterior synechiae
C0197652|ICD9CM|AB|12.33|Post synechiae lysis
C0197653|ICD9CM|PT|12.34|Lysis of corneovitreal adhesions
C0197653|ICD9CM|AB|12.34|Corneovitreal adhesiolys
C0197663|ICD9CM|PT|12.43|Destruction of lesion of ciliary body, nonexcisional
C0197663|ICD9CM|AB|12.43|Nonexc destr cil bod les
C0197672|ICD9CM|HT|13|Operations on lens
C0197717|ICD9CM|HT|13.1|Intracapsular extraction of lens
C0197723|ICD9CM|PT|13.11|Intracapsular extraction of lens by temporal inferior route
C0197723|ICD9CM|AB|13.11|Temp-inf intrcap lens ex
C0197729|ICD9CM|PT|13.2|Extracapsular extraction of lens by linear extraction technique
C0197729|ICD9CM|AB|13.2|Linear extracap lens ext
C0197736|ICD9CM|PT|13.51|Extracapsular extraction of lens by temporal inferior route
C0197736|ICD9CM|AB|13.51|Temp-inf xtracap lens ex
C0197741|ICD9CM|HT|13.0|Removal of foreign body from lens
C0197741|ICD9CM|PT|13.00|Removal of foreign body from lens, not otherwise specified
C0197741|ICD9CM|AB|13.00|Remove FB lens NOS
C0197742|ICD9CM|PT|13.02|Removal of foreign body from lens without use of magnet
C0197742|ICD9CM|AB|13.02|Nonmagnet remove FB lens
C0197743|ICD9CM|PT|13.01|Removal of foreign body from lens with use of magnet
C0197743|ICD9CM|AB|13.01|Magnet remove FB lens
C0197750|ICD9CM|PT|13.72|Secondary insertion of intraocular lens prosthesis
C0197750|ICD9CM|AB|13.72|Secondary insert lens
C0197762|ICD9CM|PT|13.66|Mechanical fragmentation of secondary membrane [after cataract]
C0197762|ICD9CM|AB|13.66|After catar fragmntation
C0197784|ICD9CM|PT|14.11|Diagnostic aspiration of vitreous
C0197784|ICD9CM|AB|14.11|Diagnost vitreous aspir
C0197786|ICD9CM|PT|14.71|Removal of vitreous, anterior approach
C0197786|ICD9CM|AB|14.71|Anterior remov vitreous
C0197792|ICD9CM|PT|14.73|Mechanical vitrectomy by anterior approach
C0197792|ICD9CM|AB|14.73|Anterior mechan vitrect
C0197802|ICD9CM|HT|14.0|Removal of foreign body from posterior segment of eye
C0197802|ICD9CM|PT|14.00|Removal of foreign body from posterior segment of eye, not otherwise specified
C0197802|ICD9CM|AB|14.00|Remov post segmnt FB NOS
C0197806|ICD9CM|PT|14.01|Removal of foreign body from posterior segment of eye with use of magnet
C0197806|ICD9CM|AB|14.01|Magnet remov post seg FB
C0197812|ICD9CM|PT|14.02|Removal of foreign body from posterior segment of eye without use of magnet
C0197812|ICD9CM|AB|14.02|Nonmag remov post seg FB
C0197827|ICD9CM|PT|14.6|Removal of surgically implanted material from posterior segment of eye
C0197827|ICD9CM|AB|14.6|Remov pros mat post seg
C0197875|ICD9CM|PT|14.52|Repair of retinal detachment with cryotherapy
C0197875|ICD9CM|AB|14.52|Detach retina-cryotherap
C0197888|ICD9CM|PT|14.33|Repair of retinal tear by xenon arc photocoagulation
C0197888|ICD9CM|AB|14.33|Retinal tear xenon coag
C0197902|ICD9CM|PT|14.21|Destruction of chorioretinal lesion by diathermy
C0197902|ICD9CM|AB|14.21|Chorioret les diathermy
C0197912|ICD9CM|PT|14.22|Destruction of chorioretinal lesion by cryotherapy
C0197912|ICD9CM|AB|14.22|Chorioretin les cryother
C0197920|ICD9CM|PT|14.23|Destruction of chorioretinal lesion by xenon arc photocoagulation
C0197920|ICD9CM|AB|14.23|Chorioret les xenon coag
C0197923|ICD9CM|PT|14.24|Destruction of chorioretinal lesion by laser photocoagulation
C0197923|ICD9CM|AB|14.24|Chorioret les laser coag
C0197926|ICD9CM|PT|14.26|Destruction of chorioretinal lesion by radiation therapy
C0197926|ICD9CM|AB|14.26|Chorioret les radiother
C0197930|ICD9CM|PT|14.27|Destruction of chorioretinal lesion by implantation of radiation source
C0197930|ICD9CM|AB|14.27|Chorioret les rad implan
C0197937|ICD9CM|HT|15|Operations on extraocular muscles
C0197943|ICD9CM|PT|15.3|Operations on two or more extraocular muscles involving temporary detachment from globe, one or both eyes
C0197943|ICD9CM|AB|15.3|Temp detach >1 xtroc mus
C0197958|ICD9CM|PT|15.13|Resection of one extraocular muscle
C0197958|ICD9CM|AB|15.13|1 extraoc muscl resect
C0197972|ICD9CM|PT|15.11|Recession of one extraocular muscle
C0197972|ICD9CM|AB|15.11|One extraoc mus recess
C0197999|ICD9CM|PT|15.6|Revision of extraocular muscle surgery
C0197999|ICD9CM|AB|15.6|Revis extraoc musc surg
C0198005|ICD9CM|PT|15.5|Transposition of extraocular muscles
C0198005|ICD9CM|AB|15.5|Extraocul mus transposit
C0198010|ICD9CM|HT|18-20.99|OPERATIONS ON THE EAR
C0198011|ICD9CM|HT|18|Operations on external ear
C0198012|ICD9CM|HT|18.1|Diagnostic procedures on external ear
C0198014|ICD9CM|HT|18.0|Incision of external ear
C0198025|ICD9CM|PT|18.02|Incision of external auditory canal
C0198025|ICD9CM|AB|18.02|Ext auditory canal incis
C0198030|ICD9CM|PT|18.12|Biopsy of external ear
C0198030|ICD9CM|AB|18.12|External ear biopsy
C0198044|ICD9CM|PT|18.31|Radical excision of lesion of external ear
C0198044|ICD9CM|AB|18.31|Rad excis ext ear les
C0198052|ICD9CM|PT|98.11|Removal of intraluminal foreign body from ear without incision
C0198052|ICD9CM|AB|98.11|Remov intralum ear FB
C0198057|ICD9CM|PT|96.11|Packing of external auditory canal
C0198057|ICD9CM|AB|96.11|Pack ext auditory canal
C0198066|ICD9CM|PT|18.5|Surgical correction of prominent ear
C0198066|ICD9CM|AB|18.5|Correction prominent ear
C0198075|ICD9CM|PT|18.4|Suture of laceration of external ear
C0198075|ICD9CM|AB|18.4|Suture ext ear lac
C0198097|ICD9CM|PT|20.23|Incision of middle ear
C0198097|ICD9CM|AB|20.23|Middle ear incision
C0198122|ICD9CM|PT|20.21|Incision of mastoid
C0198122|ICD9CM|AB|20.21|Mastoid incision
C0198132|ICD9CM|PT|20.51|Excision of lesion of middle ear
C0198132|ICD9CM|AB|20.51|Excise middle ear lesion
C0198142|ICD9CM|AB|20.91|Tympanosympathectomy
C0198142|ICD9CM|PT|20.91|Tympanosympathectomy
C0198143|ICD9CM|PT|19.11|Stapedectomy with incus replacement
C0198143|ICD9CM|AB|19.11|Stapedect w replac incus
C0198154|ICD9CM|HT|20.4|Mastoidectomy
C0198159|ICD9CM|AB|20.42|Radical mastoidectomy
C0198159|ICD9CM|PT|20.42|Radical mastoidectomy
C0198162|ICD9CM|PT|20.92|Revision of mastoidectomy
C0198162|ICD9CM|AB|20.92|Mastoidectomy revision
C0198183|ICD9CM|PT|20.94|Injection of tympanum
C0198183|ICD9CM|AB|20.94|Tympanic injection
C0198206|ICD9CM|PT|19.53|Type III tympanoplasty
C0198206|ICD9CM|AB|19.53|Type 3 tympanoplasty
C0198291|ICD9CM|PT|20.72|Injection into inner ear
C0198291|ICD9CM|AB|20.72|Inner ear injection
C0198293|ICD9CM|PT|20.95|Implantation of electromagnetic hearing device
C0198293|ICD9CM|AB|20.95|Elecmag hear dev implant
C0198308|ICD9CM|PT|20.93|Repair of oval and round windows
C0198308|ICD9CM|AB|20.93|Repair oval/round window
C0198318|ICD9CM|PT|20.62|Revision of fenestration of inner ear
C0198318|ICD9CM|AB|20.62|Revis inner ear fenestra
C0198375|ICD9CM|HT|34.7|Repair of chest wall
C0198376|ICD9CM|PT|34.71|Suture of laceration of chest wall
C0198376|ICD9CM|AB|34.71|Suture chest wall lacer
C0198378|ICD9CM|PT|34.72|Closure of thoracostomy
C0198378|ICD9CM|AB|34.72|Thoracostomy closure
C0198402|ICD9CM|AB|34.1|Incision of mediastinum
C0198402|ICD9CM|PT|34.1|Incision of mediastinum
C0198419|ICD9CM|PT|97.42|Removal of mediastinal drain
C0198419|ICD9CM|AB|97.42|Remov mediastinal drain
C0198438|ICD9CM|HT|34.8|Operations on diaphragm
C0198442|ICD9CM|AB|34.27|Biopsy of diaphragm
C0198442|ICD9CM|PT|34.27|Biopsy of diaphragm
C0198448|ICD9CM|PT|34.85|Implantation of diaphragmatic pacemaker
C0198448|ICD9CM|AB|34.85|Implant diaphra pacemake
C0198451|ICD9CM|PT|34.82|Suture of laceration of diaphragm
C0198451|ICD9CM|AB|34.82|Suture diaphragm lacerat
C0198452|ICD9CM|PT|34.83|Closure of fistula of diaphragm
C0198452|ICD9CM|AB|34.83|Close diaphragm fistula
C0198453|ICD9CM|PT|53.81|Plication of the diaphragm
C0198453|ICD9CM|AB|53.81|Diaphragmatic plication
C0198463|ICD9CM|HT|53.7|Repair of diaphragmatic hernia, abdominal approach
C0198464|ICD9CM|HT|53.8|Repair of diaphragmatic hernia, thoracic approach
C0198464|ICD9CM|PT|53.80|Repair of diaphragmatic hernia with thoracic approach, not otherwise specified
C0198464|ICD9CM|AB|53.80|Thor rep-diaph hern NOS
C0198471|ICD9CM|PT|53.82|Repair of parasternal hernia
C0198471|ICD9CM|AB|53.82|Parastern hernia repair
C0198489|ICD9CM|PT|54.0|Incision of abdominal wall
C0198489|ICD9CM|AB|54.0|Abdominal wall incision
C0198497|ICD9CM|PT|54.91|Percutaneous abdominal drainage
C0198497|ICD9CM|AB|54.91|Percu abdominal drainage
C0198525|ICD9CM|PT|54.97|Injection of locally-acting therapeutic substance into peritoneal cavity
C0198525|ICD9CM|AB|54.97|Inj therap subst periton
C0198534|ICD9CM|PT|97.81|Removal of retroperitoneal drainage device
C0198534|ICD9CM|AB|97.81|Remov retroperiton drain
C0198544|ICD9CM|PT|54.62|Delayed closure of granulating abdominal wound
C0198544|ICD9CM|AB|54.62|Delayed clos abd wound
C0198546|ICD9CM|PT|54.61|Reclosure of postoperative disruption of abdominal wall
C0198546|ICD9CM|AB|54.61|Reclose post op disrupt
C0198566|ICD9CM|AB|54.71|Repair of gastroschisis
C0198566|ICD9CM|PT|54.71|Repair of gastroschisis
C0198593|ICD9CM|PT|54.95|Incision of peritoneum
C0198593|ICD9CM|AB|54.95|Peritoneal incision
C0198609|ICD9CM|PT|54.23|Biopsy of peritoneum
C0198609|ICD9CM|AB|54.23|Peritoneal biopsy
C0198632|ICD9CM|PT|54.96|Injection of air into peritoneal cavity
C0198632|ICD9CM|AB|54.96|Injec air-periton cavity
C0198639|ICD9CM|PT|54.64|Suture of peritoneum
C0198639|ICD9CM|AB|54.64|Peritoneal suture
C0198644|ICD9CM|PT|54.93|Creation of cutaneoperitoneal fistula
C0198644|ICD9CM|AB|54.93|Create cutanperiton fist
C0198664|ICD9CM|HT|54.5|Lysis of peritoneal adhesions
C0198737|ICD9CM|PT|53.10|Bilateral repair of inguinal hernia, not otherwise specified
C0198737|ICD9CM|AB|53.10|Bilat ing hernia rep NOS
C0198742|ICD9CM|PT|53.05|Repair of inguinal hernia with graft or prosthesis, not otherwise specified
C0198742|ICD9CM|AB|53.05|Ing hernia rep-graft NOS
C0198745|ICD9CM|PT|53.17|Bilateral inguinal hernia repair with graft or prosthesis, not otherwise specified
C0198745|ICD9CM|AB|53.17|Bil ing hrn rep-grft NOS
C0198760|ICD9CM|HT|53.2|Unilateral repair of femoral hernia
C0198761|ICD9CM|HT|53.3|Bilateral repair of femoral hernia
C0198762|ICD9CM|PT|53.21|Unilateral repair of femoral hernia with graft or prosthesis
C0198762|ICD9CM|AB|53.21|Unil femor hrn rep-grft
C0198763|ICD9CM|PT|53.31|Bilateral repair of femoral hernia with graft or prosthesis
C0198763|ICD9CM|AB|53.31|Bil fem hern repair-grft
C0198793|ICD9CM|PT|96.27|Manual reduction of hernia
C0198793|ICD9CM|AB|96.27|Manual reduction hernia
C0198807|ICD9CM|PT|04.81|Injection of anesthetic into peripheral nerve for analgesia
C0198807|ICD9CM|AB|04.81|Anesth injec periph nerv
C0199177|ICD9CM|AB|89.06|Limited consultation
C0199177|ICD9CM|PT|89.06|Consultation, described as limited
C0199178|ICD9CM|PT|89.07|Consultation, described as comprehensive
C0199178|ICD9CM|AB|89.07|Comprehensive consultat
C0199182|ICD9CM|PT|89.05|Diagnostic interview and evaluation, not otherwise specified
C0199182|ICD9CM|AB|89.05|Interview & evaluat NOS
C0199403|ICD9CM|PT|94.45|Drug addiction counseling
C0199403|ICD9CM|AB|94.45|Drug addict counselling
C0199404|ICD9CM|PT|94.46|Alcoholism counseling
C0199404|ICD9CM|AB|94.46|Alcoholism counselling
C0199420|ICD9CM|AB|89.12|Nasal function study
C0199420|ICD9CM|PT|89.12|Nasal function study
C0199430|ICD9CM|PT|89.35|Transillumination of nasal sinuses
C0199430|ICD9CM|AB|89.35|Nasal sinus transillumin
C0199447|ICD9CM|AB|93.94|Nebulizer therapy
C0199447|ICD9CM|PT|93.94|Respiratory medication administered by nebulizer
C0199472|ICD9CM|AB|93.97|Decompression chamber
C0199472|ICD9CM|PT|93.97|Decompression chamber
C0199550|ICD9CM|AB|99.61|Atrial cardioversion
C0199550|ICD9CM|PT|99.61|Atrial cardioversion
C0199551|ICD9CM|PT|37.26|Catheter based invasive electrophysiologic testing
C0199551|ICD9CM|AB|37.26|Cath base invasv ep test
C0199553|ICD9CM|AB|37.27|Cardiac mapping
C0199553|ICD9CM|PT|37.27|Cardiac mapping
C0199556|ICD9CM|AB|89.51|Rhythm electrocardiogram
C0199556|ICD9CM|PT|89.51|Rhythm electrocardiogram
C0199581|ICD9CM|PT|89.56|Carotid pulse tracing with ECG lead
C0199581|ICD9CM|AB|89.56|Carotid pulse tracing
C0199597|ICD9CM|PT|89.55|Phonocardiogram with ECG lead
C0199597|ICD9CM|AB|89.55|Phonocardiogram
C0199605|ICD9CM|PT|89.53|Vectorcardiogram (with ECG)
C0199605|ICD9CM|AB|89.53|Vectorcardiogram
C0199612|ICD9CM|PT|89.57|Apexcardiogram (with ECG lead)
C0199612|ICD9CM|AB|89.57|Apexcardiogram
C0199624|ICD9CM|PT|89.67|Monitoring of cardiac output by oxygen consumption technique
C0199624|ICD9CM|AB|89.67|Oxygen consumption monit
C0199627|ICD9CM|PT|89.68|Monitoring of cardiac output by other technique
C0199627|ICD9CM|AB|89.68|Oth cardiac mon output
C0199629|ICD9CM|PT|89.63|Pulmonary artery pressure monitoring
C0199629|ICD9CM|AB|89.63|Pulmon art press monitor
C0199631|ICD9CM|PT|89.69|Monitoring of coronary blood flow
C0199631|ICD9CM|AB|89.69|Coronary bld flow monit
C0199655|ICD9CM|PT|39.64|Intraoperative cardiac pacemaker
C0199655|ICD9CM|AB|39.64|Intraop cardiac pacemak
C0199699|ICD9CM|PT|89.45|Artificial pacemaker rate check
C0199699|ICD9CM|AB|89.45|Pacemaker rate check
C0199700|ICD9CM|PT|89.46|Artificial pacemaker artifact wave form check
C0199700|ICD9CM|AB|89.46|Pacemaker wave form chck
C0199701|ICD9CM|PT|89.47|Artificial pacemaker electrode impedance check
C0199701|ICD9CM|AB|89.47|Pacemaker impedance chck
C0199779|ICD9CM|PT|99.21|Injection of antibiotic
C0199779|ICD9CM|AB|99.21|Inject antibiotic
C0199782|ICD9CM|PT|99.17|Injection of insulin
C0199782|ICD9CM|AB|99.17|Inject insulin
C0199783|ICD9CM|PT|99.26|Injection of tranquilizer
C0199783|ICD9CM|AB|99.26|Inject tranquilizer
C0199789|ICD9CM|PT|99.56|Administration of tetanus antitoxin
C0199789|ICD9CM|AB|99.56|Tetanus antitoxin admini
C0199791|ICD9CM|PT|99.57|Administration of botulism antitoxin
C0199791|ICD9CM|AB|99.57|Botulism antitoxin admin
C0199795|ICD9CM|PT|99.19|Injection of anticoagulant
C0199795|ICD9CM|AB|99.19|Inject anticoagulant
C0199804|ICD9CM|PT|99.33|Vaccination against tuberculosis
C0199804|ICD9CM|AB|99.33|Tuberculosis vaccination
C0199806|ICD9CM|PT|99.36|Administration of diphtheria toxoid
C0199806|ICD9CM|AB|99.36|Diphtheria toxoid admin
C0199807|ICD9CM|PT|99.38|Administration of tetanus toxoid
C0199807|ICD9CM|AB|99.38|Tetanus toxoid administ
C0199809|ICD9CM|PT|99.41|Administration of poliomyelitis vaccine
C0199809|ICD9CM|AB|99.41|Polio vaccine administra
C0199810|ICD9CM|PT|99.48|Administration of measles-mumps-rubella vaccine
C0199810|ICD9CM|AB|99.48|Mmr administration
C0199821|ICD9CM|PT|99.53|Prophylactic vaccination against arthropod-borne viral encephalitis
C0199821|ICD9CM|AB|99.53|Arbovirus enceph vaccin
C0199822|ICD9CM|PT|99.51|Prophylactic vaccination against the common cold
C0199822|ICD9CM|AB|99.51|Common cold vaccination
C0199823|ICD9CM|PT|99.43|Vaccination against yellow fever
C0199823|ICD9CM|AB|99.43|Yellow fever vaccination
C0199824|ICD9CM|PT|99.13|Immunization for autoimmune disease
C0199824|ICD9CM|AB|99.13|Autoimmune dis immunizat
C0199851|ICD9CM|PT|89.36|Manual examination of breast
C0199851|ICD9CM|AB|89.36|Manual exam of breast
C0199873|ICD9CM|AB|89.32|Esophageal manometry
C0199873|ICD9CM|PT|89.32|Esophageal manometry
C0199885|ICD9CM|PT|89.33|Digital examination of enterostomy stoma
C0199885|ICD9CM|AB|89.33|Digital enterostomy exam
C0199901|ICD9CM|PT|96.38|Removal of impacted feces
C0199901|ICD9CM|AB|96.38|Impacted feces removal
C0199911|ICD9CM|PT|51.15|Pressure measurement of sphincter of Oddi
C0199911|ICD9CM|AB|51.15|Sphinct of oddi measure
C0199964|ICD9CM|PT|99.08|Transfusion of blood expander
C0199964|ICD9CM|AB|99.08|Blood expander transfus
C0199967|ICD9CM|PT|99.06|Transfusion of coagulation factors
C0199967|ICD9CM|AB|99.06|Coag factor transfusion
C0199995|ICD9CM|AB|89.21|Urinary manometry
C0199995|ICD9CM|PT|89.21|Urinary manometry
C0200000|ICD9CM|AB|89.22|Cystometrogram
C0200000|ICD9CM|PT|89.22|Cystometrogram
C0200005|ICD9CM|PT|89.25|Urethral pressure profile [UPP]
C0200005|ICD9CM|AB|89.25|Urethral pressure profil
C0200007|ICD9CM|PT|89.23|Urethral sphincter electromyogram
C0200007|ICD9CM|AB|89.23|Urethral sphincter emg
C0200008|ICD9CM|AB|89.24|Uroflowmetry
C0200008|ICD9CM|PT|89.24|Uroflowmetry [UFR]
C0200038|ICD9CM|HT|68.1|Diagnostic procedures on uterus and supporting structures
C0200044|ICD9CM|PT|89.26|Gynecological examination
C0200044|ICD9CM|AB|89.26|Gynecologic examination
C0200066|ICD9CM|PT|73.4|Medical induction of labor
C0200066|ICD9CM|AB|73.4|Medical induction labor
C0200078|ICD9CM|PT|89.16|Transillumination of newborn skull
C0200078|ICD9CM|AB|89.16|Skull transilluminat
C0200104|ICD9CM|PT|89.19|Video and radio-telemetered electroencephalographic monitoring
C0200104|ICD9CM|AB|89.19|Video/radio eeg monitor
C0200149|ICD9CM|AB|95.09|Eye examination NOS
C0200149|ICD9CM|PT|95.09|Eye examination, not otherwise specified
C0200153|ICD9CM|AB|95.01|Limited eye examination
C0200153|ICD9CM|PT|95.01|Limited eye examination
C0200154|ICD9CM|PT|95.02|Comprehensive eye examination
C0200154|ICD9CM|PT|95.03|Extended ophthalmologic work-up
C0200154|ICD9CM|AB|95.03|Extended ophthal work-up
C0200154|ICD9CM|AB|95.02|Comprehensive eye exam
C0200156|ICD9CM|PT|95.04|Eye examination under anesthesia
C0200156|ICD9CM|AB|95.04|Anesthetized eye exam
C0200159|ICD9CM|AB|95.06|Color vision study
C0200159|ICD9CM|PT|95.06|Color vision study
C0200161|ICD9CM|AB|95.07|Dark adaptation study
C0200161|ICD9CM|PT|95.07|Dark adaptation study
C0200166|ICD9CM|PT|95.36|Ophthalmologic counseling and instruction
C0200166|ICD9CM|AB|95.36|Ophth counsel & instruct
C0200189|ICD9CM|AB|95.11|Fundus photography
C0200189|ICD9CM|PT|95.11|Fundus photography
C0200202|ICD9CM|AB|95.15|Ocular motility study
C0200202|ICD9CM|PT|95.15|Ocular motility study
C0200204|ICD9CM|AB|95.25|Electromyogram of eye
C0200204|ICD9CM|PT|95.25|Electromyogram of eye [EMG]
C0200223|ICD9CM|PT|95.31|Fitting and dispensing of spectacles
C0200223|ICD9CM|AB|95.31|Spectacle fit & dispense
C0200245|ICD9CM|AB|95.35|Orthoptic training
C0200245|ICD9CM|PT|95.35|Orthoptic training
C0200297|ICD9CM|AB|95.43|Audiological evaluation
C0200297|ICD9CM|PT|95.43|Audiological evaluation
C0200318|ICD9CM|AB|95.48|Fitting of hearing aid
C0200318|ICD9CM|PT|95.48|Fitting of hearing aid
C0200949|ICD9CM|AB|90.52|Culture-blood
C0200949|ICD9CM|PT|90.52|Microscopic examination of blood, culture
C0202616|ICD9CM|PT|88.31|Skeletal series
C0202616|ICD9CM|AB|88.31|Skeletal series x-ray
C0202638|ICD9CM|AB|88.83|Bone thermography
C0202638|ICD9CM|PT|88.83|Bone thermography
C0202639|ICD9CM|AB|88.84|Muscle thermography
C0202639|ICD9CM|PT|88.84|Muscle thermography
C0202673|ICD9CM|AB|88.94|Mri musculoskeletal
C0202673|ICD9CM|PT|88.94|Magnetic resonance imaging of musculoskeletal
C0202678|ICD9CM|HT|87.0|Soft tissue x-ray of face, head, and neck
C0202691|ICD9CM|PT|87.03|Computerized axial tomography of head
C0202691|ICD9CM|AB|87.03|C.A.T. scan of head
C0202704|ICD9CM|AB|88.81|Cerebral thermography
C0202704|ICD9CM|PT|88.81|Cerebral thermography
C0202725|ICD9CM|PT|87.13|Temporomandibular contrast arthrogram
C0202725|ICD9CM|AB|87.13|Tm contrast arthrogram
C0202735|ICD9CM|PT|87.15|Contrast radiogram of sinus
C0202735|ICD9CM|AB|87.15|Contrast x-ray of sinus
C0202745|ICD9CM|AB|87.05|Contrast dacryocystogram
C0202745|ICD9CM|PT|87.05|Contrast dacryocystogram
C0202750|ICD9CM|PT|87.14|Contrast radiogram of orbit
C0202750|ICD9CM|AB|87.14|Contrast x-ray of orbit
C0202752|ICD9CM|AB|88.82|Ocular thermography
C0202752|ICD9CM|PT|88.82|Ocular thermography
C0202774|ICD9CM|PT|87.06|Contrast radiogram of nasopharynx
C0202774|ICD9CM|AB|87.06|Nasophary contrast x-ray
C0202777|ICD9CM|PT|87.11|Full-mouth x-ray of teeth
C0202777|ICD9CM|AB|87.11|Full-mouth x-ray
C0202784|ICD9CM|AB|87.44|Routine chest x-ray
C0202784|ICD9CM|PT|87.44|Routine chest x-ray, so described
C0202806|ICD9CM|AB|87.31|Endotracheal bronchogram
C0202806|ICD9CM|PT|87.31|Endotracheal bronchogram
C0202812|ICD9CM|AB|87.33|Mediastinal pneumogram
C0202812|ICD9CM|PT|87.33|Mediastinal pneumogram
C0202819|ICD9CM|PT|87.43|X-ray of ribs, sternum, and clavicle
C0202819|ICD9CM|AB|87.43|Rib/sternum/clavic x-ray
C0202823|ICD9CM|PT|87.41|Computerized axial tomography of thorax
C0202823|ICD9CM|AB|87.41|C.A.T. scan of thorax
C0202827|ICD9CM|PT|88.92|Magnetic resonance imaging of chest and myocardium
C0202827|ICD9CM|AB|88.92|Mri chest & heart
C0202830|ICD9CM|HT|87.3|Soft tissue x-ray of thorax
C0202842|ICD9CM|PT|88.03|Sinogram of abdominal wall
C0202842|ICD9CM|AB|88.03|Abdominal wall sinogram
C0202843|ICD9CM|PT|88.14|Retroperitoneal fistulogram
C0202843|ICD9CM|AB|88.14|Retroperiton fistulogram
C0202845|ICD9CM|PT|88.12|Pelvic gas contrast radiography
C0202845|ICD9CM|AB|88.12|Pelvic gas contrast xray
C0202851|ICD9CM|PT|88.58|Negative-contrast cardiac roentgenography
C0202851|ICD9CM|AB|88.58|Negatve-contr cardiogram
C0202856|ICD9CM|PT|88.52|Angiocardiography of right heart structures
C0202856|ICD9CM|AB|88.52|Rt heart angiocardiogram
C0202857|ICD9CM|PT|88.53|Angiocardiography of left heart structures
C0202857|ICD9CM|AB|88.53|Lt heart angiocardiogram
C0202858|ICD9CM|PT|88.54|Combined right and left heart angiocardiography
C0202858|ICD9CM|AB|88.54|Rt & lt heart angiocard
C0202860|ICD9CM|PT|88.55|Coronary arteriography using a single catheter
C0202860|ICD9CM|AB|88.55|Coronar arteriogr-1 cath
C0202861|ICD9CM|PT|88.56|Coronary arteriography using two catheters
C0202861|ICD9CM|AB|88.56|Coronar arteriogr-2 cath
C0202892|ICD9CM|PT|88.86|Blood vessel thermography
C0202892|ICD9CM|AB|88.86|Blood vessel thermograph
C0202910|ICD9CM|PT|88.43|Arteriography of pulmonary arteries
C0202910|ICD9CM|AB|88.43|Contr pulmon arteriogram
C0202930|ICD9CM|PT|88.45|Arteriography of renal arteries
C0202930|ICD9CM|AB|88.45|Contrast renal arteriogr
C0202952|ICD9CM|PT|88.68|Impedance phlebography
C0202952|ICD9CM|AB|88.68|Impedance phlebogram
C0202968|ICD9CM|PT|88.51|Angiocardiography of venae cavae
C0202968|ICD9CM|AB|88.51|Vena cav angiocardiogram
C0202989|ICD9CM|AB|87.08|Cervical lymphangiogram
C0202989|ICD9CM|PT|87.08|Cervical lymphangiogram
C0202990|ICD9CM|PT|87.34|Intrathoracic lymphangiogram
C0202990|ICD9CM|AB|87.34|Intrathor lymphangiogram
C0202991|ICD9CM|AB|88.04|Abdominal lymphangiogram
C0202991|ICD9CM|PT|88.04|Abdominal lymphangiogram
C0202999|ICD9CM|PT|88.34|Lymphangiogram of upper limb
C0202999|ICD9CM|AB|88.34|Upper limb lymphangiogrm
C0203002|ICD9CM|PT|88.36|Lymphangiogram of lower limb
C0203002|ICD9CM|AB|88.36|Lower limb lymphangiogrm
C0203032|ICD9CM|AB|88.85|Breast thermography
C0203032|ICD9CM|PT|88.85|Breast thermography
C0203036|ICD9CM|HT|87.8|X-ray of female genital organs
C0203038|ICD9CM|AB|87.81|X-ray of gravid uterus
C0203038|ICD9CM|PT|87.81|X-ray of gravid uterus
C0203040|ICD9CM|AB|87.84|Percutaneous hysterogram
C0203040|ICD9CM|PT|87.84|Percutaneous hysterogram
C0203057|ICD9CM|AB|87.62|Upper GI series
C0203057|ICD9CM|PT|87.62|Upper GI series
C0203065|ICD9CM|AB|87.61|Barium swallow
C0203065|ICD9CM|PT|87.61|Barium swallow
C0203075|ICD9CM|AB|87.64|Lower GI series
C0203075|ICD9CM|PT|87.64|Lower GI series
C0203082|ICD9CM|PT|87.52|Intravenous cholangiogram
C0203082|ICD9CM|AB|87.52|Intraven cholangiogram
C0203083|ICD9CM|PT|87.53|Intraoperative cholangiogram
C0203083|ICD9CM|AB|87.53|Intraoper cholangiogram
C0203101|ICD9CM|HT|87.7|X-ray of urinary system
C0203108|ICD9CM|AB|87.73|Intravenous pyelogram
C0203108|ICD9CM|PT|87.73|Intravenous pyelogram
C0203110|ICD9CM|AB|87.74|Retrograde pyelogram
C0203110|ICD9CM|PT|87.74|Retrograde pyelogram
C0203122|ICD9CM|PT|88.95|Magnetic resonance imaging of pelvis, prostate, and bladder
C0203122|ICD9CM|AB|88.95|Mri pelvis,prostate,blad
C0203125|ICD9CM|PT|87.76|Retrograde cystourethrogram
C0203125|ICD9CM|AB|87.76|Retrogr cystourethrogram
C0203139|ICD9CM|HT|87.2|X-ray of spine
C0203238|ICD9CM|PT|88.22|Skeletal x-ray of elbow and forearm
C0203238|ICD9CM|AB|88.22|Skel xray-elbow/forearm
C0203243|ICD9CM|PT|88.23|Skeletal x-ray of wrist and hand
C0203243|ICD9CM|AB|88.23|Skel xray-wrist & hand
C0203286|ICD9CM|PT|88.28|Skeletal x-ray of ankle and foot
C0203286|ICD9CM|AB|88.28|Skel xray-ankle & foot
C0203407|ICD9CM|PT|88.75|Diagnostic ultrasound of urinary system
C0203407|ICD9CM|AB|88.75|Dx ultrasound-urinary
C0203419|ICD9CM|PT|88.78|Diagnostic ultrasound of gravid uterus
C0203419|ICD9CM|AB|88.78|Dx ultrasound-grav uter
C0203474|ICD9CM|PT|88.76|Diagnostic ultrasound of abdomen and retroperitoneum
C0203474|ICD9CM|AB|88.76|Dx ultrasound-abdomen
C0203541|ICD9CM|AB|92.22|Orthovoltage radiation
C0203541|ICD9CM|PT|92.22|Orthovoltage radiation
C0203598|ICD9CM|PT|99.85|Hyperthermia for treatment of cancer
C0203598|ICD9CM|AB|99.85|Hyperthermia ca therapy
C0203631|ICD9CM|PT|92.28|Injection or instillation of radioisotopes
C0203631|ICD9CM|AB|92.28|Isotope inject/instill
C0203668|ICD9CM|AB|92.14|Bone scan
C0203668|ICD9CM|PT|92.14|Bone scan
C0203669|ICD9CM|AB|92.18|Total body scan
C0203669|ICD9CM|PT|92.18|Total body scan
C0203683|ICD9CM|AB|92.15|Pulmonary scan
C0203683|ICD9CM|PT|92.15|Pulmonary scan
C0203779|ICD9CM|PT|92.01|Thyroid scan and radioisotope function studies
C0203779|ICD9CM|AB|92.01|Thyroid scan/isotop func
C0203792|ICD9CM|AB|92.13|Parathyroid scan
C0203792|ICD9CM|PT|92.13|Parathyroid scan
C0203879|ICD9CM|AB|92.17|Placental scan
C0203879|ICD9CM|PT|92.17|Placental scan
C0203886|ICD9CM|HT|93.0|Diagnostic physical therapy
C0203901|ICD9CM|PT|93.21|Manual and mechanical traction
C0203901|ICD9CM|AB|93.21|Manual & mechan traction
C0203909|ICD9CM|PT|93.38|Combined physical therapy without mention of the components
C0203909|ICD9CM|AB|93.38|Combined pt NOS
C0203910|ICD9CM|AB|93.07|Body measurement
C0203910|ICD9CM|PT|93.07|Body measurement
C0203922|ICD9CM|PT|93.06|Measurement of limb length
C0203922|ICD9CM|AB|93.06|Limb length measurement
C0203923|ICD9CM|PT|93.25|Forced extension of limb
C0203923|ICD9CM|AB|93.25|Forced limb extension
C0203924|ICD9CM|PT|93.26|Manual rupture of joint adhesions
C0203924|ICD9CM|AB|93.26|Manual rupt joint adhes
C0203938|ICD9CM|PT|93.64|Osteopathic manipulative treatment using isotonic, isometric forces
C0203938|ICD9CM|AB|93.64|Omt with isoton,isometri
C0203939|ICD9CM|PT|93.65|Osteopathic manipulative treatment using indirect forces
C0203939|ICD9CM|AB|93.65|Omt with indirect forces
C0203940|ICD9CM|PT|93.66|Osteopathic manipulative treatment to move tissue fluids
C0203940|ICD9CM|AB|93.66|Omt to move tissue fluid
C0203967|ICD9CM|AB|93.14|Joint movement training
C0203967|ICD9CM|PT|93.14|Training in joint movements
C0203968|ICD9CM|PT|93.22|Ambulation and gait training
C0203968|ICD9CM|AB|93.22|Ambulat & gait training
C0203981|ICD9CM|AB|93.36|Cardiac retraining
C0203981|ICD9CM|PT|93.36|Cardiac retraining
C0203989|ICD9CM|AB|93.11|Assisting exercise
C0203989|ICD9CM|PT|93.11|Assisting exercise
C0203991|ICD9CM|AB|93.13|Resistive exercise
C0203991|ICD9CM|PT|93.13|Resistive exercise
C0204026|ICD9CM|AB|93.32|Whirlpool treatment
C0204026|ICD9CM|PT|93.32|Whirlpool treatment
C0204051|ICD9CM|PT|93.04|Manual testing of muscle function
C0204051|ICD9CM|AB|93.04|Manual muscle funct test
C0204061|ICD9CM|AB|93.05|Range of motion testing
C0204061|ICD9CM|PT|93.05|Range of motion testing
C0204067|ICD9CM|AB|93.02|Orthotic evaluation
C0204067|ICD9CM|PT|93.02|Orthotic evaluation
C0204072|ICD9CM|PT|93.23|Fitting of orthotic device
C0204072|ICD9CM|AB|93.23|Orthotic device fitting
C0204077|ICD9CM|AB|93.03|Prosthetic evaluation
C0204077|ICD9CM|PT|93.03|Prosthetic evaluation
C0204088|ICD9CM|AB|93.72|Dysphasia training
C0204088|ICD9CM|PT|93.72|Dysphasia training
C0204089|ICD9CM|AB|93.74|Speech defect training
C0204089|ICD9CM|PT|93.74|Speech defect training
C0204090|ICD9CM|AB|93.71|Dyslexia training
C0204090|ICD9CM|PT|93.71|Dyslexia training
C0204093|ICD9CM|HT|93.3|Other physical therapy therapeutic procedures
C0204145|ICD9CM|PT|23.01|Extraction of deciduous tooth
C0204145|ICD9CM|AB|23.01|Deciduous tooth extract
C0204479|ICD9CM|HT|94|Procedures related to the psyche
C0204525|ICD9CM|HT|94.3|Individual psychotherapy
C0204540|ICD9CM|PT|94.38|Supportive verbal psychotherapy
C0204540|ICD9CM|AB|94.38|Suppor verbal psychother
C0204542|ICD9CM|PT|94.37|Exploratory verbal psychotherapy
C0204542|ICD9CM|AB|94.37|Explor verbal psychother
C0204583|ICD9CM|AB|93.82|Educational therapy
C0204583|ICD9CM|PT|93.82|Educational therapy
C0204589|ICD9CM|PT|94.26|Subconvulsive electroshock therapy
C0204589|ICD9CM|AB|94.26|Subconvulsive est
C0204592|ICD9CM|AB|94.22|Lithium therapy
C0204592|ICD9CM|PT|94.22|Lithium therapy
C0204597|ICD9CM|AB|94.62|Alcohol detoxification
C0204597|ICD9CM|PT|94.62|Alcohol detoxification
C0204598|ICD9CM|AB|94.61|Alcohol rehabilitation
C0204598|ICD9CM|PT|94.61|Alcohol rehabilitation
C0204599|ICD9CM|PT|94.63|Alcohol rehabilitation and detoxification
C0204599|ICD9CM|AB|94.63|Alcohol rehab/detox
C0204600|ICD9CM|AB|94.65|Drug detoxification
C0204600|ICD9CM|PT|94.65|Drug detoxification
C0204601|ICD9CM|AB|94.64|Drug rehabilitation
C0204601|ICD9CM|PT|94.64|Drug rehabilitation
C0204602|ICD9CM|PT|94.66|Drug rehabilitation and detoxification
C0204602|ICD9CM|AB|94.66|Drug rehab/detox
C0204603|ICD9CM|PT|94.68|Combined alcohol and drug detoxification
C0204603|ICD9CM|AB|94.68|Comb alcohol/drug detox
C0204604|ICD9CM|PT|94.67|Combined alcohol and drug rehabilitation
C0204604|ICD9CM|AB|94.67|Comb alcohol/drug rehab
C0204605|ICD9CM|PT|94.69|Combined alcohol and drug rehabilitation and detoxification
C0204605|ICD9CM|AB|94.69|Comb alco/drug reha/deto
C0204727|ICD9CM|AB|99.84|Isolation
C0204727|ICD9CM|PT|99.84|Isolation
C0204785|ICD9CM|AB|96.44|Vaginal douche
C0204785|ICD9CM|PT|96.44|Vaginal douche
C0204786|ICD9CM|PT|97.71|Removal of intrauterine contraceptive device
C0204786|ICD9CM|AB|97.71|Removal iud
C0204816|ICD9CM|PT|97.23|Replacement of tracheostomy tube
C0204816|ICD9CM|AB|97.23|Replace trach tube
C0204854|ICD9CM|AB|81.91|Arthrocentesis
C0204854|ICD9CM|PT|81.91|Arthrocentesis
C0204861|ICD9CM|AB|93.54|Application of splint
C0204861|ICD9CM|PT|93.54|Application of splint
C0204916|ICD9CM|PT|89.64|Pulmonary artery wedge monitoring
C0204916|ICD9CM|AB|89.64|Pulmon art wedge monitor
C0205792|ICD9CM|PT|618.6|Vaginal enterocele, congenital or acquired
C0205792|ICD9CM|AB|618.6|Vaginal enterocele
C0205858|ICD9CM|AB|094.1|General paresis
C0205858|ICD9CM|PT|094.1|General paresis
C0205929|ICD9CM|AB|565.1|Anal fistula
C0205929|ICD9CM|PT|565.1|Anal fistula
C0205930|ICD9CM|AB|733.7|Algoneurodystrophy
C0205930|ICD9CM|PT|733.7|Algoneurodystrophy
C0206042|ICD9CM|PT|046.72|Fatal familial insomnia
C0206042|ICD9CM|AB|046.72|Fatal familial insomnia
C0206078|ICD9CM|PT|80.51|Excision of intervertebral disc
C0206078|ICD9CM|AB|80.51|Excision intervert disc
C0206180|ICD9CM|HT|200.6|Anaplastic large cell lymphoma
C0206368|ICD9CM|PT|365.52|Pseudoexfoliation glaucoma
C0206368|ICD9CM|AB|365.52|Pseudoexfoliat glaucoma
C0206373|ICD9CM|PT|99.88|Therapeutic photopheresis
C0206373|ICD9CM|AB|99.88|Therapeutc photopheresis
C0206504|ICD9CM|HT|384.2|Perforation of tympanic membrane
C0206504|ICD9CM|PT|384.20|Perforation of tympanic membrane, unspecified
C0206504|ICD9CM|AB|384.20|Perforat tympan memb NOS
C0206754|ICD9CM|HT|209-209.99|NEUROENDOCRINE TUMORS
C0206754|ICD9CM|HT|209|Neuroendocrine tumors
C0206762|ICD9CM|PT|755.9|Unspecified anomaly of unspecified limb
C0206762|ICD9CM|AB|755.9|Congen limb anomaly NOS
C0220636|ICD9CM|PT|142.9|Malignant neoplasm of salivary gland, unspecified
C0220636|ICD9CM|AB|142.9|Mal neo salivary NOS
C0220656|ICD9CM|PT|789.51|Malignant ascites
C0220656|ICD9CM|AB|789.51|Malignant ascites
C0220704|ICD9CM|PT|758.32|Velo-cardio-facial syndrome
C0220704|ICD9CM|AB|758.32|Velo-cardio-facial synd
C0220887|ICD9CM|HT|666.1|Other immediate postpartum hemorrhage
C0220887|ICD9CM|PT|666.14|Other immediate postpartum hemorrhage, postpartum condition or complication
C0220887|ICD9CM|AB|666.14|Postpart hem NEC-postpar
C0220977|ICD9CM|HT|115.1|Infection by Histoplasma duboisii
C0221002|ICD9CM|PT|252.01|Primary hyperparathyroidism
C0221002|ICD9CM|AB|252.01|Primary hyperparathyroid
C0221023|ICD9CM|PT|288.02|Cyclic neutropenia
C0221023|ICD9CM|AB|288.02|Cyclic neutropenia
C0221046|ICD9CM|PT|337.01|Carotid sinus syndrome
C0221046|ICD9CM|AB|337.01|Carotid sinus syndrome
C0221103|ICD9CM|PT|368.31|Suppression of binocular vision
C0221103|ICD9CM|AB|368.31|Binocular vis suppress
C0221217|ICD9CM|AB|744.5|Webbing of neck
C0221217|ICD9CM|PT|744.5|Webbing of neck
C0221244|ICD9CM|AB|690.11|Seborrhea capitis
C0221244|ICD9CM|PT|690.11|Seborrhea capitis
C0221352|ICD9CM|PT|755.11|Syndactyly of fingers without fusion of bone
C0221352|ICD9CM|AB|755.11|Syndactyl fing-no fusion
C0221468|ICD9CM|AB|268.0|Rickets, active
C0221468|ICD9CM|PT|268.0|Rickets, active
C0221520|ICD9CM|HT|295.0|Simple type schizophrenia
C0221520|ICD9CM|PT|295.00|Simple type schizophrenia, unspecified
C0221520|ICD9CM|AB|295.00|Simpl schizophren-unspec
C0221539|ICD9CM|PT|780.02|Transient alteration of awareness
C0221539|ICD9CM|AB|780.02|Trans alter awareness
C0221540|ICD9CM|PT|780.09|Other alteration of consciousness
C0221540|ICD9CM|AB|780.09|Other alter consciousnes
C0221565|ICD9CM|PT|V17.7|Family history of arthritis
C0221565|ICD9CM|AB|V17.7|Family hx-arthritis
C0221757|ICD9CM|PT|273.4|Alpha-1-antitrypsin deficiency
C0221757|ICD9CM|AB|273.4|Alpha-1-antitrypsin def
C0231311|ICD9CM|PT|327.35|Circadian rhythm sleep disorder, jet lag type
C0231311|ICD9CM|AB|327.35|Circadian rhythm-jetlag
C0231471|ICD9CM|AB|781.92|Abnormal posture
C0231471|ICD9CM|PT|781.92|Abnormal posture
C0231666|ICD9CM|AB|736.05|Wrist drop
C0231666|ICD9CM|PT|736.05|Wrist drop (acquired)
C0231835|ICD9CM|AB|786.06|Tachypnea
C0231835|ICD9CM|PT|786.06|Tachypnea
C0232286|ICD9CM|AB|786.51|Precordial pain
C0232286|ICD9CM|PT|786.51|Precordial pain
C0232488|ICD9CM|PT|789.7|Colic
C0232488|ICD9CM|AB|789.7|Colic
C0232493|ICD9CM|PT|789.06|Abdominal pain, epigastric
C0232493|ICD9CM|AB|789.06|Abdmnal pain epigastric
C0232498|ICD9CM|HT|789.6|Abdominal tenderness
C0232498|ICD9CM|PT|789.60|Abdominal tenderness, unspecified site
C0232498|ICD9CM|AB|789.60|Abdmnal tndr unspcf site
C0232599|ICD9CM|AB|787.04|Bilious emesis
C0232599|ICD9CM|PT|787.04|Bilious emesis
C0232854|ICD9CM|PT|788.62|Slowing of urinary stream
C0232854|ICD9CM|AB|788.62|Slowing urinary stream
C0232855|ICD9CM|PT|788.61|Splitting of urinary stream
C0232855|ICD9CM|AB|788.61|Splitting urinary stream
C0232857|ICD9CM|AB|306.53|Psychogenic dysuria
C0232857|ICD9CM|PT|306.53|Psychogenic dysuria
C0232867|ICD9CM|AB|593.6|Postural proteinuria
C0232867|ICD9CM|PT|593.6|Postural proteinuria
C0233757|ICD9CM|AB|307.54|Psychogenic vomiting
C0233757|ICD9CM|PT|307.54|Psychogenic vomiting
C0233880|ICD9CM|PT|302.0|Ego-dystonic sexual orientation
C0233880|ICD9CM|AB|302.0|Ego-dystonic sex orient
C0234398|ICD9CM|HT|377.7|Disorders of visual cortex
C0234428|ICD9CM|HT|780.0|Alteration of consciousness
C0235029|ICD9CM|PT|997.00|Nervous system complication, unspecified
C0235029|ICD9CM|AB|997.00|Nervous syst complc NOS
C0235065|ICD9CM|PT|770.87|Respiratory arrest of newborn
C0235065|ICD9CM|AB|770.87|NB respiratory arrest
C0235093|ICD9CM|AB|596.53|Paralysis of bladder
C0235093|ICD9CM|PT|596.53|Paralysis of bladder
C0235238|ICD9CM|AB|367.51|Paresis of accommodation
C0235238|ICD9CM|PT|367.51|Paresis of accommodation
C0235299|ICD9CM|PT|789.01|Abdominal pain, right upper quadrant
C0235299|ICD9CM|AB|789.01|Abdmnal pain rt upr quad
C0235326|ICD9CM|PT|455.7|Unspecified thrombosed hemorrhoids
C0235326|ICD9CM|AB|455.7|Thrombos hemorrhoids NOS
C0235604|ICD9CM|PT|287.1|Qualitative platelet defects
C0235604|ICD9CM|AB|287.1|Thrombocytopathy
C0235653|ICD9CM|HT|174|Malignant neoplasm of female breast
C0235653|ICD9CM|PT|174.9|Malignant neoplasm of breast (female), unspecified
C0235653|ICD9CM|AB|174.9|Malign neopl breast NOS
C0235660|ICD9CM|PT|611.6|Galactorrhea not associated with childbirth
C0235660|ICD9CM|AB|611.6|Galactorrhea-nonobstet
C0235756|ICD9CM|PT|792.2|Nonspecific abnormal findings in semen
C0235756|ICD9CM|AB|792.2|Abn findings-semen
C0235815|ICD9CM|PT|771.82|Urinary tract infection of newborn
C0235815|ICD9CM|AB|771.82|NB urinary tract infectn
C0235880|ICD9CM|AB|355.9|Mononeuritis NOS
C0235880|ICD9CM|PT|355.9|Mononeuritis of unspecified site
C0235904|ICD9CM|PT|564.7|Megacolon, other than Hirschsprung's
C0235904|ICD9CM|AB|564.7|Megacolon NEC
C0235963|ICD9CM|PT|478.11|Nasal mucositis (ulcerative)
C0235963|ICD9CM|AB|478.11|Nasal mucositis (ulcer)
C0236000|ICD9CM|PT|784.92|Jaw pain
C0236000|ICD9CM|AB|784.92|Jaw pain
C0236127|ICD9CM|PT|530.21|Ulcer of esophagus with bleeding
C0236127|ICD9CM|AB|530.21|Ulcer esophagus w bleed
C0236140|ICD9CM|PT|794.31|Nonspecific abnormal electrocardiogram [ECG] [EKG]
C0236140|ICD9CM|AB|794.31|Abnorm electrocardiogram
C0236151|ICD9CM|PT|794.4|Nonspecific abnormal results of function study of kidney
C0236151|ICD9CM|AB|794.4|Abn kidney funct study
C0236642|ICD9CM|AB|331.11|Pick's disease
C0236642|ICD9CM|PT|331.11|Pick's disease
C0236650|ICD9CM|PT|290.40|Vascular dementia, uncomplicated
C0236650|ICD9CM|AB|290.40|Vascular dementia,uncomp
C0236651|ICD9CM|PT|290.41|Vascular dementia, with delirium
C0236651|ICD9CM|AB|290.41|Vasc dementia w delirium
C0236652|ICD9CM|PT|290.42|Vascular dementia, with delusions
C0236652|ICD9CM|AB|290.42|Vasc dementia w delusion
C0236653|ICD9CM|PT|290.43|Vascular dementia, with depressed mood
C0236653|ICD9CM|AB|290.43|Vasc dementia w depressn
C0236656|ICD9CM|PT|291.2|Alcohol-induced persisting dementia
C0236656|ICD9CM|AB|291.2|Alcohol persist dementia
C0236658|ICD9CM|PT|291.5|Alcohol-induced psychotic disorder with delusions
C0236658|ICD9CM|AB|291.5|Alcoh psych dis w delus
C0236662|ICD9CM|PT|291.82|Alcohol induced sleep disorders
C0236662|ICD9CM|AB|291.82|Alcoh induce sleep disor
C0236663|ICD9CM|AB|291.81|Alcohol withdrawal
C0236663|ICD9CM|PT|291.81|Alcohol withdrawal
C0236756|ICD9CM|PT|296.00|Bipolar I disorder, single manic episode, unspecified
C0236756|ICD9CM|HT|296.0|Bipolar I disorder, single manic episode
C0236756|ICD9CM|AB|296.00|Bipol I single manic NOS
C0236757|ICD9CM|PT|296.01|Bipolar I disorder, single manic episode, mild
C0236757|ICD9CM|AB|296.01|Bipol I single manc-mild
C0236758|ICD9CM|PT|296.02|Bipolar I disorder, single manic episode, moderate
C0236758|ICD9CM|AB|296.02|Bipol I single manic-mod
C0236762|ICD9CM|PT|296.06|Bipolar I disorder, single manic episode, in full remission
C0236762|ICD9CM|AB|296.06|Bipol I single manic rem
C0236773|ICD9CM|PT|296.50|Bipolar I disorder, most recent episode (or current) depressed, unspecified
C0236773|ICD9CM|AB|296.50|Bipol I cur depres NOS
C0236780|ICD9CM|PT|296.60|Bipolar I disorder, most recent episode (or current) mixed, unspecified
C0236780|ICD9CM|AB|296.60|Bipol I currnt mixed NOS
C0236791|ICD9CM|HT|299.1|Childhood disintegrative disorder
C0236794|ICD9CM|PT|300.01|Panic disorder without agoraphobia
C0236794|ICD9CM|AB|300.01|Panic dis w/o agorphobia
C0236795|ICD9CM|AB|300.12|Dissociative amnesia
C0236795|ICD9CM|PT|300.12|Dissociative amnesia
C0236800|ICD9CM|PT|300.21|Agoraphobia with panic disorder
C0236800|ICD9CM|AB|300.21|Agoraphobia w panic dis
C0236802|ICD9CM|PT|302.6|Gender identity disorder in children
C0236802|ICD9CM|AB|302.6|Gendr identity dis-child
C0236816|ICD9CM|HT|308|Acute reaction to stress
C0236816|ICD9CM|PT|308.9|Unspecified acute reaction to stress
C0236816|ICD9CM|AB|308.9|Acute stress react NOS
C0236826|ICD9CM|PT|315.31|Expressive language disorder
C0236826|ICD9CM|AB|315.31|Expressive language dis
C0236827|ICD9CM|PT|315.32|Mixed receptive-expressive language disorder
C0236827|ICD9CM|AB|315.32|Recp-expres language dis
C0236859|ICD9CM|AB|995.81|Adult physical abuse
C0236859|ICD9CM|PT|995.81|Adult physical abuse
C0236860|ICD9CM|AB|995.83|Adult sexual abuse
C0236860|ICD9CM|PT|995.83|Adult sexual abuse
C0236861|ICD9CM|AB|995.54|Child physical abuse
C0236861|ICD9CM|PT|995.54|Child physical abuse
C0236989|ICD9CM|HT|302|Sexual and gender identity disorders
C0238009|ICD9CM|PT|036.82|Meningococcal arthropathy
C0238009|ICD9CM|AB|036.82|Meningococc arthropathy
C0238015|ICD9CM|AB|337.3|Autonomic dysreflexia
C0238015|ICD9CM|PT|337.3|Autonomic dysreflexia
C0238027|ICD9CM|PT|040.41|Infant botulism
C0238027|ICD9CM|AB|040.41|Infant botulism
C0238074|ICD9CM|HT|416|Chronic pulmonary heart disease
C0238074|ICD9CM|PT|416.9|Chronic pulmonary heart disease, unspecified
C0238074|ICD9CM|AB|416.9|Chr pulmon heart dis NOS
C0238124|ICD9CM|AB|728.86|Necrotizing fasciitis
C0238124|ICD9CM|PT|728.86|Necrotizing fasciitis
C0238190|ICD9CM|AB|359.71|Inclusion body myositis
C0238190|ICD9CM|PT|359.71|Inclusion body myositis
C0238378|ICD9CM|PT|516.37|Desquamative interstitial pneumonia
C0238378|ICD9CM|PT|516.34|Respiratory bronchiolitis interstitial lung disease
C0238378|ICD9CM|AB|516.37|Desquamatv interst pneu
C0238378|ICD9CM|AB|516.34|Resp brncio interst lung
C0238425|ICD9CM|PT|282.62|Hb-SS disease with crisis
C0238425|ICD9CM|AB|282.62|Hb-SS disease w crisis
C0238502|ICD9CM|AB|618.03|Urethrocele
C0238502|ICD9CM|PT|618.03|Urethrocele
C0238528|ICD9CM|PT|008.44|Intestinal infection due to yersinia enterocolitica
C0238528|ICD9CM|AB|008.44|Int inf yrsnia entrcltca
C0238551|ICD9CM|PT|789.04|Abdominal pain, left lower quadrant
C0238551|ICD9CM|AB|789.04|Abdmnal pain lt lwr quad
C0238552|ICD9CM|PT|789.02|Abdominal pain, left upper quadrant
C0238552|ICD9CM|AB|789.02|Abdmnal pain lft up quad
C0238566|ICD9CM|PT|789.62|Abdominal tenderness, left upper quadrant
C0238566|ICD9CM|AB|789.62|Abdmnal tndr lft up quad
C0238570|ICD9CM|PT|789.63|Abdominal tenderness, right lower quadrant
C0238570|ICD9CM|AB|789.63|Abdmnal tndr rt lwr quad
C0238571|ICD9CM|PT|789.61|Abdominal tenderness, right upper quadrant
C0238571|ICD9CM|AB|789.61|Abdmnal tndr rt upr quad
C0238875|ICD9CM|PT|795.82|Elevated cancer antigen 125 [CA 125]
C0238875|ICD9CM|AB|795.82|Elev ca antigen 125
C0239167|ICD9CM|AB|787.61|Incomplete defecation
C0239167|ICD9CM|PT|787.61|Incomplete defecation
C0239233|ICD9CM|AB|780.94|Early satiety
C0239233|ICD9CM|PT|780.94|Early satiety
C0239280|ICD9CM|PT|789.66|Abdominal tenderness, epigastric
C0239280|ICD9CM|AB|789.66|Abdmnal tndr epigastric
C0239293|ICD9CM|AB|530.82|Esophageal hemorrhage
C0239293|ICD9CM|PT|530.82|Esophageal hemorrhage
C0239295|ICD9CM|AB|112.84|Candidal esophagitis
C0239295|ICD9CM|PT|112.84|Candidal esophagitis
C0239937|ICD9CM|PT|599.72|Microscopic hematuria
C0239937|ICD9CM|AB|599.72|Microscopic hematuria
C0240310|ICD9CM|AB|524.03|Maxillary hypoplasia
C0240310|ICD9CM|PT|524.03|Major anomalies of jaw size, maxillary hypoplasia
C0240802|ICD9CM|AB|V72.42|Pregnancy test-positive
C0240802|ICD9CM|PT|V72.42|Pregnancy examination or test, positive result
C0240896|ICD9CM|AB|743.52|Fundus coloboma
C0240896|ICD9CM|PT|743.52|Fundus coloboma
C0241790|ICD9CM|PT|747.32|Pulmonary arteriovenous malformation
C0241790|ICD9CM|AB|747.32|Pulmonary AV malformatn
C0241910|ICD9CM|AB|571.42|Autoimmune hepatitis
C0241910|ICD9CM|PT|571.42|Autoimmune hepatitis
C0242172|ICD9CM|PT|614.9|Unspecified inflammatory disease of female pelvic organs and tissues
C0242172|ICD9CM|HT|614-616.99|INFLAMMATORY DISEASE OF FEMALE PELVIC ORGANS
C0242172|ICD9CM|AB|614.9|Fem pelv inflam dis NOS
C0242225|ICD9CM|HT|368.5|Color vision deficiencies
C0242343|ICD9CM|AB|253.2|Panhypopituitarism
C0242343|ICD9CM|PT|253.2|Panhypopituitarism
C0242383|ICD9CM|AB|362.50|Macular degeneration NOS
C0242383|ICD9CM|PT|362.50|Macular degeneration (senile), unspecified
C0242407|ICD9CM|PT|429.82|Hyperkinetic heart disease
C0242407|ICD9CM|AB|429.82|Hyperkinetic heart dis
C0242420|ICD9CM|AB|362.83|Retinal edema
C0242420|ICD9CM|PT|362.83|Retinal edema
C0242427|ICD9CM|AB|37.12|Pericardiotomy
C0242427|ICD9CM|PT|37.12|Pericardiotomy
C0242429|ICD9CM|AB|784.1|Throat pain
C0242429|ICD9CM|PT|784.1|Throat pain
C0242490|ICD9CM|PT|726.90|Enthesopathy of unspecified site
C0242490|ICD9CM|HT|726.9|Unspecified enthesopathy
C0242490|ICD9CM|AB|726.90|Enthesopathy, site NOS
C0242670|ICD9CM|PT|780.03|Persistent vegetative state
C0242670|ICD9CM|AB|780.03|Persistent vegtv state
C0242770|ICD9CM|PT|516.36|Cryptogenic organizing pneumonia
C0242770|ICD9CM|AB|516.36|Cryptogenic organiz pneu
C0242787|ICD9CM|HT|175|Malignant neoplasm of male breast
C0242855|ICD9CM|PT|746.01|Atresia of pulmonary valve, congenital
C0242855|ICD9CM|AB|746.01|Cong pulmon valv atresia
C0242966|ICD9CM|AB|995.90|SIRS, NOS
C0242966|ICD9CM|HT|995.9|Systemic inflammatory response syndrome (SIRS)
C0242966|ICD9CM|PT|995.90|Systemic inflammatory response syndrome, unspecified
C0243026|ICD9CM|PT|995.91|Sepsis
C0243026|ICD9CM|AB|995.91|Sepsis
C0259768|ICD9CM|HT|998.3|Disruption of wound
C0259768|ICD9CM|AB|998.30|Wound disruption NOS
C0259768|ICD9CM|PT|998.30|Disruption of wound, unspecified
C0259797|ICD9CM|AB|E906.0|Dog bite
C0259797|ICD9CM|PT|E906.0|Dog bite
C0259799|ICD9CM|AB|370.21|Punctate keratitis
C0259799|ICD9CM|PT|370.21|Punctate keratitis
C0259800|ICD9CM|HT|360.0|Purulent endophthalmitis
C0259800|ICD9CM|PT|360.00|Purulent endophthalmitis, unspecified
C0259800|ICD9CM|AB|360.00|Purulent endophthalm NOS
C0260334|ICD9CM|AB|507.0|Food/vomit pneumonitis
C0260334|ICD9CM|PT|507.0|Pneumonitis due to inhalation of food or vomitus
C0260335|ICD9CM|HT|636.9|Illegally induced abortion without mention of complication
C0260335|ICD9CM|PT|636.90|Illegally induced abortion, without mention of complication, unspecified
C0260335|ICD9CM|AB|636.90|Illeg abort uncompl-unsp
C0260338|ICD9CM|HT|642.6|Eclampsia complicating pregnancy, childbirth or the puerperium
C0260339|ICD9CM|HT|V01|Contact with or exposure to communicable diseases
C0260339|ICD9CM|PT|V01.9|Contact with or exposure to unspecified communicable disease
C0260339|ICD9CM|AB|V01.9|Communic dis contact NOS
C0260340|ICD9CM|PT|V01.0|Contact with or exposure to cholera
C0260340|ICD9CM|AB|V01.0|Cholera contact
C0260341|ICD9CM|PT|V01.1|Contact with or exposure to tuberculosis
C0260341|ICD9CM|AB|V01.1|Tuberculosis contact
C0260342|ICD9CM|PT|V01.2|Contact with or exposure to poliomyelitis
C0260342|ICD9CM|AB|V01.2|Poliomyelitis contact
C0260343|ICD9CM|PT|V01.3|Contact with or exposure to smallpox
C0260343|ICD9CM|AB|V01.3|Smallpox contact
C0260344|ICD9CM|PT|V01.4|Contact with or exposure to rubella
C0260344|ICD9CM|AB|V01.4|Rubella contact
C0260345|ICD9CM|PT|V01.5|Contact with or exposure to rabies
C0260345|ICD9CM|AB|V01.5|Rabies contact
C0260346|ICD9CM|PT|V01.6|Contact with or exposure to venereal diseases
C0260346|ICD9CM|AB|V01.6|Venereal dis contact
C0260347|ICD9CM|HT|V01.7|Contact with or exposure to other viral diseases
C0260347|ICD9CM|PT|V01.79|Contact with or exposure to other viral diseases
C0260347|ICD9CM|AB|V01.79|Viral dis contact NEC
C0260348|ICD9CM|HT|V01.8|Contact with or exposure to other communicable diseases
C0260348|ICD9CM|PT|V01.89|Contact with or exposure to other communicable diseases
C0260348|ICD9CM|AB|V01.89|Communic dis contact NEC
C0260351|ICD9CM|PT|V02.0|Carrier or suspected carrier of cholera
C0260351|ICD9CM|AB|V02.0|Cholera carrier
C0260352|ICD9CM|PT|V02.1|Carrier or suspected carrier of typhoid
C0260352|ICD9CM|AB|V02.1|Typhoid carrier
C0260354|ICD9CM|PT|V02.3|Carrier or suspected carrier of other gastrointestinal pathogens
C0260354|ICD9CM|AB|V02.3|GI pathogen carrier NEC
C0260355|ICD9CM|PT|V02.4|Carrier or suspected carrier of diphtheria
C0260355|ICD9CM|AB|V02.4|Diphtheria carrier
C0260356|ICD9CM|HT|V02.5|Carrier or suspected carrier of other specified bacterial diseases
C0260356|ICD9CM|PT|V02.59|Carrier or suspected carrier of other specified bacterial diseases
C0260356|ICD9CM|AB|V02.59|Bacteria dis carrier NEC
C0260359|ICD9CM|PT|V02.8|Carrier or suspected carrier of other venereal diseases
C0260359|ICD9CM|AB|V02.8|Venereal dis carrier NEC
C0260360|ICD9CM|PT|V02.9|Carrier or suspected carrier of other specified infectious organism
C0260360|ICD9CM|AB|V02.9|Carrier NEC
C0260361|ICD9CM|HT|V03|Need for prophylactic vaccination and inoculation against bacterial diseases
C0260362|ICD9CM|PT|V03.0|Need for prophylactic vaccination and inoculation against cholera alone
C0260362|ICD9CM|AB|V03.0|Vaccin for cholera
C0260363|ICD9CM|PT|V03.1|Need for prophylactic vaccination and inoculation against typhoid-paratyphoid alone [TAB]
C0260363|ICD9CM|AB|V03.1|Vacc-typhoid-paratyphoid
C0260364|ICD9CM|PT|V03.2|Need for prophylactic vaccination and inoculation against tuberculosis [BCG]
C0260364|ICD9CM|AB|V03.2|Vaccin for tuberculosis
C0260367|ICD9CM|PT|V03.5|Need for prophylactic vaccination and inoculation against diphtheria alone
C0260367|ICD9CM|AB|V03.5|Vaccin for diphtheria
C0260368|ICD9CM|PT|V03.6|Need for prophylactic vaccination and inoculation against pertussis alone
C0260368|ICD9CM|AB|V03.6|Vaccin for pertussis
C0260371|ICD9CM|PT|V03.9|Need for prophylactic vaccination and inoculation against unspecified single bacterial disease
C0260371|ICD9CM|AB|V03.9|Vaccin for bact dis NOS
C0260374|ICD9CM|PT|V04.1|Need for prophylactic vaccination and inoculation against smallpox
C0260374|ICD9CM|AB|V04.1|Vaccin for smallpox
C0260380|ICD9CM|PT|V04.7|Need for prophylactic vaccination and inoculation against common cold
C0260380|ICD9CM|AB|V04.7|Vaccin for common cold
C0260384|ICD9CM|PT|V05.1|Need for prophylactic vaccination and inoculation against other arthropod-borne viral diseases
C0260384|ICD9CM|AB|V05.1|Vacc arboviral dis NEC
C0260386|ICD9CM|PT|V05.8|Need for prophylactic vaccination and inoculation against other specified disease
C0260386|ICD9CM|AB|V05.8|Vaccin for disease NEC
C0260387|ICD9CM|PT|V05.9|Need for prophylactic vaccination and inoculation against unspecified single disease
C0260387|ICD9CM|AB|V05.9|Vaccin for singl dis NOS
C0260388|ICD9CM|HT|V06|Need for prophylactic vaccination and inoculation against combinations of diseases
C0260389|ICD9CM|PT|V06.0|Need for prophylactic vaccination and inoculation against cholera with typhoid-paratyphoid [cholera + TAB]
C0260389|ICD9CM|AB|V06.0|Vaccin for cholera + tab
C0260390|ICD9CM|PT|V06.1|Need for prophylactic vaccination and inoculation against diphtheria-tetanus-pertussis, combined [DTP] [DTaP]
C0260390|ICD9CM|AB|V06.1|Vaccination for DTP-DTaP
C0260391|ICD9CM|PT|V06.2|Need for prophylactic vaccination and inoculation against diptheria-tetanus- pertussis with typhoid-paratyphoid (DTP + TAB)
C0260391|ICD9CM|AB|V06.2|Vaccin for dtp + tab
C0260392|ICD9CM|PT|V06.3|Need for prophylactic vaccination and inoculation against diptheria-tetanus- pertussis with poliomyelitis [DTP + polio]
C0260392|ICD9CM|AB|V06.3|Vaccin for dtp + polio
C0260394|ICD9CM|PT|V06.8|Need for prophylactic vaccination and inoculation against other combinations of diseases
C0260394|ICD9CM|AB|V06.8|Vac-dis combinations NEC
C0260395|ICD9CM|PT|V06.9|Unspecified combined vaccine
C0260395|ICD9CM|AB|V06.9|Vac-dis combinations NOS
C0260397|ICD9CM|PT|V07.0|Need for isolation
C0260397|ICD9CM|AB|V07.0|Prophylactic isolation
C0260398|ICD9CM|PT|V07.1|Need for desensitization to allergens
C0260398|ICD9CM|AB|V07.1|Desensitiza to allergens
C0260399|ICD9CM|PT|V07.2|Need for prophylactic immunotherapy
C0260399|ICD9CM|AB|V07.2|Prophylact immunotherapy
C0260400|ICD9CM|HT|V07.3|Need for other prophylactic chemotherapy
C0260400|ICD9CM|PT|V07.39|Need for other prophylactic chemotherapy
C0260400|ICD9CM|AB|V07.39|Other prophylac chemothr
C0260402|ICD9CM|PT|V07.9|Unspecified prophylactic or treatment measure
C0260402|ICD9CM|AB|V07.9|Prophyl or tx meas NOS
C0260405|ICD9CM|PT|V10.00|Personal history of malignant neoplasm of gastrointestinal tract, unspecified
C0260405|ICD9CM|HT|V10.0|Personal history of malignant neoplasm of gastrointestinal tract
C0260405|ICD9CM|AB|V10.00|Hx of GI malignancy NOS
C0260406|ICD9CM|PT|V10.01|Personal history of malignant neoplasm of tongue
C0260406|ICD9CM|AB|V10.01|Hx of tongue malignancy
C0260407|ICD9CM|PT|V10.02|Personal history of malignant neoplasm of other and unspecified oral cavity and pharynx
C0260407|ICD9CM|AB|V10.02|Hx-oral/pharynx malg NEC
C0260408|ICD9CM|PT|V10.03|Personal history of malignant neoplasm of esophagus
C0260408|ICD9CM|AB|V10.03|Hx-esophageal malignancy
C0260409|ICD9CM|PT|V10.04|Personal history of malignant neoplasm of stomach
C0260409|ICD9CM|AB|V10.04|Hx of gastric malignancy
C0260410|ICD9CM|PT|V10.05|Personal history of malignant neoplasm of large intestine
C0260410|ICD9CM|AB|V10.05|Hx of colonic malignancy
C0260411|ICD9CM|PT|V10.06|Personal history of malignant neoplasm of rectum, rectosigmoid junction, and anus
C0260411|ICD9CM|AB|V10.06|Hx-rectal & anal malign
C0260412|ICD9CM|PT|V10.07|Personal history of malignant neoplasm of liver
C0260412|ICD9CM|AB|V10.07|Hx of liver malignancy
C0260413|ICD9CM|PT|V10.09|Personal history of malignant neoplasm of other gastrointestinal tract
C0260413|ICD9CM|AB|V10.09|Hx of GI malignancy NEC
C0260414|ICD9CM|HT|V10.1|Personal history of malignant neoplasm of trachea, bronchus, and lung
C0260415|ICD9CM|PT|V10.11|Personal history of malignant neoplasm of bronchus and lung
C0260415|ICD9CM|AB|V10.11|Hx-bronchogenic malignan
C0260416|ICD9CM|PT|V10.12|Personal history of malignant neoplasm of trachea
C0260416|ICD9CM|AB|V10.12|Hx-tracheal malignancy
C0260417|ICD9CM|HT|V10.2|Personal history of malignant neoplasm of other respiratory and intrathoracic organs
C0260417|ICD9CM|PT|V10.29|Personal history of malignant neoplasm of other respiratory and intrathoracic organs
C0260417|ICD9CM|AB|V10.29|Hx-intrathoracic mal NEC
C0260418|ICD9CM|PT|V10.20|Personal history of malignant neoplasm of respiratory organ, unspecified
C0260418|ICD9CM|AB|V10.20|Hx-resp org malignan NOS
C0260419|ICD9CM|PT|V10.21|Personal history of malignant neoplasm of larynx
C0260419|ICD9CM|AB|V10.21|Hx-laryngeal malignancy
C0260420|ICD9CM|PT|V10.22|Personal history of malignant neoplasm of nasal cavities, middle ear, and accessory sinuses
C0260420|ICD9CM|AB|V10.22|Hx-nose/ear/sinus malig
C0260421|ICD9CM|PT|V10.3|Personal history of malignant neoplasm of breast
C0260421|ICD9CM|AB|V10.3|Hx of breast malignancy
C0260422|ICD9CM|HT|V10.4|Personal history of malignant neoplasm of genital organs
C0260423|ICD9CM|PT|V10.40|Personal history of malignant neoplasm of female genital organ, unspecified
C0260423|ICD9CM|AB|V10.40|Hx-female genit malg NOS
C0260424|ICD9CM|PT|V10.41|Personal history of malignant neoplasm of cervix uteri
C0260424|ICD9CM|AB|V10.41|Hx-cervical malignancy
C0260425|ICD9CM|PT|V10.42|Personal history of malignant neoplasm of other parts of uterus
C0260425|ICD9CM|AB|V10.42|Hx-uterus malignancy NEC
C0260426|ICD9CM|PT|V10.43|Personal history of malignant neoplasm of ovary
C0260426|ICD9CM|AB|V10.43|Hx of ovarian malignancy
C0260427|ICD9CM|PT|V10.44|Personal history of malignant neoplasm of other female genital organs
C0260427|ICD9CM|AB|V10.44|Hx-female genit malg NEC
C0260428|ICD9CM|PT|V10.45|Personal history of malignant neoplasm of male genital organ, unspecified
C0260428|ICD9CM|AB|V10.45|Hx-male genit malig NOS
C0260429|ICD9CM|PT|V10.46|Personal history of malignant neoplasm of prostate
C0260429|ICD9CM|AB|V10.46|Hx-prostatic malignancy
C0260430|ICD9CM|PT|V10.47|Personal history of malignant neoplasm of testis
C0260430|ICD9CM|AB|V10.47|Hx-testicular malignancy
C0260431|ICD9CM|PT|V10.49|Personal history of malignant neoplasm of other male genital organs
C0260431|ICD9CM|AB|V10.49|Hx-male genit malig NEC
C0260432|ICD9CM|HT|V10.5|Personal history of malignant neoplasm of urinary organs
C0260433|ICD9CM|PT|V10.50|Personal history of malignant neoplasm of urinary organ, unspecified
C0260433|ICD9CM|AB|V10.50|Hx-urinary malignan NOS
C0260434|ICD9CM|PT|V10.51|Personal history of malignant neoplasm of bladder
C0260434|ICD9CM|AB|V10.51|Hx of bladder malignancy
C0260435|ICD9CM|PT|V10.52|Personal history of malignant neoplasm of kidney
C0260435|ICD9CM|AB|V10.52|Hx of kidney malignancy
C0260437|ICD9CM|HT|V10.6|Personal history of leukemia
C0260439|ICD9CM|PT|V10.61|Personal history of lymphoid leukemia
C0260439|ICD9CM|AB|V10.61|Hx of lymphoid leukemia
C0260440|ICD9CM|PT|V10.62|Personal history of myeloid leukemia
C0260440|ICD9CM|AB|V10.62|Hx of myeloid leukemia
C0260441|ICD9CM|PT|V10.63|Personal history of monocytic leukemia
C0260441|ICD9CM|AB|V10.63|Hx of monocytic leukemia
C0260442|ICD9CM|PT|V10.69|Personal history of other leukemia
C0260442|ICD9CM|AB|V10.69|Hx of leukemia NEC
C0260444|ICD9CM|PT|V10.71|Personal history of lymphosarcoma and reticulosarcoma
C0260444|ICD9CM|AB|V10.71|Hx-lymphosarcoma
C0260445|ICD9CM|PT|V10.72|Personal history of hodgkin's disease
C0260445|ICD9CM|AB|V10.72|Hx-hodgkin's disease
C0260446|ICD9CM|HT|V10.8|Personal history of malignant neoplasm of other sites
C0260446|ICD9CM|PT|V10.89|Personal history of malignant neoplasm of other sites
C0260446|ICD9CM|AB|V10.89|Hx of malignancy NEC
C0260447|ICD9CM|PT|V10.81|Personal history of malignant neoplasm of bone
C0260447|ICD9CM|AB|V10.81|Hx of bone malignancy
C0260448|ICD9CM|PT|V10.82|Personal history of malignant melanoma of skin
C0260448|ICD9CM|AB|V10.82|Hx-malig skin melanoma
C0260449|ICD9CM|PT|V10.83|Personal history of other malignant neoplasm of skin
C0260449|ICD9CM|AB|V10.83|Hx-skin malignancy NEC
C0260450|ICD9CM|PT|V10.84|Personal history of malignant neoplasm of eye
C0260450|ICD9CM|AB|V10.84|Hx of eye malignancy
C0260451|ICD9CM|PT|V10.85|Personal history of malignant neoplasm of brain
C0260451|ICD9CM|AB|V10.85|Hx of brain malignancy
C0260452|ICD9CM|PT|V10.86|Personal history of malignant neoplasm of other parts of nervous system
C0260452|ICD9CM|AB|V10.86|Hx-malign nerve syst NEC
C0260453|ICD9CM|PT|V10.87|Personal history of malignant neoplasm of thyroid
C0260453|ICD9CM|AB|V10.87|Hx of thyroid malignancy
C0260454|ICD9CM|PT|V10.88|Personal history of malignant neoplasm of other endocrine glands and related structures
C0260454|ICD9CM|AB|V10.88|Hx-endocrine malign NEC
C0260455|ICD9CM|PT|V10.90|Personal history of unspecified malignant neoplasm
C0260455|ICD9CM|HT|V10|Personal history of malignant neoplasm
C0260455|ICD9CM|AB|V10.90|Hx malig neoplasm NOS
C0260457|ICD9CM|PT|V11.0|Personal history of schizophrenia
C0260457|ICD9CM|AB|V11.0|Hx of schizophrenia
C0260458|ICD9CM|PT|V11.1|Personal history of affective disorders
C0260458|ICD9CM|AB|V11.1|Hx of affective disorder
C0260459|ICD9CM|PT|V11.2|Personal history of neurosis
C0260459|ICD9CM|AB|V11.2|Hx of neurosis
C0260460|ICD9CM|PT|V11.3|Personal history of alcoholism
C0260460|ICD9CM|AB|V11.3|Hx of alcoholism
C0260461|ICD9CM|PT|V11.8|Personal history of other mental disorders
C0260461|ICD9CM|AB|V11.8|Hx-mental disorder NEC
C0260462|ICD9CM|PT|V11.9|Personal history of unspecified mental disorder
C0260462|ICD9CM|HT|V11|Personal history of mental disorder
C0260462|ICD9CM|AB|V11.9|Hx-mental disorder NOS
C0260463|ICD9CM|HT|V12|Personal history of certain other diseases
C0260464|ICD9CM|HT|V12.0|Personal history of infectious and parasitic diseases
C0260465|ICD9CM|PT|V12.1|Personal history of nutritional deficiency
C0260465|ICD9CM|AB|V12.1|Hx-nutrition deficiency
C0260466|ICD9CM|HT|V12.2|Personal history of endocrine, metabolic, and immunity disorders
C0260467|ICD9CM|PT|V12.3|Personal history of diseases of blood and blood-forming organs
C0260467|ICD9CM|AB|V12.3|Hx-blood diseases
C0260469|ICD9CM|HT|V12.5|Personal history of diseases of circulatory system
C0260470|ICD9CM|HT|V12.6|Personal history of diseases of respiratory system
C0260471|ICD9CM|HT|V12.7|Personal history of diseases of digestive system
C0260472|ICD9CM|HT|V13|Personal history of other diseases
C0260473|ICD9CM|PT|V13.00|Personal history of unspecified urinary disorder
C0260473|ICD9CM|AB|V13.00|Prsnl hst urnr dsrd unsp
C0260474|ICD9CM|PT|V13.1|Personal history of trophoblastic disease
C0260474|ICD9CM|AB|V13.1|Hx-trophoblastic disease
C0260475|ICD9CM|HT|V13.2|Personal history of other genital system and obstetric disorders
C0260475|ICD9CM|PT|V13.29|Personal history of other genital system and obstetric disorders
C0260475|ICD9CM|AB|V13.29|Hx-genital/obs dis NEC
C0260476|ICD9CM|PT|V13.3|Personal history of diseases of skin and subcutaneous tissue
C0260476|ICD9CM|AB|V13.3|Hx-skin/subcutan tis dis
C0260477|ICD9CM|PT|V13.4|Personal history of arthritis
C0260477|ICD9CM|AB|V13.4|Hx of arthritis
C0260478|ICD9CM|HT|V13.5|Personal history of other musculoskeletal disorders
C0260478|ICD9CM|PT|V13.59|Personal history of other musculoskeletal disorders
C0260478|ICD9CM|AB|V13.59|Hx musculoskletl dis NEC
C0260480|ICD9CM|PT|V13.7|Personal history of perinatal problems
C0260480|ICD9CM|AB|V13.7|Hx-perinatal problems
C0260481|ICD9CM|HT|V13.8|Personal history of other specified diseases
C0260481|ICD9CM|PT|V13.89|Personal history of other specified diseases
C0260481|ICD9CM|AB|V13.89|Hx diseases NEC
C0260482|ICD9CM|PT|V13.9|Personal history of unspecified disease
C0260482|ICD9CM|AB|V13.9|Hx of disease NOS
C0260483|ICD9CM|HT|V14|Personal history of allergy to medicinal agents
C0260484|ICD9CM|PT|V14.0|Personal history of allergy to penicillin
C0260484|ICD9CM|AB|V14.0|Hx-penicillin allergy
C0260485|ICD9CM|PT|V14.1|Personal history of allergy to other antibiotic agent
C0260485|ICD9CM|AB|V14.1|Hx-antibiot allergy NEC
C0260486|ICD9CM|PT|V14.2|Personal history of allergy to sulfonamides
C0260486|ICD9CM|AB|V14.2|Hx-sulfonamides allergy
C0260487|ICD9CM|PT|V14.3|Personal history of allergy to other anti-infective agent
C0260487|ICD9CM|AB|V14.3|Hx-anti-infect allergy
C0260488|ICD9CM|PT|V14.4|Personal history of allergy to anesthetic agent
C0260488|ICD9CM|AB|V14.4|Hx-anesthetic allergy
C0260489|ICD9CM|PT|V14.5|Personal history of allergy to narcotic agent
C0260489|ICD9CM|AB|V14.5|Hx-narcotic allergy
C0260490|ICD9CM|PT|V14.6|Personal history of allergy to analgesic agent
C0260490|ICD9CM|AB|V14.6|Hx-analgesic allergy
C0260491|ICD9CM|PT|V14.7|Personal history of allergy to serum or vaccine
C0260491|ICD9CM|AB|V14.7|Hx-vaccine allergy
C0260492|ICD9CM|PT|V14.8|Personal history of allergy to other specified medicinal agents
C0260492|ICD9CM|AB|V14.8|Hx-drug allergy NEC
C0260493|ICD9CM|PT|V14.9|Personal history of allergy to unspecified medicinal agent
C0260493|ICD9CM|AB|V14.9|Hx-drug allergy NOS
C0260494|ICD9CM|HT|V15|Other personal history presenting hazards to health
C0260495|ICD9CM|PT|V15.1|Personal history of surgery to heart and great vessels, presenting hazards to health
C0260495|ICD9CM|AB|V15.1|Hx-major cardiovasc surg
C0260496|ICD9CM|PT|V15.29|Personal history of surgery to other organs
C0260496|ICD9CM|AB|V15.29|Hx surgery to organs NEC
C0260496|ICD9CM|HT|V15.2|Personal history of surgery to other organs, presenting hazards to health
C0260497|ICD9CM|PT|V15.3|Personal history of irradiation, presenting hazards to health
C0260497|ICD9CM|AB|V15.3|Hx of irradiation
C0260498|ICD9CM|HT|V15.4|Personal history of psychological trauma, presenting hazards to health
C0260499|ICD9CM|HT|V15.5|Personal history of injury, presenting hazards to health
C0260500|ICD9CM|PT|V15.6|Personal history of poisoning, presenting hazards to health
C0260500|ICD9CM|AB|V15.6|Hx of poisoning
C0260501|ICD9CM|PT|V15.7|Personal history of contraception, presenting hazards to health
C0260501|ICD9CM|AB|V15.7|Hx of contraception
C0260502|ICD9CM|HT|V15.8|Other specified personal history presenting hazards to health
C0260502|ICD9CM|PT|V15.89|Other specified personal history presenting hazards to health
C0260502|ICD9CM|AB|V15.89|Hx-health hazards NEC
C0260503|ICD9CM|PT|V15.81|Personal history of noncompliance with medical treatment, presenting hazards to health
C0260503|ICD9CM|AB|V15.81|Hx of past noncompliance
C0260504|ICD9CM|PT|V15.9|Unspecified personal history presenting hazards to health
C0260504|ICD9CM|AB|V15.9|Hx-health hazard NOS
C0260506|ICD9CM|PT|V16.0|Family history of malignant neoplasm of gastrointestinal tract
C0260506|ICD9CM|AB|V16.0|Family hx-gi malignancy
C0260507|ICD9CM|PT|V16.1|Family history of malignant neoplasm of trachea, bronchus, and lung
C0260507|ICD9CM|AB|V16.1|Fm hx-trach/bronchog mal
C0260508|ICD9CM|PT|V16.2|Family history of malignant neoplasm of other respiratory and intrathoracic organs
C0260508|ICD9CM|AB|V16.2|Fam hx-intrathoracic mal
C0260510|ICD9CM|HT|V16.4|Family history of malignant neoplasm of genital organs
C0260510|ICD9CM|PT|V16.40|Family history of malignant neoplasm of genital organ, unspecified
C0260510|ICD9CM|AB|V16.40|Fm hx genital malig NOS
C0260511|ICD9CM|HT|V16.5|Family history of malignant neoplasm of urinary organs
C0260512|ICD9CM|PT|V16.6|Family history of leukemia
C0260512|ICD9CM|AB|V16.6|Family hx-leukemia
C0260514|ICD9CM|PT|V16.8|Family history of other specified malignant neoplasm
C0260514|ICD9CM|AB|V16.8|Family hx-malignancy NEC
C0260516|ICD9CM|HT|V17|Family history of certain chronic disabling diseases
C0260517|ICD9CM|PT|V17.0|Family history of psychiatric condition
C0260517|ICD9CM|AB|V17.0|Fam hx-psychiatric cond
C0260518|ICD9CM|PT|V17.1|Family history of stroke (cerebrovascular)
C0260518|ICD9CM|AB|V17.1|Family hx-stroke
C0260519|ICD9CM|PT|V17.2|Family history of other neurological diseases
C0260519|ICD9CM|AB|V17.2|Fam hx-neurolog dis NEC
C0260520|ICD9CM|PT|V17.3|Family history of ischemic heart disease
C0260520|ICD9CM|AB|V17.3|Fam hx-ischem heart dis
C0260522|ICD9CM|PT|V17.5|Family history of asthma
C0260522|ICD9CM|AB|V17.5|Family hx-asthma
C0260523|ICD9CM|PT|V17.6|Family history of other chronic respiratory conditions
C0260523|ICD9CM|AB|V17.6|Fam hx-chr resp cond NEC
C0260524|ICD9CM|HT|V17.8|Family history of other musculoskeletal diseases
C0260524|ICD9CM|PT|V17.89|Family history of other musculoskeletal diseases
C0260524|ICD9CM|AB|V17.89|Fam hx musculosk dis NEC
C0260525|ICD9CM|HT|V18|Family history of certain other specific conditions
C0260526|ICD9CM|PT|V18.0|Family history of diabetes mellitus
C0260526|ICD9CM|AB|V18.0|Fam hx-diabetes mellitus
C0260528|ICD9CM|PT|V18.2|Family history of anemia
C0260528|ICD9CM|AB|V18.2|Family hx-anemia
C0260529|ICD9CM|PT|V18.3|Family history of other blood disorders
C0260529|ICD9CM|AB|V18.3|Fam hx-blood disord NEC
C0260530|ICD9CM|AB|V18.4|Fm hx-intellect disablty
C0260530|ICD9CM|PT|V18.4|Family history of intellectual disabilities
C0260533|ICD9CM|PT|V18.7|Family history of other genitourinary diseases
C0260533|ICD9CM|AB|V18.7|Family hx-gu disease NEC
C0260534|ICD9CM|PT|V18.8|Family history of infectious and parasitic diseases
C0260534|ICD9CM|AB|V18.8|Fm hx-infect/parasit dis
C0260535|ICD9CM|PT|V19.8|Family history of other condition
C0260535|ICD9CM|HT|V19|Family history of other conditions
C0260535|ICD9CM|AB|V19.8|Family hx-condition NEC
C0260537|ICD9CM|HT|V19.1|Family history of other eye disorders
C0260538|ICD9CM|PT|V19.2|Family history of deafness or hearing loss
C0260538|ICD9CM|AB|V19.2|Family hx-deafness
C0260539|ICD9CM|PT|V19.3|Family history of other ear disorders
C0260539|ICD9CM|AB|V19.3|Family hx-ear disord NEC
C0260540|ICD9CM|PT|V19.4|Family history of skin conditions
C0260540|ICD9CM|AB|V19.4|Family hx-skin condition
C0260541|ICD9CM|PT|V19.5|Family history of congenital anomalies
C0260541|ICD9CM|AB|V19.5|Fam hx-congen anomalies
C0260542|ICD9CM|PT|V19.6|Family history of allergic disorders
C0260542|ICD9CM|AB|V19.6|Family hx-allergic dis
C0260543|ICD9CM|HT|V20|Health supervision of infant or child
C0260545|ICD9CM|PT|V20.2|Routine infant or child health check
C0260545|ICD9CM|AB|V20.2|Routin child health exam
C0260546|ICD9CM|HT|V21|Constitutional states in development
C0260548|ICD9CM|PT|V21.8|Other specified constitutional states in development
C0260548|ICD9CM|AB|V21.8|Constit state in dev NEC
C0260549|ICD9CM|PT|V21.9|Unspecified constitutional state in development
C0260549|ICD9CM|AB|V21.9|Constit state in dev NOS
C0260550|ICD9CM|PT|V22.0|Supervision of normal first pregnancy
C0260550|ICD9CM|AB|V22.0|Supervis normal 1st preg
C0260551|ICD9CM|HT|V23|Supervision of high-risk pregnancy
C0260552|ICD9CM|PT|V23.0|Supervision of high-risk pregnancy with history of infertility
C0260552|ICD9CM|AB|V23.0|Preg w hx of infertility
C0260553|ICD9CM|PT|V23.1|Supervision of high-risk pregnancy with history of trophoblastic disease
C0260553|ICD9CM|AB|V23.1|Preg w hx-trophoblas dis
C0260554|ICD9CM|PT|V23.2|Supervision of high-risk pregnancy with history of abortion
C0260554|ICD9CM|AB|V23.2|Preg w hx of abortion
C0260555|ICD9CM|PT|V23.3|Supervision of high-risk pregnancy with grand multiparity
C0260555|ICD9CM|AB|V23.3|Grand multiparity
C0260556|ICD9CM|HT|V23.4|Supervision of high-risk pregnancy with other poor obstetric history
C0260557|ICD9CM|PT|V23.5|Supervision of high-risk pregnancy with other poor reproductive history
C0260557|ICD9CM|AB|V23.5|Preg w poor reproduct hx
C0260559|ICD9CM|HT|V23.8|Supervision of other high-risk pregnancy
C0260559|ICD9CM|PT|V23.89|Supervision of other high-risk pregnancy
C0260559|ICD9CM|AB|V23.89|Suprv high-risk preg NEC
C0260561|ICD9CM|HT|V24|Postpartum care and examination
C0260563|ICD9CM|PT|V24.1|Postpartum care and examination of lactating mother
C0260563|ICD9CM|AB|V24.1|Postpart care-lactation
C0260564|ICD9CM|PT|V24.2|Routine postpartum follow-up
C0260564|ICD9CM|AB|V24.2|Rout postpart follow-up
C0260572|ICD9CM|PT|V25.42|Surveillance of intrauterine contraceptive device
C0260572|ICD9CM|AB|V25.42|Iud surveillance
C0260574|MTH|PN|NOCODE|Contraceptive mangmt NEC in ICD9CM_2014
C0260574|ICD9CM|PT|V25.8|Other specified contraceptive management
C0260574|ICD9CM|AB|V25.8|Contraceptive mangmt NEC
C0260576|ICD9CM|PT|V26.9|Unspecified procreative management
C0260576|ICD9CM|HT|V26|Procreative management
C0260576|ICD9CM|AB|V26.9|Procreative mangmt NOS
C0260581|ICD9CM|HT|V27|Outcome of delivery
C0260587|ICD9CM|PT|V27.5|Outcome of delivery, other multiple birth, all liveborn
C0260587|ICD9CM|AB|V27.5|Del-mult birth, all live
C0260588|ICD9CM|PT|V27.6|Outcome of delivery, other multiple birth, some liveborn
C0260588|ICD9CM|AB|V27.6|Del-mult brth, some live
C0260590|ICD9CM|AB|V27.9|Outcome of delivery NOS
C0260590|ICD9CM|PT|V27.9|Outcome of delivery, unspecified outcome of delivery
C0260591|ICD9CM|AB|V28.9|Antenatal screening NOS
C0260591|ICD9CM|PT|V28.9|Unspecified antenatal screening
C0260594|ICD9CM|PT|V28.2|Other antenatal screening based on amniocentesis
C0260594|ICD9CM|AB|V28.2|Screen by amniocent NEC
C0260596|ICD9CM|PT|V28.4|Antenatal screening for fetal growth retardation using ultrasonics
C0260596|ICD9CM|AB|V28.4|Screen-fetal retardation
C0260597|ICD9CM|PT|V28.5|Antenatal screening for isoimmunization
C0260597|ICD9CM|AB|V28.5|Screen-isoimmunization
C0260598|ICD9CM|HT|V28.8|Other specified antenatal screening
C0260598|ICD9CM|PT|V28.89|Other specified antenatal screening
C0260598|ICD9CM|AB|V28.89|Antenatal screening NEC
C0260601|ICD9CM|HT|V30.0|Single liveborn, born in hospital
C0260602|ICD9CM|PT|V30.00|Single liveborn, born in hospital, delivered without mention of cesarean section
C0260602|ICD9CM|AB|V30.00|Single lb in-hosp w/o cs
C0260603|ICD9CM|PT|V30.01|Single liveborn, born in hospital, delivered by cesarean section
C0260603|ICD9CM|AB|V30.01|Single lb in-hosp w cs
C0260604|ICD9CM|PT|V30.1|Single liveborn, born before admission to hospital
C0260604|ICD9CM|AB|V30.1|Singl livebrn-before adm
C0260607|ICD9CM|HT|V31.0|Twin, mate liveborn, born in hospital
C0260608|ICD9CM|PT|V31.00|Twin birth, mate liveborn, born in hospital, delivered without mention of cesarean section
C0260608|ICD9CM|AB|V31.00|Twin-mate lb-hosp w/o cs
C0260609|ICD9CM|PT|V31.01|Twin birth, mate liveborn, born in hospital, delivered by cesarean section
C0260609|ICD9CM|AB|V31.01|Twin-mate lb-in hos w cs
C0260610|ICD9CM|PT|V31.1|Twin birth, mate liveborn, born before admission to hospital
C0260610|ICD9CM|AB|V31.1|Twin, mate lb-before adm
C0260611|ICD9CM|PT|V31.2|Twin birth, mate liveborn, born outside hospital and not hospitalized
C0260611|ICD9CM|AB|V31.2|Twin, mate lb-nonhosp
C0260612|ICD9CM|HT|V32|Twin birth, mate stillborn
C0260613|ICD9CM|HT|V32.0|Twin, mate stillborn, born in hospital
C0260614|ICD9CM|PT|V32.00|Twin birth, mate stillborn, born in hospital, delivered without mention of cesarean section
C0260614|ICD9CM|AB|V32.00|Twin-mate sb-hosp w/o cs
C0260615|ICD9CM|PT|V32.01|Twin birth, mate stillborn, born in hospital, delivered by cesarean section
C0260615|ICD9CM|AB|V32.01|Twin-mate sb-hosp w cs
C0260616|ICD9CM|PT|V32.1|Twin birth, mate stillborn, born before admission to hospital
C0260616|ICD9CM|AB|V32.1|Twin, mate sb-before adm
C0260617|ICD9CM|PT|V32.2|Twin birth, mate stillborn, born outside hospital and not hospitalized
C0260617|ICD9CM|AB|V32.2|Twin, mate sb-nonhosp
C0260619|ICD9CM|PT|V33.00|Twin birth, unspecified whether mate liveborn or stillborn, born in hospital, delivered without mention of cesarean section
C0260619|ICD9CM|AB|V33.00|Twin-NOS-in hosp w/o cs
C0260620|ICD9CM|PT|V33.01|Twin birth, unspecified whether mate liveborn or stillborn, born in hospital, delivered by cesarean section
C0260620|ICD9CM|AB|V33.01|Twin-NOS-in hosp w cs
C0260621|ICD9CM|PT|V33.1|Twin birth, unspecified whether mate liveborn or stillborn, born before admission to hospital
C0260621|ICD9CM|AB|V33.1|Twin NOS-before admissn
C0260622|ICD9CM|PT|V33.2|Twin birth, unspecified whether mate liveborn or stillborn, born outside hospital and not hospitalized
C0260622|ICD9CM|AB|V33.2|Twin NOS-nonhosp
C0260623|ICD9CM|HT|V34|Other multiple birth (three or more), mates all liveborn
C0260624|ICD9CM|HT|V34.0|Other multiple, mates all liveborn, born in hospital
C0260625|ICD9CM|PT|V34.00|Other multiple birth (three or more), mates all liveborn, born in hospital, delivered without mention of cesarean section
C0260625|ICD9CM|AB|V34.00|Oth mult lb-hosp w/o cs
C0260626|ICD9CM|PT|V34.01|Other multiple birth (three or more), mates all liveborn, born in hospital, delivered by cesarean section
C0260626|ICD9CM|AB|V34.01|Oth mult lb-in hosp w cs
C0260627|ICD9CM|PT|V34.1|Other multiple birth (three or more), mates all liveborn, born before admission to hospital
C0260627|ICD9CM|AB|V34.1|Oth mult nb-before adm
C0260628|ICD9CM|PT|V34.2|Other multiple birth (three or more), mates all liveborn, born outside hospital and not hospitalized
C0260628|ICD9CM|AB|V34.2|Oth multiple nb-nonhosp
C0260629|ICD9CM|HT|V35|Other multiple birth (three or more), mates all stillborn
C0260630|ICD9CM|HT|V35.0|Other multiple, mates all stillborn, born in hospital
C0260631|ICD9CM|PT|V35.00|Other multiple birth (three or more), mates all still born, born in hospital, delivered without mention of cesarean section
C0260631|ICD9CM|AB|V35.00|Oth mult sb-hosp w/o cs
C0260632|ICD9CM|PT|V35.01|Other multiple birth (three or more), mates all still born, born in hospital, delivered by cesarean section
C0260632|ICD9CM|AB|V35.01|Oth mult sb-in hosp w cs
C0260633|ICD9CM|PT|V35.1|Other multiple birth (three or more), mates all stillborn, born before admission to hospital
C0260633|ICD9CM|AB|V35.1|Oth mult sb-before adm
C0260634|ICD9CM|PT|V35.2|Other multiple birth (three or more), mates all stillborn, born outside of hospital and not hospitalized
C0260634|ICD9CM|AB|V35.2|Oth multiple sb-nonhosp
C0260635|ICD9CM|HT|V36|Other multiple birth (three or more), mates liveborn and stillborn
C0260636|ICD9CM|HT|V36.0|Other multiple, mates liveborn and stillborn, born in hospital
C0260637|ICD9CM|PT|V36.00|Other multiple birth (three or more), mates liveborn and stillborn, born in hospital, delivered without mention of cesarean section
C0260637|ICD9CM|AB|V36.00|Mult lb/sb-in hos w/o cs
C0260638|ICD9CM|PT|V36.01|Other multiple birth (three or more), mates liveborn and stillborn, born in hospital, delivered without mention of cesarean section
C0260638|ICD9CM|AB|V36.01|Mult lb/sb-in hosp w cs
C0260639|ICD9CM|PT|V36.1|Other multiple birth (three or more), mates liveborn and stillborn, born before admission to hospital
C0260639|ICD9CM|AB|V36.1|Mult nb/sb-before adm
C0260640|ICD9CM|PT|V36.2|Other multiple birth (three or more), mates liveborn and stillborn, born outside hospital and not hospitalized
C0260640|ICD9CM|AB|V36.2|Multiple nb/sb-nonhosp
C0260641|ICD9CM|HT|V37|Other multiple birth (three or more), unspecified whether mates liveborn or stillborn
C0260642|ICD9CM|HT|V37.0|Other multiple, unspecified, born in hospital
C0260643|ICD9CM|PT|V37.00|Other multiple birth (three or more), unspecified whether mates liveborn or stillborn, born in hospital, delivered without mention of cesarean section
C0260643|ICD9CM|AB|V37.00|Mult brth NOS-hos w/o cs
C0260644|ICD9CM|PT|V37.01|Other multiple birth (three or more), unspecified whether mates liveborn or stillborn, born in hospital, delivered by cesarean section
C0260644|ICD9CM|AB|V37.01|Mult birth NOS-hosp w cs
C0260645|ICD9CM|PT|V37.1|Other multiple birth (three or more), unspecified whether mates liveborn or stillborn, born before admission to hospital
C0260645|ICD9CM|AB|V37.1|Mult brth NOS-before adm
C0260646|ICD9CM|PT|V37.2|Other multiple birth (three or more), unspecified whether mates liveborn or stillborn, born outside of hospital
C0260646|ICD9CM|AB|V37.2|Mult birth NOS-nonhosp
C0260647|ICD9CM|HT|V39|Liveborn, unspecified whether single, twin, or multiple
C0260648|ICD9CM|HT|V39.0|Other liveborn, unspecified, born in hospital
C0260649|ICD9CM|PT|V39.00|Liveborn, unspecified whether single, twin or multiple, born in hospital, delivered without mention of cesarean section
C0260649|ICD9CM|AB|V39.00|Liveborn NOS-hosp w/o cs
C0260650|ICD9CM|PT|V39.01|Liveborn, unspecified whether single, twin or multiple, born in hospital, delivered by cesarean section
C0260650|ICD9CM|AB|V39.01|Liveborn NOS-hosp w cs
C0260651|ICD9CM|PT|V39.1|Liveborn, unspecified whether single, twin or multiple, born before admission to hospital
C0260651|ICD9CM|AB|V39.1|Liveborn NOS-before adm
C0260652|ICD9CM|PT|V39.2|Liveborn, unspecified whether single, twin or multiple, born outside hospital and not hospitalized
C0260652|ICD9CM|AB|V39.2|Liveborn NOS-nonhosp
C0260654|MTH|PN|NOCODE|Mental and behavioral problems with learning in ICD9CM
C0260654|ICD9CM|PT|V40.0|Mental and behavioral problems with learning
C0260654|ICD9CM|AB|V40.0|Problems with learning
C0260655|ICD9CM|PT|V40.1|Mental and behavioral problems with communication [including speech]
C0260655|ICD9CM|AB|V40.1|Prob with communication
C0260656|ICD9CM|PT|V40.2|Other mental problems
C0260656|ICD9CM|AB|V40.2|Mental problems NEC
C0260657|ICD9CM|HT|V40.3|Other behavioral problems
C0260658|ICD9CM|PT|V40.9|Unspecified mental or behavioral problem
C0260658|ICD9CM|HT|V40|Mental and behavioral problems
C0260658|ICD9CM|AB|V40.9|Mental/behavior prob NOS
C0260659|ICD9CM|HT|V41|Problems with special senses and other special functions
C0260661|ICD9CM|PT|V41.1|Other eye problems
C0260661|ICD9CM|AB|V41.1|Eye problems NEC
C0260663|ICD9CM|PT|V41.3|Other ear problems
C0260663|ICD9CM|AB|V41.3|Ear problems NEC
C0260664|ICD9CM|AB|V41.4|Voice production problem
C0260664|ICD9CM|PT|V41.4|Problems with voice production
C0260665|ICD9CM|PT|V41.5|Problems with smell and taste
C0260665|ICD9CM|AB|V41.5|Smell and taste problem
C0260667|ICD9CM|AB|V41.7|Sexual function problem
C0260667|ICD9CM|PT|V41.7|Problems with sexual function
C0260668|ICD9CM|PT|V41.8|Other problems with special functions
C0260668|ICD9CM|AB|V41.8|Probl w special func NEC
C0260669|ICD9CM|PT|V41.9|Unspecified problem with special functions
C0260669|ICD9CM|AB|V41.9|Probl w special func NOS
C0260672|ICD9CM|HT|V43|Organ or tissue replaced by other means
C0260673|ICD9CM|PT|V43.0|Eye globe replaced by other means
C0260673|ICD9CM|AB|V43.0|Eye replacement NEC
C0260674|ICD9CM|HT|V43.2|Heart replaced by other means
C0260675|ICD9CM|PT|V43.3|Heart valve replaced by other means
C0260675|ICD9CM|AB|V43.3|Heart valve replac NEC
C0260676|ICD9CM|PT|V43.4|Blood vessel replaced by other means
C0260676|ICD9CM|AB|V43.4|Blood vessel replac NEC
C0260678|ICD9CM|HT|V43.6|Joint replaced by other means
C0260679|ICD9CM|PT|V43.7|Limb replaced by other means
C0260679|ICD9CM|AB|V43.7|Limb replacement NEC
C0260680|ICD9CM|HT|V43.8|Other organ or tissue replaced by other means
C0260680|ICD9CM|PT|V43.89|Other organ or tissue replaced by other means
C0260680|ICD9CM|AB|V43.89|Organ/tiss replacmnt NEC
C0260682|ICD9CM|AB|V44.0|Tracheostomy status
C0260682|ICD9CM|PT|V44.0|Tracheostomy status
C0260683|ICD9CM|AB|V44.1|Gastrostomy status
C0260683|ICD9CM|PT|V44.1|Gastrostomy status
C0260684|ICD9CM|AB|V44.2|Ileostomy status
C0260684|ICD9CM|PT|V44.2|Ileostomy status
C0260685|ICD9CM|AB|V44.3|Colostomy status
C0260685|ICD9CM|PT|V44.3|Colostomy status
C0260686|ICD9CM|PT|V44.4|Status of other artificial opening of gastrointestinal tract
C0260686|ICD9CM|AB|V44.4|Enterostomy status NEC
C0260687|ICD9CM|HT|V44.5|Cystostomy status
C0260687|ICD9CM|AB|V44.50|Cystostomy status NOS
C0260687|ICD9CM|PT|V44.50|Cystostomy, unspecified
C0260688|ICD9CM|PT|V44.6|Other artificial opening of urinary tract status
C0260688|ICD9CM|AB|V44.6|Urinostomy status NEC
C0260689|ICD9CM|AB|V44.7|Artificial vagina status
C0260689|ICD9CM|PT|V44.7|Artificial vagina status
C0260690|ICD9CM|PT|V44.8|Other artificial opening status
C0260690|ICD9CM|AB|V44.8|Artif open status NEC
C0260691|ICD9CM|HT|V44|Artificial opening status
C0260691|ICD9CM|PT|V44.9|Unspecified artificial opening status
C0260691|ICD9CM|AB|V44.9|Artif open status NOS
C0260694|ICD9CM|HT|V45.1|Postsurgical renal dialysis status
C0260698|ICD9CM|HT|V45.8|Other postprocedural status
C0260698|ICD9CM|PT|V45.89|Other postprocedural status
C0260698|ICD9CM|HT|V45|Other postprocedural states
C0260698|ICD9CM|AB|V45.89|Post-proc states NEC
C0260700|ICD9CM|AB|V46.0|Dependence on aspirator
C0260700|ICD9CM|PT|V46.0|Dependence on aspirator
C0260702|ICD9CM|PT|V46.8|Dependence on other enabling machines
C0260702|ICD9CM|AB|V46.8|Machine dependence NEC
C0260703|ICD9CM|AB|V46.9|Machine dependence NOS
C0260703|ICD9CM|PT|V46.9|Unspecified machine dependence
C0260704|ICD9CM|HT|V47|Other problems with internal organs
C0260705|ICD9CM|PT|V47.0|Deficiencies of internal organs
C0260705|ICD9CM|AB|V47.0|Intern organ deficiency
C0260706|ICD9CM|PT|V47.1|Mechanical and motor problems with internal organs
C0260706|ICD9CM|AB|V47.1|Mech prob w internal org
C0260707|ICD9CM|PT|V47.2|Other cardiorespiratory problems
C0260707|ICD9CM|AB|V47.2|Cardiorespirat probl NEC
C0260708|ICD9CM|PT|V47.3|Other digestive problems
C0260708|ICD9CM|AB|V47.3|Digestive problems NEC
C0260709|ICD9CM|PT|V47.4|Other urinary problems
C0260709|ICD9CM|AB|V47.4|Urinary problems NEC
C0260710|ICD9CM|PT|V47.5|Other genital problems
C0260710|ICD9CM|AB|V47.5|Genital problems NEC
C0260711|ICD9CM|PT|V47.9|Unspecified problems with internal organs
C0260711|ICD9CM|AB|V47.9|Probl w internal org NOS
C0260712|ICD9CM|HT|V48|Problems with head, neck, and trunk
C0260713|ICD9CM|AB|V48.0|Deficiencies of head
C0260713|ICD9CM|PT|V48.0|Deficiencies of head
C0260714|ICD9CM|PT|V48.1|Deficiencies of neck and trunk
C0260714|ICD9CM|AB|V48.1|Deficiencies neck/trunk
C0260715|ICD9CM|PT|V48.2|Mechanical and motor problems with head
C0260715|ICD9CM|AB|V48.2|Mechanical prob w head
C0260716|ICD9CM|PT|V48.3|Mechanical and motor problems with neck and trunk
C0260716|ICD9CM|AB|V48.3|Mech prob w neck & trunk
C0260717|ICD9CM|PT|V48.4|Sensory problem with head
C0260717|ICD9CM|AB|V48.4|Sensory problem w head
C0260718|ICD9CM|PT|V48.5|Sensory problem with neck and trunk
C0260718|ICD9CM|AB|V48.5|Sensor prob w neck/trunk
C0260719|ICD9CM|AB|V48.6|Disfigurements of head
C0260719|ICD9CM|PT|V48.6|Disfigurements of head
C0260720|ICD9CM|PT|V48.7|Disfigurements of neck and trunk
C0260720|ICD9CM|AB|V48.7|Disfigurement neck/trunk
C0260721|ICD9CM|PT|V48.8|Other problems with head, neck, and trunk
C0260721|ICD9CM|AB|V48.8|Prob-head/neck/trunk NEC
C0260722|ICD9CM|PT|V48.9|Unspecified problem with head, neck, or trunk
C0260722|ICD9CM|AB|V48.9|Prob-head/neck/trunk NOS
C0260724|ICD9CM|AB|V49.0|Deficiencies of limbs
C0260724|ICD9CM|PT|V49.0|Deficiencies of limbs
C0260725|ICD9CM|PT|V49.1|Mechanical problems with limbs
C0260725|ICD9CM|AB|V49.1|Mechanical prob w limbs
C0260726|ICD9CM|PT|V49.2|Motor problems with limbs
C0260726|ICD9CM|AB|V49.2|Motor problems w limbs
C0260727|ICD9CM|PT|V49.3|Sensory problems with limbs
C0260727|ICD9CM|AB|V49.3|Sensory problems w limbs
C0260728|ICD9CM|AB|V49.4|Disfigurements of limbs
C0260728|ICD9CM|PT|V49.4|Disfigurements of limbs
C0260729|ICD9CM|PT|V49.9|Unspecified problems with limbs and other problems
C0260729|ICD9CM|AB|V49.9|Probl influ health NOS
C0260731|ICD9CM|HT|V50|Elective surgery for purposes other than remedying health states
C0260734|ICD9CM|PT|V50.8|Other elective surgery for purposes other than remedying health states
C0260734|ICD9CM|AB|V50.8|Elective surgery NEC
C0260735|ICD9CM|PT|V50.9|Unspecified elective surgery for purposes other than remedying health states
C0260735|ICD9CM|AB|V50.9|Elective surgery NOS
C0260736|ICD9CM|HT|V51|Aftercare involving the use of plastic surgery
C0260738|ICD9CM|PT|V52.0|Fitting and adjustment of artificial arm (complete) (partial)
C0260738|ICD9CM|AB|V52.0|Fitting artificial arm
C0260739|ICD9CM|PT|V52.1|Fitting and adjustment of artificial leg (complete) (partial)
C0260739|ICD9CM|AB|V52.1|Fitting artificial leg
C0260743|ICD9CM|PT|V52.8|Fitting and adjustment of other specified prosthetic device
C0260743|ICD9CM|AB|V52.8|Fitting prosthesis NEC
C0260744|ICD9CM|PT|V52.9|Fitting and adjustment of unspecified prosthetic device
C0260744|ICD9CM|AB|V52.9|Fitting prosthesis NOS
C0260745|ICD9CM|PT|V53.99|Fitting and adjustment, other device
C0260745|ICD9CM|HT|V53|Fitting and adjustment of other device
C0260745|ICD9CM|AB|V53.99|Fit/adjust device NEC
C0260746|ICD9CM|HT|V53.0|Fitting and adjustment of devices related to nervous system and special senses
C0260747|ICD9CM|PT|V53.1|Fitting and adjustment of spectacles and contact lenses
C0260747|ICD9CM|AB|V53.1|Fit contact lens/glasses
C0260748|ICD9CM|PT|V53.2|Fitting and adjustment of hearing aid
C0260748|ICD9CM|AB|V53.2|Adjustment hearing aid
C0260749|ICD9CM|HT|V53.3|Fitting and adjustment of cardiac pacemaker
C0260749|ICD9CM|PT|V53.31|Fitting and adjustment of cardiac pacemaker
C0260749|ICD9CM|AB|V53.31|Ftng cardiac pacemaker
C0260750|ICD9CM|PT|V53.4|Fitting and adjustment of orthodontic devices
C0260750|ICD9CM|AB|V53.4|Fit orthodontic device
C0260752|ICD9CM|PT|V53.6|Fitting and adjustment of urinary devices
C0260752|ICD9CM|AB|V53.6|Fitting urinary devices
C0260753|ICD9CM|PT|V53.7|Fitting and adjustment of orthopedic devices
C0260753|ICD9CM|AB|V53.7|Fit orthopedic devices
C0260755|ICD9CM|HT|V53.9|Fitting and adjustment of other and unspecified device
C0260756|ICD9CM|HT|V54|Other orthopedic aftercare
C0260756|ICD9CM|HT|V54.8|Other orthopedic aftercare
C0260756|ICD9CM|PT|V54.89|Other orthopedic aftercare
C0260756|ICD9CM|AB|V54.89|Orthopedic aftercare NEC
C0260757|ICD9CM|HT|V54.0|Aftercare involving internal fixation device
C0260758|ICD9CM|PT|V54.9|Unspecified orthopedic aftercare
C0260758|ICD9CM|AB|V54.9|Orthopedic aftercare NOS
C0260760|ICD9CM|PT|V55.0|Attention to tracheostomy
C0260760|ICD9CM|AB|V55.0|Atten to tracheostomy
C0260761|ICD9CM|PT|V55.1|Attention to gastrostomy
C0260761|ICD9CM|AB|V55.1|Atten to gastrostomy
C0260762|ICD9CM|PT|V55.2|Attention to ileostomy
C0260762|ICD9CM|AB|V55.2|Atten to ileostomy
C0260763|ICD9CM|PT|V55.3|Attention to colostomy
C0260763|ICD9CM|AB|V55.3|Atten to colostomy
C0260764|ICD9CM|PT|V55.4|Attention to other artificial opening of digestive tract
C0260764|ICD9CM|AB|V55.4|Atten to enterostomy NEC
C0260765|ICD9CM|PT|V55.5|Attention to cystostomy
C0260765|ICD9CM|AB|V55.5|Atten to cystostomy
C0260766|ICD9CM|PT|V55.6|Attention to other artificial opening of urinary tract
C0260766|ICD9CM|AB|V55.6|Atten to urinostomy NEC
C0260767|ICD9CM|PT|V55.7|Attention to artificial vagina
C0260767|ICD9CM|AB|V55.7|Atten artificial vagina
C0260768|ICD9CM|PT|V55.8|Attention to other specified artificial opening
C0260768|ICD9CM|AB|V55.8|Attn to artif open NEC
C0260771|ICD9CM|PT|V56.0|Encounter for extracorporeal dialysis
C0260771|ICD9CM|AB|V56.0|Renal dialysis encounter
C0260774|ICD9CM|PT|V57.4|Care involving orthoptic training
C0260774|ICD9CM|AB|V57.4|Orthoptic training
C0260775|ICD9CM|HT|V57.8|Care involving other specified rehabilitation procedure
C0260775|ICD9CM|PT|V57.89|Care involving other specified rehabilitation procedure
C0260775|ICD9CM|AB|V57.89|Rehabilitation proc NEC
C0260776|ICD9CM|PT|V57.81|Care involving orthotic training
C0260776|ICD9CM|AB|V57.81|Orthotic training
C0260777|ICD9CM|HT|V58|Encounter for other and unspecified procedures and aftercare
C0260778|ICD9CM|PT|V58.0|Encounter for radiotherapy
C0260778|ICD9CM|AB|V58.0|Radiotherapy encounter
C0260780|ICD9CM|PT|V58.2|Blood transfusion, without reported diagnosis
C0260780|ICD9CM|AB|V58.2|Blood transfusion, no dx
C0260782|ICD9CM|HT|V58.4|Other aftercare following surgery
C0260783|ICD9CM|PT|V58.89|Other specified aftercare
C0260783|ICD9CM|AB|V58.89|Other specfied aftercare
C0260784|ICD9CM|PT|V58.9|Unspecified aftercare
C0260784|ICD9CM|AB|V58.9|Aftercare NOS
C0260785|ICD9CM|AB|V59.1|Skin donor
C0260785|ICD9CM|PT|V59.1|Skin donors
C0260789|ICD9CM|AB|V59.5|Cornea donor
C0260789|ICD9CM|PT|V59.5|Cornea donors
C0260790|ICD9CM|PT|V59.8|Donors of other specified organ or tissue
C0260790|ICD9CM|AB|V59.8|Org or tissue donor NEC
C0260791|ICD9CM|HT|V60|Housing, household, and economic circumstances
C0260793|ICD9CM|AB|V60.1|Inadequate housing
C0260793|ICD9CM|PT|V60.1|Inadequate housing
C0260794|ICD9CM|AB|V60.3|Person living alone
C0260794|ICD9CM|PT|V60.3|Person living alone
C0260795|ICD9CM|PT|V60.4|No other household member able to render care
C0260795|ICD9CM|AB|V60.4|No family able to care
C0260796|ICD9CM|AB|V60.5|Holiday relief care
C0260796|ICD9CM|PT|V60.5|Holiday relief care
C0260797|ICD9CM|PT|V60.6|Person living in residential institution
C0260797|ICD9CM|AB|V60.6|Person in resident inst
C0260798|ICD9CM|HT|V60.8|Other specified housing or economic circumstances
C0260799|ICD9CM|PT|V60.9|Unspecified housing or economic circumstance
C0260799|ICD9CM|AB|V60.9|Housing/econo circum NOS
C0260801|ICD9CM|PT|V61.3|Problems with aged parents or in-laws
C0260801|ICD9CM|AB|V61.3|Problem w aged parent
C0260804|ICD9CM|PT|V61.49|Other health problems within the family
C0260804|ICD9CM|AB|V61.49|Family health probl NEC
C0260805|ICD9CM|HT|V62|Other psychosocial circumstances
C0260806|ICD9CM|PT|V62.1|Adverse effects of work environment
C0260806|ICD9CM|AB|V62.1|Adverse eff-work environ
C0260807|ICD9CM|AB|V62.5|Legal circumstances
C0260807|ICD9CM|PT|V62.5|Legal circumstances
C0260808|ICD9CM|PT|V62.9|Unspecified psychosocial circumstance
C0260808|ICD9CM|AB|V62.9|Psychosocial circum NOS
C0260809|ICD9CM|HT|V63|Unavailability of other medical facilities for care
C0260810|ICD9CM|PT|V63.0|Residence remote from hospital or other health care facility
C0260810|ICD9CM|AB|V63.0|Home remote from hospitl
C0260812|ICD9CM|PT|V63.2|Person awaiting admission to adequate facility elsewhere
C0260812|ICD9CM|AB|V63.2|Wait adm to oth facility
C0260813|ICD9CM|PT|V63.8|Other specified reasons for unavailability of medical facilities
C0260813|ICD9CM|AB|V63.8|No med facilities NEC
C0260814|ICD9CM|PT|V63.9|Unspecified reason for unavailability of medical facilities
C0260814|ICD9CM|AB|V63.9|No med facilities NOS
C0260815|ICD9CM|HT|V64|Persons encountering health services for specific procedures, not carried out
C0260817|ICD9CM|PT|V64.1|Surgical or other procedure not carried out because of contraindication
C0260817|ICD9CM|AB|V64.1|No proc/contraindication
C0260818|ICD9CM|PT|V64.2|Surgical or other procedure not carried out because of patient's decision
C0260818|ICD9CM|AB|V64.2|No proc/patient decision
C0260819|ICD9CM|PT|V64.3|Procedure not carried out for other reasons
C0260819|ICD9CM|AB|V64.3|No proc for reasons NEC
C0260820|ICD9CM|HT|V65|Other persons seeking consultation
C0260821|ICD9CM|PT|V65.0|Healthy person accompanying sick person
C0260821|ICD9CM|AB|V65.0|Healthy person w sick
C0260822|ICD9CM|HT|V65.1|Person consulting on behalf of another person
C0260823|ICD9CM|PT|V65.3|Dietary surveillance and counseling
C0260823|ICD9CM|AB|V65.3|Dietary surveil/counsel
C0260825|ICD9CM|PT|V65.8|Other reasons for seeking consultation
C0260825|ICD9CM|AB|V65.8|Reason for consult NEC
C0260826|ICD9CM|PT|V66.0|Convalescence following surgery
C0260826|ICD9CM|AB|V66.0|Surgical convalescence
C0260827|ICD9CM|PT|V66.1|Convalescence following radiotherapy
C0260827|ICD9CM|AB|V66.1|Radiotherapy convalescen
C0260828|ICD9CM|PT|V66.2|Convalescence following chemotherapy
C0260828|ICD9CM|AB|V66.2|Chemotherapy convalescen
C0260830|ICD9CM|PT|V66.4|Convalescence following treatment of fracture
C0260830|ICD9CM|AB|V66.4|Fracture treatmnt conval
C0260832|ICD9CM|HT|V67|Follow-up examination
C0260832|ICD9CM|PT|V67.9|Unspecified follow-up examination
C0260832|ICD9CM|AB|V67.9|Follow-up exam NOS
C0260833|ICD9CM|HT|V67.0|Follow-up examination following surgery
C0260834|ICD9CM|AB|V67.1|Radiotherapy follow-up
C0260834|ICD9CM|PT|V67.1|Follow-up examination, following radiotherapy
C0260836|ICD9CM|AB|V67.3|Psychiatric follow-up
C0260836|ICD9CM|PT|V67.3|Follow-up examination, following psychotherapy and other treatment for mental disorder
C0260838|ICD9CM|HT|V67.5|Follow-up examination following other treatment
C0260840|ICD9CM|PT|V67.59|Other follow-up examination
C0260840|ICD9CM|AB|V67.59|Follow-up exam NEC
C0260841|ICD9CM|PT|V67.6|Follow-up examination, following combined treatment
C0260841|ICD9CM|AB|V67.6|Comb treatment follow-up
C0260843|ICD9CM|HT|V68|Encounters for administrative purposes
C0260844|ICD9CM|HT|V68.0|Issue of medical certificates
C0260845|ICD9CM|PT|V68.1|Issue of repeat prescriptions
C0260845|ICD9CM|AB|V68.1|Issue repeat prescript
C0260846|ICD9CM|PT|V68.2|Request for expert evidence
C0260846|ICD9CM|AB|V68.2|Request expert evidence
C0260847|ICD9CM|HT|V68.8|Encounters for other specified administrative purpose
C0260847|ICD9CM|PT|V68.89|Encounters for other specified administrative purpose
C0260847|ICD9CM|AB|V68.89|Administrtve encount NEC
C0260848|ICD9CM|PT|V68.81|Referral of patient without examination or treatment
C0260848|ICD9CM|AB|V68.81|Referral-no exam/treat
C0260849|ICD9CM|PT|V68.9|Encounters for unspecified administrative purpose
C0260849|ICD9CM|AB|V68.9|Administrtve encount NOS
C0260851|ICD9CM|PT|V70.0|Routine general medical examination at a health care facility
C0260851|ICD9CM|AB|V70.0|Routine medical exam
C0260852|ICD9CM|PT|V70.1|General psychiatric examination, requested by the authority
C0260852|ICD9CM|AB|V70.1|Psych exam-authority req
C0260855|ICD9CM|PT|V70.4|Examination for medicolegal reasons
C0260855|ICD9CM|AB|V70.4|Exam-medicolegal reasons
C0260856|ICD9CM|PT|V70.5|Health examination of defined subpopulations
C0260856|ICD9CM|AB|V70.5|Health exam-group survey
C0260857|ICD9CM|PT|V70.6|Health examination in population surveys
C0260857|ICD9CM|AB|V70.6|Health exam-pop survey
C0260859|ICD9CM|PT|V70.8|Other specified general medical examinations
C0260859|ICD9CM|AB|V70.8|General medical exam NEC
C0260860|ICD9CM|HT|V70|General medical examination
C0260860|ICD9CM|PT|V70.9|Unspecified general medical examination
C0260860|ICD9CM|AB|V70.9|General medical exam NOS
C0260862|ICD9CM|HT|V71.0|Observation for suspected mental condition
C0260863|ICD9CM|PT|V71.01|Observation for adult antisocial behavior
C0260863|ICD9CM|AB|V71.01|Obsv-adult antisoc behav
C0260864|ICD9CM|PT|V71.02|Observation for childhood or adolescent antisocial behavior
C0260864|ICD9CM|AB|V71.02|Obsv-adolesc antisoc beh
C0260865|ICD9CM|PT|V71.09|Observation for other suspected mental condition
C0260865|ICD9CM|AB|V71.09|Observ-mental cond NEC
C0260866|ICD9CM|PT|V71.1|Observation for suspected malignant neoplasm
C0260866|ICD9CM|AB|V71.1|Obsv-suspct mal neoplasm
C0260867|ICD9CM|PT|V71.2|Observation for suspected tuberculosis
C0260867|ICD9CM|AB|V71.2|Observ-suspect TB
C0260868|ICD9CM|PT|V71.3|Observation following accident at work
C0260868|ICD9CM|AB|V71.3|Observ-work accident
C0260869|ICD9CM|PT|V71.4|Observation following other accident
C0260869|ICD9CM|AB|V71.4|Observ-accident NEC
C0260870|ICD9CM|PT|V71.5|Observation following alleged rape or seduction
C0260870|ICD9CM|AB|V71.5|Observ following rape
C0260871|ICD9CM|PT|V71.6|Observation following other inflicted injury
C0260871|ICD9CM|AB|V71.6|Observ-inflicted inj NEC
C0260872|ICD9CM|PT|V71.7|Observation for suspected cardiovascular disease
C0260872|ICD9CM|AB|V71.7|Obs-susp cardiovasc dis
C0260875|ICD9CM|HT|V72|Special investigations and examinations
C0260876|ICD9CM|PT|V72.40|Pregnancy examination or test, pregnancy unconfirmed
C0260876|ICD9CM|AB|V72.40|Pregnancy test unconfirm
C0260877|ICD9CM|HT|V72.6|Laboratory examination
C0260879|ICD9CM|PT|V72.85|Other specified examination
C0260879|ICD9CM|HT|V72.8|Other specified examinations
C0260879|ICD9CM|AB|V72.85|Oth specified exam
C0260880|ICD9CM|PT|V72.9|Unspecified examination
C0260880|ICD9CM|AB|V72.9|Examination NOS
C0260882|ICD9CM|PT|V73.0|Screening examination for poliomyelitis
C0260882|ICD9CM|AB|V73.0|Screening-poliomyelitis
C0260883|MTH|PN|NOCODE|Screening examination for smallpox in ICD9CM
C0260883|ICD9CM|PT|V73.1|Screening examination for smallpox
C0260883|ICD9CM|AB|V73.1|Screening for smallpox
C0260884|MTH|PN|NOCODE|Screening examination for measles in ICD9CM
C0260884|ICD9CM|PT|V73.2|Screening examination for measles
C0260884|ICD9CM|AB|V73.2|Screening for measles
C0260887|ICD9CM|PT|V73.5|Screening examination for other arthropod-borne viral diseases
C0260887|ICD9CM|AB|V73.5|Screening-arbovirus dis
C0260889|ICD9CM|PT|V73.89|Special screening examination for other specified viral diseases
C0260889|ICD9CM|AB|V73.89|Scrn oth spcf viral dis
C0260892|MTH|PN|NOCODE|Screening examination for cholera in ICD9CM
C0260892|ICD9CM|PT|V74.0|Screening examination for cholera
C0260892|ICD9CM|AB|V74.0|Screening for cholera
C0260894|MTH|PN|NOCODE|Screening examination for diphtheria in ICD9CM
C0260894|ICD9CM|PT|V74.3|Screening examination for diphtheria
C0260894|ICD9CM|AB|V74.3|Screening for diphtheria
C0260895|ICD9CM|PT|V74.4|Screening examination for bacterial conjunctivitis
C0260895|ICD9CM|AB|V74.4|Screen-bact conjunctivit
C0260897|ICD9CM|AB|V74.6|Screening for yaws
C0260897|ICD9CM|PT|V74.6|Screening examination for yaws
C0260898|ICD9CM|PT|V74.8|Screening examination for other specified bacterial and spirochetal diseases
C0260898|ICD9CM|AB|V74.8|Screen-bacterial dis NEC
C0260899|ICD9CM|HT|V74|Special screening examination for bacterial and spirochetal diseases
C0260899|ICD9CM|PT|V74.9|Screening examination for unspecified bacterial and spirochetal diseases
C0260899|ICD9CM|AB|V74.9|Screen-bacterial dis NOS
C0260900|ICD9CM|HT|V75|Special screening examination for other infectious diseases
C0260901|ICD9CM|PT|V75.0|Screening examination for rickettsial diseases
C0260901|ICD9CM|AB|V75.0|Screen-rickettsial dis
C0260902|MTH|PN|NOCODE|Screening examination for malaria in ICD9CM
C0260902|ICD9CM|PT|V75.1|Screening examination for malaria
C0260902|ICD9CM|AB|V75.1|Screening for malaria
C0260905|ICD9CM|PT|V75.4|Screening examination for mycotic infections
C0260905|ICD9CM|AB|V75.4|Screen-mycotic infect
C0260906|ICD9CM|PT|V75.5|Screening examination for schistosomiasis
C0260906|ICD9CM|AB|V75.5|Screen-schistosomiasis
C0260907|ICD9CM|PT|V75.6|Screening examination for filariasis
C0260907|ICD9CM|AB|V75.6|Screen for filariasis
C0260909|ICD9CM|PT|V75.8|Screening examination for other specified parasitic infections
C0260909|ICD9CM|AB|V75.8|Screen-parasitic dis NEC
C0260910|ICD9CM|PT|V75.9|Screening examination for unspecified infectious disease
C0260910|ICD9CM|AB|V75.9|Screen for infec dis NOS
C0260914|ICD9CM|PT|V76.2|Screening for malignant neoplasms of cervix
C0260914|ICD9CM|AB|V76.2|Screen mal neop-cervix
C0260915|ICD9CM|PT|V76.3|Screening for malignant neoplasms of bladder
C0260915|ICD9CM|AB|V76.3|Screen mal neop-bladder
C0260917|ICD9CM|PT|V76.41|Screening for malignant neoplasms of rectum
C0260917|ICD9CM|AB|V76.41|Screen mal neop-rectum
C0260918|ICD9CM|PT|V76.42|Screening for malignant neoplasms of oral cavity
C0260918|ICD9CM|AB|V76.42|Screen mal neop-oral cav
C0260919|ICD9CM|PT|V76.43|Screening for malignant neoplasms of skin
C0260919|ICD9CM|AB|V76.43|Screen mal neop-skin
C0260922|ICD9CM|HT|V76|Special screening for malignant neoplasms
C0260922|ICD9CM|AB|V76.9|Screen-neoplasm NOS
C0260922|ICD9CM|PT|V76.9|Special screening for unspecified malignant neoplasms
C0260923|ICD9CM|HT|V77|Special screening for endocrine, nutritional, metabolic, and immunity disorders
C0260924|ICD9CM|PT|V77.0|Screening for thyroid disorders
C0260924|ICD9CM|AB|V77.0|Screen-thyroid disorder
C0260925|ICD9CM|PT|V77.1|Screening for diabetes mellitus
C0260925|ICD9CM|AB|V77.1|Screen-diabetes mellitus
C0260926|ICD9CM|PT|V77.2|Screening for malnutrition
C0260926|ICD9CM|AB|V77.2|Screen for malnutrition
C0260927|ICD9CM|PT|V77.3|Screening for phenylketonuria (PKU)
C0260927|ICD9CM|AB|V77.3|Screen-phenylketonuria
C0260928|ICD9CM|PT|V77.4|Screening for galactosemia
C0260928|ICD9CM|AB|V77.4|Screen for galactosemia
C0260929|ICD9CM|AB|V77.5|Screening for gout
C0260929|ICD9CM|PT|V77.5|Screening for gout
C0260930|ICD9CM|PT|V77.6|Screening for cystic fibrosis
C0260930|ICD9CM|AB|V77.6|Screen-cystic fibrosis
C0260931|ICD9CM|PT|V77.7|Screening for other inborn errors of metabolism
C0260931|ICD9CM|AB|V77.7|Screen-inborn err metab
C0260932|ICD9CM|AB|V77.8|Screening for obesity
C0260932|ICD9CM|PT|V77.8|Screening for obesity
C0260934|ICD9CM|HT|V78|Special screening for disorders of blood and blood-forming organs
C0260935|ICD9CM|PT|V78.0|Screening for iron deficiency anemia
C0260935|ICD9CM|AB|V78.0|Screen-iron defic anemia
C0260936|ICD9CM|PT|V78.1|Screening for other and unspecified deficiency anemia
C0260936|ICD9CM|AB|V78.1|Screen-defic anemia NEC
C0260937|ICD9CM|PT|V78.2|Screening for sickle-cell disease or trait
C0260937|ICD9CM|AB|V78.2|Screen-sickle cell dis
C0260939|ICD9CM|PT|V78.8|Screening for other disorders of blood and blood-forming organs
C0260939|ICD9CM|AB|V78.8|Screen-blood dis NEC
C0260940|ICD9CM|PT|V78.9|Screening for unspecified disorder of blood and blood-forming organs
C0260940|ICD9CM|AB|V78.9|Screen-blood dis NOS
C0260941|ICD9CM|HT|V79|Special screening for mental disorders and developmental handicaps
C0260942|ICD9CM|AB|V79.0|Screening for depression
C0260942|ICD9CM|PT|V79.0|Screening for depression
C0260943|ICD9CM|AB|V79.1|Screening for alcoholism
C0260943|ICD9CM|PT|V79.1|Screening for alcoholism
C0260944|ICD9CM|PT|V79.2|Special screening for intellectual disabilities
C0260944|ICD9CM|AB|V79.2|Scrn intellect disabilty
C0260945|ICD9CM|PT|V79.3|Screening for developmental handicaps in early childhood
C0260945|ICD9CM|AB|V79.3|Screen-development prob
C0260946|ICD9CM|PT|V79.8|Screening for other specified mental disorders and developmental handicaps
C0260946|ICD9CM|AB|V79.8|Screen-mental dis NEC
C0260948|ICD9CM|HT|V80|Special screening for neurological, eye, and ear diseases
C0260949|ICD9CM|HT|V80.0|Screening for neurological conditions
C0260950|ICD9CM|AB|V80.1|Screening for glaucoma
C0260950|ICD9CM|PT|V80.1|Screening for glaucoma
C0260951|ICD9CM|PT|V80.2|Screening for other eye conditions
C0260951|ICD9CM|AB|V80.2|Screening-eye cond NEC
C0260952|ICD9CM|PT|V80.3|Screening for ear diseases
C0260952|ICD9CM|AB|V80.3|Screening for ear dis
C0260953|ICD9CM|HT|V81|Special screening for cardiovascular, respiratory, and genitourinary diseases
C0260954|ICD9CM|PT|V81.0|Screening for ischemic heart disease
C0260954|ICD9CM|AB|V81.0|Scrn-ischemic heart dis
C0260955|ICD9CM|PT|V81.1|Screening for hypertension
C0260955|ICD9CM|AB|V81.1|Screen for hypertension
C0260956|ICD9CM|PT|V81.2|Screening for other and unspecified cardiovascular conditions
C0260956|ICD9CM|AB|V81.2|Screen-cardiovasc NEC
C0260957|ICD9CM|PT|V81.3|Screening for chronic bronchitis and emphysema
C0260957|ICD9CM|AB|V81.3|Screen-bronch/emphysema
C0260958|ICD9CM|PT|V81.4|Screening for other and unspecified respiratory conditions
C0260958|ICD9CM|AB|V81.4|Screen-respir cond NEC
C0260959|ICD9CM|PT|V81.5|Screening for nephropathy
C0260959|ICD9CM|AB|V81.5|Screen for nephropathy
C0260960|ICD9CM|PT|V81.6|Screening for other and unspecified genitourinary conditions
C0260960|ICD9CM|AB|V81.6|Screen for gu cond NEC
C0260961|ICD9CM|HT|V82|Special screening for other conditions
C0260962|ICD9CM|PT|V82.0|Screening for skin conditions
C0260962|ICD9CM|AB|V82.0|Screen for skin cond
C0260963|ICD9CM|PT|V82.1|Screening for rheumatoid arthritis
C0260963|ICD9CM|AB|V82.1|Screen-rheumatoid arthr
C0260964|ICD9CM|PT|V82.2|Screening for other rheumatic disorders
C0260964|ICD9CM|AB|V82.2|Screen-rheumat dis NEC
C0260965|ICD9CM|PT|V82.3|Screening for congenital dislocation of hip
C0260965|ICD9CM|AB|V82.3|Screen-cong hip dislocat
C0260967|ICD9CM|PT|V82.5|Screening for chemical poisoning and other contamination
C0260967|ICD9CM|AB|V82.5|Screen-contamination NEC
C0260968|ICD9CM|PT|V82.9|Screening for unspecified condition
C0260968|ICD9CM|AB|V82.9|Screen for condition NOS
C0260969|ICD9CM|HT|E800|Railway accident involving collision with rolling stock
C0260970|ICD9CM|PT|E800.0|Railway accident involving collision with rolling stock and injuring railway employee
C0260970|ICD9CM|AB|E800.0|RR collision NOS-employ
C0260971|ICD9CM|PT|E800.1|Railway accident involving collision with rolling stock and injuring passenger on railway
C0260971|ICD9CM|AB|E800.1|RR coll NOS-passenger
C0260972|ICD9CM|PT|E800.2|Railway accident involving collision with rolling stock and injuring pedestrian
C0260972|ICD9CM|AB|E800.2|RR coll NOS-pedestrian
C0260973|ICD9CM|PT|E800.3|Railway accident involving collision with rolling stock and injuring pedal cyclist
C0260973|ICD9CM|AB|E800.3|RR coll NOS-ped cyclist
C0260974|ICD9CM|PT|E800.8|Railway accident involving collision with rolling stock and injuring other specified person
C0260974|ICD9CM|AB|E800.8|RR coll NOS-person NEC
C0260975|ICD9CM|PT|E800.9|Railway accident involving collision with rolling stock and injuring unspecified person
C0260975|ICD9CM|AB|E800.9|RR coll NOS-person NOS
C0260976|ICD9CM|HT|E801|Railway accident involving collision with other object
C0260977|ICD9CM|PT|E801.0|Railway accident involving collision with other object and injuring railway employee
C0260977|ICD9CM|AB|E801.0|RR coll w oth obj-employ
C0260978|ICD9CM|PT|E801.1|Railway accident involving collision with other object and injuring passenger on railway
C0260978|ICD9CM|AB|E801.1|RR coll w oth obj-pasngr
C0260979|ICD9CM|PT|E801.2|Railway accident involving collision with other object and injuring pedestrian
C0260979|ICD9CM|AB|E801.2|RR coll w oth obj-pedest
C0260980|ICD9CM|PT|E801.3|Railway accident involving collision with other object and injuring pedal cyclist
C0260980|ICD9CM|AB|E801.3|RR coll w oth obj-cycl
C0260981|ICD9CM|PT|E801.8|Railway accident involving collision with other object and injuring other specified person
C0260981|ICD9CM|AB|E801.8|RR col w oth obj-per NEC
C0260982|ICD9CM|PT|E801.9|Railway accident involving collision with other object and injuring unspecified person
C0260982|ICD9CM|AB|E801.9|RR col w oth obj-per NOS
C0260983|ICD9CM|HT|E802|Railway accident involving derailment without antecedent collision
C0260984|ICD9CM|PT|E802.0|Railway accident involving derailment without antecedent collision injuring railway employee
C0260984|ICD9CM|AB|E802.0|RR acc w derail-employee
C0260985|ICD9CM|PT|E802.1|Railway accident involving derailment without antecedent collision injuring passenger on railway
C0260985|ICD9CM|AB|E802.1|RR acc w derail-passeng
C0260986|ICD9CM|PT|E802.2|Railway accident involving derailment without antecedent collision injuring pedestrian
C0260986|ICD9CM|AB|E802.2|RR acc w derail-pedest
C0260987|ICD9CM|PT|E802.3|Railway accident involving derailment without antecedent collision injuring pedal cyclist
C0260987|ICD9CM|AB|E802.3|RR acc w derail-ped cycl
C0260988|ICD9CM|PT|E802.8|Railway accident involving derailment without antecedent collision injuring other specified person
C0260988|ICD9CM|AB|E802.8|RR acc w derail-pers NEC
C0260989|ICD9CM|PT|E802.9|Railway accident involving derailment without antecedent collision injuring unspecified person
C0260989|ICD9CM|AB|E802.9|RR acc w derail-pers NOS
C0260990|ICD9CM|HT|E803|Railway accident involving explosion, fire, or burning
C0260991|ICD9CM|PT|E803.0|Railway accident involving explosion, fire, or burning injuring railway employee
C0260991|ICD9CM|AB|E803.0|RR acc w explosion-empl
C0260992|ICD9CM|PT|E803.1|Railway accident involving explosion, fire, or burning injuring passenger on railway
C0260992|ICD9CM|AB|E803.1|RR acc w explos-pasngr
C0260993|ICD9CM|PT|E803.2|Railway accident involving explosion, fire, or burning injuring pedestrian
C0260993|ICD9CM|AB|E803.2|RR acc w explos-pedest
C0260994|ICD9CM|PT|E803.3|Railway accident involving explosion, fire, or burning injuring pedal cyclist
C0260994|ICD9CM|AB|E803.3|RR acc w explos-ped cycl
C0260995|ICD9CM|PT|E803.8|Railway accident involving explosion, fire, or burning injuring other specified person
C0260995|ICD9CM|AB|E803.8|RR acc w explos-pers NEC
C0260996|ICD9CM|PT|E803.9|Railway accident involving explosion, fire, or burning injuring unspecified person
C0260996|ICD9CM|AB|E803.9|RR acc w explos-pers NOS
C0260999|ICD9CM|PT|E804.1|Fall in, on, or from railway train injuring passenger on railway
C0260999|ICD9CM|AB|E804.1|Fall from train-passengr
C0261005|ICD9CM|PT|E805.0|Railway employee hit by rolling stock
C0261005|ICD9CM|AB|E805.0|Hit by train-employee
C0261006|ICD9CM|PT|E805.1|Passenger on railway hit by rolling stock
C0261006|ICD9CM|AB|E805.1|Hit by train-passenger
C0261007|ICD9CM|PT|E805.2|Pedestrian hit by rolling stock
C0261007|ICD9CM|AB|E805.2|Hit by train-pedestrian
C0261008|ICD9CM|PT|E805.3|Pedal cyclist hit by rolling stock
C0261008|ICD9CM|AB|E805.3|Hit by train-ped cyclist
C0261009|ICD9CM|PT|E805.8|Other specified person hit by rolling stock
C0261009|ICD9CM|AB|E805.8|Hit by train-person NEC
C0261010|ICD9CM|PT|E805.9|Unspecified person hit by rolling stock
C0261010|ICD9CM|AB|E805.9|Hit by train-person NOS
C0261011|ICD9CM|HT|E806|Other specified railway accident
C0261012|ICD9CM|PT|E806.0|Other specified railway accident injuring railway employee
C0261012|ICD9CM|AB|E806.0|RR acc NEC-employee
C0261013|ICD9CM|PT|E806.1|Other specified railway accident injuring passenger on railway
C0261013|ICD9CM|AB|E806.1|RR acc NEC-passenger
C0261014|ICD9CM|PT|E806.2|Other specified railway accident injuring pedestrian
C0261014|ICD9CM|AB|E806.2|RR acc NEC-pedestrian
C0261015|ICD9CM|PT|E806.3|Other specified railway accident injuring pedal cyclist
C0261015|ICD9CM|AB|E806.3|RR acc NEC-ped cyclist
C0261016|ICD9CM|PT|E806.8|Other specified railway accident injuring other specified person
C0261016|ICD9CM|AB|E806.8|RR acc NEC-person NEC
C0261017|ICD9CM|PT|E806.9|Other specified railway accident injuring unspecified person
C0261017|ICD9CM|AB|E806.9|RR acc NEC-person NOS
C0261019|ICD9CM|PT|E807.0|Railway accident of unspecified nature injuring railway employee
C0261019|ICD9CM|AB|E807.0|RR accident NOS-employee
C0261020|ICD9CM|PT|E807.1|Railway accident of unspecified nature injuring passenger on railway
C0261020|ICD9CM|AB|E807.1|RR acc NOS-passenger
C0261021|ICD9CM|PT|E807.2|Railway accident of unspecified nature injuring pedestrian
C0261021|ICD9CM|AB|E807.2|RR acc NOS-pedestrian
C0261022|ICD9CM|PT|E807.3|Railway accident of unspecified nature injuring pedal cyclist
C0261022|ICD9CM|AB|E807.3|RR acc NOS-ped cyclist
C0261023|ICD9CM|PT|E807.8|Railway accident of unspecified nature injuring other specified person
C0261023|ICD9CM|AB|E807.8|RR acc NOS-person NEC
C0261024|ICD9CM|PT|E807.9|Railway accident of unspecified nature injuring unspecified person
C0261024|ICD9CM|AB|E807.9|RR acc NOS-person NOS
C0261026|ICD9CM|PT|E810.0|Motor vehicle traffic accident involving collision with train injuring driver of motor vehicle other than motorcycle
C0261026|ICD9CM|AB|E810.0|Mv-train coll-driver
C0261027|ICD9CM|PT|E810.1|Motor vehicle traffic accident involving collision with train injuring passenger in motor vehicle other than motorcycle
C0261027|ICD9CM|AB|E810.1|Mv-train coll-pasngr
C0261028|ICD9CM|PT|E810.2|Motor vehicle traffic accident involving collision with train injuring motorcyclist
C0261028|ICD9CM|AB|E810.2|Mv-train coll-motorcycl
C0261029|ICD9CM|PT|E810.3|Motor vehicle traffic accident involving collision with train injuring passenger on motorcycle
C0261029|ICD9CM|AB|E810.3|Mv-train coll-mcycl psgr
C0261030|ICD9CM|PT|E810.4|Motor vehicle traffic accident involving collision with train injuring occupant of streetcar
C0261030|ICD9CM|AB|E810.4|Mv-train coll-st car
C0261031|ICD9CM|PT|E810.5|Motor vehicle traffic accident involving collision with train injuring rider of animal; occupant of animal-drawn vehicle
C0261031|ICD9CM|AB|E810.5|Mv-train coll-anim rid
C0261036|ICD9CM|HT|E811|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle
C0261037|ICD9CM|PT|E811.0|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle injuring driver of motor vehicle other than motorcycle
C0261037|ICD9CM|AB|E811.0|Reentrant mv coll-driver
C0261038|ICD9CM|PT|E811.1|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle injuring passenger in motor vehicle other than motorcycle
C0261038|ICD9CM|AB|E811.1|Reentrant mv coll-pasngr
C0261039|ICD9CM|PT|E811.2|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle injuring motorcyclist
C0261039|ICD9CM|AB|E811.2|Reentrant coll-motcycl
C0261040|ICD9CM|PT|E811.3|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle injuring passenger on motorcycle
C0261040|ICD9CM|AB|E811.3|Reentrant coll-mcyc psgr
C0261041|ICD9CM|PT|E811.4|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle injuring occupant of streetcar
C0261041|ICD9CM|AB|E811.4|Reentrant coll-st car
C0261042|ICD9CM|PT|E811.5|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle injuring rider of animal; occupant of animal-drawn vehicle
C0261042|ICD9CM|AB|E811.5|Reentrant coll-anim rid
C0261043|ICD9CM|PT|E811.6|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle injuring pedal cyclist
C0261043|ICD9CM|AB|E811.6|Reentrant coll-ped cycl
C0261045|ICD9CM|PT|E811.8|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle injuring other specified person
C0261045|ICD9CM|AB|E811.8|Reentrant coll-pers NEC
C0261046|ICD9CM|PT|E811.9|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle injuring unspecified person
C0261046|ICD9CM|AB|E811.9|Reentrant coll-pers NOS
C0261047|ICD9CM|HT|E812|Other motor vehicle traffic accident involving collision with motor vehicle
C0261048|ICD9CM|PT|E812.0|Other motor vehicle traffic accident involving collision with motor vehicle injuring driver of motor vehicle other than motorcycle
C0261048|ICD9CM|AB|E812.0|Mv collision NOS-driver
C0261049|ICD9CM|PT|E812.1|Other motor vehicle traffic accident involving collision with motor vehicle injuring passenger in motor vehicle other than motorcycle
C0261049|ICD9CM|AB|E812.1|Mv collision NOS-pasngr
C0261050|ICD9CM|PT|E812.2|Other motor vehicle traffic accident involving collision with motor vehicle injuring motorcyclist
C0261050|ICD9CM|AB|E812.2|Mv collis NOS-motorcycl
C0261051|ICD9CM|PT|E812.3|Other motor vehicle traffic accident involving collision with motor vehicle injuring passenger on motorcycle
C0261051|ICD9CM|AB|E812.3|Mv coll NOS-mcycl psngr
C0261052|ICD9CM|PT|E812.4|Other motor vehicle traffic accident involving collision with motor vehicle injuring occupant of streetcar
C0261052|ICD9CM|AB|E812.4|Mv collision NOS-st car
C0261053|ICD9CM|PT|E812.5|Other motor vehicle traffic accident involving collision with motor vehicle injuring rider of animal; occupant of animal-drawn vehicle
C0261053|ICD9CM|AB|E812.5|Mv coll NOS-anim rid
C0261054|ICD9CM|PT|E812.6|Other motor vehicle traffic accident involving collision with motor vehicle injuring pedal cyclist
C0261054|ICD9CM|AB|E812.6|Mv coll NOS-ped cycl
C0261055|ICD9CM|PT|E812.7|Other motor vehicle traffic accident involving collision with motor vehicle injuring pedestrian
C0261055|ICD9CM|AB|E812.7|Mv collision NOS-pedest
C0261056|ICD9CM|PT|E812.8|Other motor vehicle traffic accident involving collision with motor vehicle injuring other specified person
C0261056|ICD9CM|AB|E812.8|Mv collis NOS-pers NEC
C0261057|ICD9CM|PT|E812.9|Other motor vehicle traffic accident involving collision with motor vehicle injuring unspecified person
C0261057|ICD9CM|AB|E812.9|Mv collis NOS-pers NOS
C0261058|ICD9CM|HT|E813|Motor vehicle traffic accident involving collision with other vehicle
C0261059|ICD9CM|PT|E813.0|Motor vehicle traffic accident involving collision with other vehicle injuring driver of motor vehicle other than motorcycle
C0261059|ICD9CM|AB|E813.0|Mv-oth veh coll-driver
C0261060|ICD9CM|PT|E813.1|Motor vehicle traffic accident involving collision with other vehicle injuring passenger in motor vehicle other than motorcycle
C0261060|ICD9CM|AB|E813.1|Mv-oth veh coll-pasngr
C0261061|ICD9CM|PT|E813.2|Motor vehicle traffic accident involving collision with other vehicle injuring motorcyclist
C0261061|ICD9CM|AB|E813.2|Mv-oth veh coll-motcycl
C0261062|ICD9CM|PT|E813.3|Motor vehicle traffic accident involving collision with other vehicle injuring passenger on motorcycle
C0261062|ICD9CM|AB|E813.3|Mv-oth veh coll-mcyc psg
C0261063|ICD9CM|PT|E813.4|Motor vehicle traffic accident involving collision with other vehicle injuring occupant of streetcar
C0261063|ICD9CM|AB|E813.4|Mv-oth veh coll-st car
C0261064|ICD9CM|PT|E813.5|Motor vehicle traffic accident involving collision with other vehicle injuring rider of animal; occupant of animal-drawn vehicle
C0261064|ICD9CM|AB|E813.5|Mv-oth veh coll-anim rid
C0261065|ICD9CM|PT|E813.6|Motor vehicle traffic accident involving collision with other vehicle injuring pedal cyclist
C0261065|ICD9CM|AB|E813.6|Mv-oth veh coll-ped cycl
C0261066|ICD9CM|PT|E813.7|Motor vehicle traffic accident involving collision with other vehicle injuring pedestrian
C0261066|ICD9CM|AB|E813.7|Mv-oth veh coll-pedest
C0261067|ICD9CM|PT|E813.8|Motor vehicle traffic accident involving collision with other vehicle injuring other specified person
C0261067|ICD9CM|AB|E813.8|Mv-oth veh coll-pers NEC
C0261069|ICD9CM|HT|E814|Motor vehicle traffic accident involving collision with pedestrian
C0261070|ICD9CM|PT|E814.0|Motor vehicle traffic accident involving collision with pedestrian injuring driver of motor vehicle other than motorcycle
C0261070|ICD9CM|AB|E814.0|Mv coll w pedest-driver
C0261071|ICD9CM|PT|E814.1|Motor vehicle traffic accident involving collision with pedestrian injuring passenger in motor vehicle other than motorcycle
C0261071|ICD9CM|AB|E814.1|Mv coll w pedest-pasngr
C0261072|ICD9CM|PT|E814.2|Motor vehicle traffic accident involving collision with pedestrian injuring motorcyclist
C0261072|ICD9CM|AB|E814.2|Mv coll w pedest-motcycl
C0261073|ICD9CM|PT|E814.3|Motor vehicle traffic accident involving collision with pedestrian injuring passenger on motorcycle
C0261073|ICD9CM|AB|E814.3|Mv coll w ped-mcycl psgr
C0261074|ICD9CM|PT|E814.4|Motor vehicle traffic accident involving collision with pedestrian injuring occupant of streetcar
C0261074|ICD9CM|AB|E814.4|Mv coll w pedest-st car
C0261075|ICD9CM|PT|E814.5|Motor vehicle traffic accident involving collision with pedestrian injuring rider of animal; occupant of animal drawn vehicle
C0261075|ICD9CM|AB|E814.5|Mv coll w ped-anim rid
C0261076|ICD9CM|PT|E814.6|Motor vehicle traffic accident involving collision with pedestrian injuring pedal cyclist
C0261076|ICD9CM|AB|E814.6|Mv coll w ped-ped cycl
C0261077|ICD9CM|PT|E814.7|Motor vehicle traffic accident involving collision with pedestrian injuring pedestrian
C0261077|ICD9CM|AB|E814.7|Mv coll w pedest-pedest
C0261078|ICD9CM|PT|E814.8|Motor vehicle traffic accident involving collision with pedestrian injuring other specified person
C0261078|ICD9CM|AB|E814.8|Mv coll w pedes-pers NEC
C0261079|ICD9CM|PT|E814.9|Motor vehicle traffic accident involving collision with pedestrian injuring unspecified person
C0261079|ICD9CM|AB|E814.9|Mv coll w pedes-pers NOS
C0261080|ICD9CM|HT|E815|Other motor vehicle traffic accident involving collision on the highway
C0261081|ICD9CM|PT|E815.0|Other motor vehicle traffic accident involving collision on the highway injuring driver of motor vehicle other than motorcycle
C0261081|ICD9CM|AB|E815.0|Mv coll w oth obj-driver
C0261082|ICD9CM|PT|E815.1|Other motor vehicle traffic accident involving collision on the highway injuring passenger in motor vehicle other than motorcycle
C0261082|ICD9CM|AB|E815.1|Mv coll w oth obj-pasngr
C0261083|ICD9CM|PT|E815.2|Other motor vehicle traffic accident involving collision on the highway injuring motorcyclist
C0261083|ICD9CM|AB|E815.2|Mv coll w oth obj-mocycl
C0261084|ICD9CM|PT|E815.3|Other motor vehicle traffic accident involving collision on the highway injuring passenger on motorcycle
C0261084|ICD9CM|AB|E815.3|Mv coll w obj-mcycl psgr
C0261085|ICD9CM|PT|E815.4|Other motor vehicle traffic accident involving collision on the highway injuring occupant of streetcar
C0261085|ICD9CM|AB|E815.4|Mv coll w obj-st car
C0261086|ICD9CM|PT|E815.5|Other motor vehicle traffic accident involving collision on the highway injuring rider of animal; occupant of animal-drawn vehicle
C0261086|ICD9CM|AB|E815.5|Mv coll w obj-anim rider
C0261087|ICD9CM|PT|E815.6|Other motor vehicle traffic accident involving collision on the highway injuring pedal cyclist
C0261087|ICD9CM|AB|E815.6|Mv coll w obj-ped cycl
C0261088|ICD9CM|PT|E815.7|Other motor vehicle traffic accident involving collision on the highway injuring pedestrian
C0261088|ICD9CM|AB|E815.7|Mv coll w obj-pedest
C0261089|ICD9CM|PT|E815.8|Other motor vehicle traffic accident involving collision on the highway injuring other specified person
C0261089|ICD9CM|AB|E815.8|Mv coll w obj-pers NEC
C0261090|ICD9CM|PT|E815.9|Other motor vehicle traffic accident involving collision on the highway injuring unspecified person
C0261090|ICD9CM|AB|E815.9|Mv coll w obj-pers NOS
C0261091|ICD9CM|HT|E816|Motor vehicle traffic accident due to loss of control, without collision on the highway
C0261092|ICD9CM|PT|E816.0|Motor vehicle traffic accident due to loss of control, without collision on the highway, injuring driver of motor vehicle other than motorcycle
C0261092|ICD9CM|AB|E816.0|Loss control mv acc-driv
C0261093|ICD9CM|PT|E816.1|Motor vehicle traffic accident due to loss of control, without collision on the highway, injuring passenger in motor vehicle other than motorcycle
C0261093|ICD9CM|AB|E816.1|Loss control mv acc-psgr
C0261095|ICD9CM|PT|E816.3|Motor vehicle traffic accident due to loss of control, without collision on the highway, injuring passenger on motorcycle
C0261095|ICD9CM|AB|E816.3|Loss control mv-mcyc psg
C0261096|ICD9CM|PT|E816.4|Motor vehicle traffic accident due to loss of control, without collision on the highway, injuring occupant of streetcar
C0261096|ICD9CM|AB|E816.4|Loss cont mv acc-st car
C0261097|ICD9CM|PT|E816.5|Motor vehicle traffic accident due to loss of control, without collision on the highway, injuring rider of animal; occupant of animal-drawn vehicle
C0261097|ICD9CM|AB|E816.5|Loss cont mv-anim rider
C0261102|ICD9CM|HT|E817|Noncollision motor vehicle traffic accident while boarding or alighting
C0261103|ICD9CM|PT|E817.0|Noncollision motor vehicle traffic accident while boarding or alighting injuring driver of motor vehicle other than motorcycle
C0261103|ICD9CM|AB|E817.0|Mv acc board/alight-driv
C0261104|ICD9CM|PT|E817.1|Noncollision motor vehicle traffic accident while boarding or alighting injuring passenger in motor vehicle other than motorcycle
C0261104|ICD9CM|AB|E817.1|Mv acc board/alight-psgr
C0261105|ICD9CM|PT|E817.2|Noncollision motor vehicle traffic accident while boarding or alighting injuring motorcyclist
C0261105|ICD9CM|AB|E817.2|Mv board/alight-motcycl
C0261106|ICD9CM|PT|E817.3|Noncollision motor vehicle traffic accident while boarding or alighting injuring passenger on motorcycle
C0261106|ICD9CM|AB|E817.3|Mv brd/alight-mcycl psgr
C0261107|ICD9CM|PT|E817.4|Noncollision motor vehicle traffic accident while boarding or alighting injuring occupant of streetcar
C0261107|ICD9CM|AB|E817.4|Mv acc brd/alight-st car
C0261108|ICD9CM|PT|E817.5|Noncollision motor vehicle traffic accident while boarding or alighting injuring rider of animal; occupant of animal-drawn vehicle
C0261108|ICD9CM|AB|E817.5|Mv brd/alight-anim rider
C0261109|ICD9CM|PT|E817.6|Noncollision motor vehicle traffic accident while boarding or alighting injuring pedal cyclist
C0261109|ICD9CM|AB|E817.6|Mv brd/alight-ped cycl
C0261110|ICD9CM|PT|E817.7|Noncollision motor vehicle traffic accident while boarding or alighting injuring pedestrian
C0261110|ICD9CM|AB|E817.7|Mv brd/alight-pedestrian
C0261111|ICD9CM|PT|E817.8|Noncollision motor vehicle traffic accident while boarding or alighting injuring other specified person
C0261111|ICD9CM|AB|E817.8|Mv board/alight-pers NEC
C0261112|ICD9CM|PT|E817.9|Noncollision motor vehicle traffic accident while boarding or alighting injuring unspecified person
C0261112|ICD9CM|AB|E817.9|Mv board/alight-pers NOS
C0261113|ICD9CM|HT|E818|Other noncollision motor vehicle traffic accident
C0261114|ICD9CM|PT|E818.0|Other noncollision motor vehicle traffic accident injuring driver of motor vehicle other than motorcycle
C0261114|ICD9CM|AB|E818.0|Mv traff acc NEC-driver
C0261115|ICD9CM|PT|E818.1|Other noncollision motor vehicle traffic accident injuring passenger in motor vehicle other than motorcycle
C0261115|ICD9CM|AB|E818.1|Mv traff acc NEC-pasngr
C0261116|ICD9CM|PT|E818.2|Other noncollision motor vehicle traffic accident injuring motorcyclist
C0261116|ICD9CM|AB|E818.2|Mv traff acc NEC-mocycl
C0261117|ICD9CM|PT|E818.3|Other noncollision motor vehicle traffic accident injuring passenger on motorcycle
C0261117|ICD9CM|AB|E818.3|Mv traff acc-mcycl psgr
C0261118|ICD9CM|PT|E818.4|Other noncollision motor vehicle traffic accident injuring occupant of streetcar
C0261118|ICD9CM|AB|E818.4|Mv traff acc NEC-st car
C0261119|ICD9CM|PT|E818.5|Other noncollision motor vehicle traffic accident injuring rider of animal; occupant of animal-drawn vehicle
C0261119|ICD9CM|AB|E818.5|Mv traff acc-anim rider
C0261120|ICD9CM|PT|E818.6|Other noncollision motor vehicle traffic accident injuring pedal cyclist
C0261120|ICD9CM|AB|E818.6|Mv traff acc-ped cyc
C0261121|ICD9CM|PT|E818.7|Other noncollision motor vehicle traffic accident injuring pedestrian
C0261121|ICD9CM|AB|E818.7|Mv traff acc NEC-pedest
C0261122|ICD9CM|PT|E818.8|Other noncollision motor vehicle traffic accident injuring other specified person
C0261122|ICD9CM|AB|E818.8|Mv traff acc-pers NEC
C0261123|ICD9CM|PT|E818.9|Other noncollision motor vehicle traffic accident injuring unspecified person
C0261123|ICD9CM|AB|E818.9|Mv traff acc-pers NOS
C0261124|ICD9CM|PT|E819.0|Motor vehicle traffic accident of unspecified nature injuring driver of motor vehicle other than motorcycle
C0261124|ICD9CM|AB|E819.0|Traffic acc NOS-driver
C0261125|ICD9CM|PT|E819.1|Motor vehicle traffic accident of unspecified nature injuring passenger in motor vehicle other than motorcycle
C0261125|ICD9CM|AB|E819.1|Traffic acc NOS-pasngr
C0261126|ICD9CM|PT|E819.2|Motor vehicle traffic accident of unspecified nature injuring motorcyclist
C0261126|ICD9CM|AB|E819.2|Traffic acc NOS-motcycl
C0261127|ICD9CM|PT|E819.3|Motor vehicle traffic accident of unspecified nature injuring passenger on motorcycle
C0261127|ICD9CM|AB|E819.3|Traff acc NOS-mcycl psgr
C0261128|ICD9CM|PT|E819.4|Motor vehicle traffic accident of unspecified nature injuring occupant of streetcar
C0261128|ICD9CM|AB|E819.4|Traffic acc NOS-st car
C0261129|ICD9CM|PT|E819.5|Motor vehicle traffic accident of unspecified nature injuring rider of animal; occupant of animal-drawn vehicle
C0261129|ICD9CM|AB|E819.5|Traff acc NOS-anim rider
C0261130|ICD9CM|PT|E819.6|Motor vehicle traffic accident of unspecified nature injuring pedal cyclist
C0261130|ICD9CM|AB|E819.6|Traffic acc NOS-ped cycl
C0261131|ICD9CM|PT|E819.7|Motor vehicle traffic accident of unspecified nature injuring pedestrian
C0261131|ICD9CM|AB|E819.7|Traffic acc NOS-pedest
C0261132|ICD9CM|PT|E819.8|Motor vehicle traffic accident of unspecified nature injuring other specified person
C0261132|ICD9CM|AB|E819.8|Traffic acc NOS-pers NEC
C0261133|ICD9CM|PT|E819.9|Motor vehicle traffic accident of unspecified nature injuring unspecified person
C0261133|ICD9CM|AB|E819.9|Traffic acc NOS-pers NOS
C0261135|ICD9CM|PT|E820.0|Nontraffic accident involving motor-driven snow vehicle injuring driver of motor vehicle other than motorcycle
C0261135|ICD9CM|AB|E820.0|Snow veh acc-driver
C0261136|ICD9CM|PT|E820.1|Nontraffic accident involving motor-driven snow vehicle injuring passenger in motor vehicle other than motorcycle
C0261136|ICD9CM|AB|E820.1|Snow veh acc-pasngr
C0261137|ICD9CM|PT|E820.2|Nontraffic accident involving motor-driven snow vehicle injuring motorcyclist
C0261137|ICD9CM|AB|E820.2|Snow veh acc-motorcycl
C0261138|ICD9CM|PT|E820.3|Nontraffic accident involving motor-driven snow vehicle injuring passenger on motorcycle
C0261138|ICD9CM|AB|E820.3|Snow veh acc-mcycl psgr
C0261139|ICD9CM|PT|E820.4|Nontraffic accident involving motor-driven snow vehicle injuring occupant of streetcar
C0261139|ICD9CM|AB|E820.4|Snow veh acc-st car
C0261140|ICD9CM|PT|E820.5|Nontraffic accident involving motor-driven snow vehicle injuring rider of animal; occupant of animal-drawn vehicle
C0261140|ICD9CM|AB|E820.5|Snow veh acc-anim rider
C0261141|ICD9CM|PT|E820.6|Nontraffic accident involving motor-driven snow vehicle injuring pedal cyclist
C0261141|ICD9CM|AB|E820.6|Snow veh acc-ped cycl
C0261142|ICD9CM|PT|E820.7|Nontraffic accident involving motor-driven snow vehicle injuring pedestrian
C0261142|ICD9CM|AB|E820.7|Snow veh acc-pedest
C0261143|ICD9CM|PT|E820.8|Nontraffic accident involving motor-driven snow vehicle injuring other specified person
C0261143|ICD9CM|AB|E820.8|Snow veh acc-pers NEC
C0261144|ICD9CM|PT|E820.9|Nontraffic accident involving motor-driven snow vehicle injuring unspecified person
C0261144|ICD9CM|AB|E820.9|Snow veh acc-pers NOS
C0261145|ICD9CM|HT|E821|Nontraffic accident involving other off-road motor vehicle
C0261146|ICD9CM|PT|E821.0|Nontraffic accident involving other off-road motor vehicle injuring driver of motor vehicle other than motorcycle
C0261146|ICD9CM|AB|E821.0|Oth off-road mv acc-driv
C0261147|ICD9CM|PT|E821.1|Nontraffic accident involving other off-road motor vehicle injuring passenger in motor vehicle other than motorcycle
C0261147|ICD9CM|AB|E821.1|Oth off-road mv acc-psgr
C0261148|ICD9CM|PT|E821.2|Nontraffic accident involving other off-road motor vehicle injuring motorcyclist
C0261148|ICD9CM|AB|E821.2|Oth off-road mv-mocycl
C0261149|ICD9CM|PT|E821.3|Nontraffic accident involving other off-road motor vehicle injuring passenger on motorcycle
C0261149|ICD9CM|AB|E821.3|Oth off-road mv-mcyc psg
C0261150|ICD9CM|PT|E821.4|Nontraffic accident involving other off-road motor vehicle injuring occupant of streetcar
C0261150|ICD9CM|AB|E821.4|Oth off-road mv-st car
C0261151|ICD9CM|PT|E821.5|Nontraffic accident involving other off-road motor vehicle injuring rider of animal; occupant of animal-drawn vehicle
C0261151|ICD9CM|AB|E821.5|Oth off-road mv-anim rid
C0261152|ICD9CM|PT|E821.6|Nontraffic accident involving other off-road motor vehicle injuring pedal cyclist
C0261152|ICD9CM|AB|E821.6|Oth off-road mv-ped cycl
C0261153|ICD9CM|PT|E821.7|Nontraffic accident involving other off-road motor vehicle injuring pedestrian
C0261153|ICD9CM|AB|E821.7|Oth off-road mv-pedest
C0261154|ICD9CM|PT|E821.8|Nontraffic accident involving other off-road motor vehicle injuring other specified person
C0261154|ICD9CM|AB|E821.8|Oth off-road mv-pers NEC
C0261155|ICD9CM|PT|E821.9|Nontraffic accident involving other off-road motor vehicle injuring unspecified person
C0261155|ICD9CM|AB|E821.9|Oth off-road mv-pers NOS
C0261156|ICD9CM|HT|E822|Other motor vehicle nontraffic accident involving collision with moving object
C0261157|ICD9CM|PT|E822.0|Other motor vehicle nontraffic accident involving collision with moving object injuring driver of motor vehicle other than motorcycle
C0261157|ICD9CM|AB|E822.0|Oth coll w mov obj-driv
C0261158|ICD9CM|PT|E822.1|Other motor vehicle nontraffic accident involving collision with moving object injuring passenger in motor vehicle other than motorcycle
C0261158|ICD9CM|AB|E822.1|Oth coll w mov obj-psgr
C0261159|ICD9CM|PT|E822.2|Other motor vehicle nontraffic accident involving collision with moving object injuring motorcyclist
C0261159|ICD9CM|AB|E822.2|Oth coll mov obj-mocycl
C0261160|ICD9CM|PT|E822.3|Other motor vehicle nontraffic accident involving collision with moving object injuring passenger on motorcycle
C0261160|ICD9CM|AB|E822.3|Oth coll mov obj-cyc psg
C0261161|ICD9CM|PT|E822.4|Other motor vehicle nontraffic accident involving collision with moving object injuring occupant of streetcar
C0261161|ICD9CM|AB|E822.4|Oth coll mov obj-st car
C0261162|ICD9CM|PT|E822.5|Other motor vehicle nontraffic accident involving collision with moving object injuring rider of animal; occupant of animal-drawn vehicle
C0261162|ICD9CM|AB|E822.5|Oth coll mov obj-rider
C0261163|ICD9CM|PT|E822.6|Other motor vehicle nontraffic accident involving collision with moving object injuring pedal cyclist
C0261163|ICD9CM|AB|E822.6|Oth coll mov obj-ped cyc
C0261164|ICD9CM|PT|E822.7|Other motor vehicle nontraffic accident involving collision with moving object injuring pedestrian
C0261164|ICD9CM|AB|E822.7|Oth coll mov obj-pedest
C0261165|ICD9CM|PT|E822.8|Other motor vehicle nontraffic accident involving collision with moving object injuring other specified person
C0261165|ICD9CM|AB|E822.8|Oth coll mov obj-per NEC
C0261166|ICD9CM|PT|E822.9|Other motor vehicle nontraffic accident involving collision with moving object injuring unspecified person
C0261166|ICD9CM|AB|E822.9|Oth coll mov obj-per NOS
C0261167|ICD9CM|HT|E823|Other motor vehicle nontraffic accident involving collision with stationary object
C0261168|ICD9CM|PT|E823.0|Other motor vehicle nontraffic accident involving collision with stationary object injuring driver of motor vehicle other than motorcycle
C0261168|ICD9CM|AB|E823.0|Oth coll stndng obj-driv
C0261169|ICD9CM|PT|E823.1|Other motor vehicle nontraffic accident involving collision with stationary object injuring passenger in motor vehicle other than motorcycle
C0261169|ICD9CM|AB|E823.1|Oth coll stndng obj-psgr
C0261170|ICD9CM|PT|E823.2|Other motor vehicle nontraffic accident involving collision with stationary object injuring motorcyclist
C0261170|ICD9CM|AB|E823.2|Oth coll stnd obj-mocycl
C0261171|ICD9CM|PT|E823.3|Other motor vehicle nontraffic accident involving collision with stationary object injuring passenger on motorcycle
C0261171|ICD9CM|AB|E823.3|Oth coll stn obj-cyc psg
C0261172|ICD9CM|PT|E823.4|Other motor vehicle nontraffic accident involving collision with stationary object injuring occupant of streetcar
C0261172|ICD9CM|AB|E823.4|Oth coll stnd obj-st car
C0261173|ICD9CM|PT|E823.5|Other motor vehicle nontraffic accident involving collision with stationary object injuring rider of animal; occupant of animal-drawn vehicle
C0261173|ICD9CM|AB|E823.5|Oth coll stnd obj-rider
C0261174|ICD9CM|PT|E823.6|Other motor vehicle nontraffic accident involving collision with stationary object injuring pedal cyclist
C0261174|ICD9CM|AB|E823.6|Oth coll stn obj-ped cyc
C0261175|ICD9CM|PT|E823.7|Other motor vehicle nontraffic accident involving collision with stationary object injuring pedestrian
C0261175|ICD9CM|AB|E823.7|Oth coll stnd obj-pedest
C0261176|ICD9CM|PT|E823.8|Other motor vehicle nontraffic accident involving collision with stationary object injuring other specified person
C0261176|ICD9CM|AB|E823.8|Oth coll stn obj-per NEC
C0261177|ICD9CM|PT|E823.9|Other motor vehicle nontraffic accident involving collision with stationary object injuring unspecified person
C0261177|ICD9CM|AB|E823.9|Oth col-stnd-obj-per NOS
C0261178|ICD9CM|HT|E824|Other motor vehicle nontraffic accident while boarding and alighting
C0261179|ICD9CM|PT|E824.0|Other motor vehicle nontraffic accident while boarding and alighting injuring driver of motor vehicle other than motorcycle
C0261179|ICD9CM|AB|E824.0|N-traf board/alight-driv
C0261180|ICD9CM|PT|E824.1|Other motor vehicle nontraffic accident while boarding and alighting injuring passenger in motor vehicle other than motorcycle
C0261180|ICD9CM|AB|E824.1|N-traf board/alight-psgr
C0261181|ICD9CM|PT|E824.2|Other motor vehicle nontraffic accident while boarding and alighting injuring motorcyclist
C0261181|ICD9CM|AB|E824.2|N-traf brd/alight-mocycl
C0261182|ICD9CM|PT|E824.3|Other motor vehicle nontraffic accident while boarding and alighting injuring passenger on motorcycle
C0261182|ICD9CM|AB|E824.3|N-traf brd/alit-mcyc psg
C0261183|ICD9CM|PT|E824.4|Other motor vehicle nontraffic accident while boarding and alighting injuring occupant of streetcar
C0261183|ICD9CM|AB|E824.4|N-traf brd/alit-st car
C0261184|ICD9CM|PT|E824.5|Other motor vehicle nontraffic accident while boarding and alighting injuring rider of animal; occupant of animal-drawn vehicle
C0261184|ICD9CM|AB|E824.5|N-traf brd/alit-anim rid
C0261185|ICD9CM|PT|E824.6|Other motor vehicle nontraffic accident while boarding and alighting injuring pedal cyclist
C0261185|ICD9CM|AB|E824.6|N-traf brd/alit-ped cycl
C0261186|ICD9CM|PT|E824.7|Other motor vehicle nontraffic accident while boarding and alighting injuring pedestrian
C0261186|ICD9CM|AB|E824.7|N-traf brd/alit-pedest
C0261187|ICD9CM|PT|E824.8|Other motor vehicle nontraffic accident while boarding and alighting injuring other specified person
C0261187|ICD9CM|AB|E824.8|N-traf brd/alit-pers NEC
C0261188|ICD9CM|PT|E824.9|Other motor vehicle nontraffic accident while boarding and alighting injuring unspecified person
C0261188|ICD9CM|AB|E824.9|N-traf brd/alit-pers NOS
C0261189|ICD9CM|HT|E825|Other motor vehicle nontraffic accident of other and unspecified nature
C0261190|ICD9CM|PT|E825.0|Other motor vehicle nontraffic accident of other and unspecified nature injuring driver of motor vehicle other than motorcycle
C0261190|ICD9CM|AB|E825.0|Mv n-traff acc NEC-driv
C0261191|ICD9CM|PT|E825.1|Other motor vehicle nontraffic accident of other and unspecified nature injuring passenger in motor vehicle other than motorcycle
C0261191|ICD9CM|AB|E825.1|Mv n-traff NEC/NOS-psgr
C0261192|ICD9CM|PT|E825.2|Other motor vehicle nontraffic accident of other and unspecified nature injuring motorcyclist
C0261192|ICD9CM|AB|E825.2|Mv n-traf acc NEC-mocycl
C0261193|ICD9CM|PT|E825.3|Other motor vehicle nontraffic accident of other and unspecified nature injuring passenger on motorcycle
C0261193|ICD9CM|AB|E825.3|Mv n-traff NEC-mcyc psgr
C0261194|ICD9CM|PT|E825.4|Other motor vehicle nontraffic accident of other and unspecified nature injuring occupant of streetcar
C0261194|ICD9CM|AB|E825.4|Mv n-traff NEC-st car
C0261195|ICD9CM|PT|E825.5|Other motor vehicle nontraffic accident of other and unspecified nature injuring rider of animal; occupant of animal-drawn vehicle
C0261195|ICD9CM|AB|E825.5|Mv n-traf NEC-anim rider
C0261196|ICD9CM|PT|E825.6|Other motor vehicle nontraffic accident of other and unspecified nature injuring pedal cyclist
C0261196|ICD9CM|AB|E825.6|Mv n-traff NEC-ped cycl
C0261197|ICD9CM|PT|E825.7|Other motor vehicle nontraffic accident of other and unspecified nature injuring pedestrian
C0261197|ICD9CM|AB|E825.7|Mv n-traff NEC-pedest
C0261198|ICD9CM|PT|E825.8|Other motor vehicle nontraffic accident of other and unspecified nature injuring other specified person
C0261198|ICD9CM|AB|E825.8|Mv n-traff NEC-pers NEC
C0261199|ICD9CM|PT|E825.9|Other motor vehicle nontraffic accident of other and unspecified nature injuring unspecified person
C0261199|ICD9CM|AB|E825.9|Mv n-traff NEC-pers NOS
C0261200|ICD9CM|HT|E826|Pedal cycle accident
C0261201|ICD9CM|PT|E826.0|Pedal cycle accident injuring pedestrian
C0261201|ICD9CM|AB|E826.0|Pedal cycle acc-pedest
C0261202|ICD9CM|PT|E826.1|Pedal cycle accident injuring pedal cyclist
C0261202|ICD9CM|AB|E826.1|Ped cycl acc-ped cyclist
C0261203|ICD9CM|PT|E826.2|Pedal cycle accident injuring rider of animal
C0261203|ICD9CM|AB|E826.2|Ped cycle acc-anim rider
C0261205|ICD9CM|PT|E826.4|Pedal cycle accident injuring occupant of streetcar
C0261205|ICD9CM|AB|E826.4|Ped cycle acc-occ st car
C0261206|ICD9CM|PT|E826.8|Pedal cycle accident injuring other specified person
C0261206|ICD9CM|AB|E826.8|Ped cycle acc-pers NEC
C0261207|ICD9CM|PT|E826.9|Pedal cycle accident injuring unspecified person
C0261207|ICD9CM|AB|E826.9|Ped cycle acc-pers NOS
C0261208|ICD9CM|HT|E827|Animal-drawn vehicle accident
C0261209|ICD9CM|PT|E827.0|Animal-drawn vehicle accident injuring pedestrian
C0261209|ICD9CM|AB|E827.0|Animal drawn veh-pedest
C0261210|ICD9CM|PT|E827.2|Animal-drawn vehicle accident injuring rider of animal
C0261210|ICD9CM|AB|E827.2|Anim drawn veh-anim rid
C0261211|ICD9CM|PT|E827.3|Animal-drawn vehicle accident injuring occupant of animal drawn vehicle
C0261211|ICD9CM|AB|E827.3|Animal drawn veh-occupan
C0261212|ICD9CM|PT|E827.4|Animal-drawn vehicle accident injuring occupant of streetcar
C0261212|ICD9CM|AB|E827.4|Anim drawn-occ st car
C0261213|ICD9CM|PT|E827.8|Animal-drawn vehicle accident injuring other specified person
C0261213|ICD9CM|AB|E827.8|Anim drawn veh-pers NEC
C0261214|ICD9CM|PT|E827.9|Animal-drawn vehicle accident injuring unspecified person
C0261214|ICD9CM|AB|E827.9|Anim drawn veh-pers NOS
C0261215|ICD9CM|HT|E828|Accident involving animal being ridden
C0261218|ICD9CM|PT|E828.4|Accident involving animal being ridden injuring occupant of streetcar
C0261218|ICD9CM|AB|E828.4|Ridden animal acc-st car
C0261219|ICD9CM|PT|E828.8|Accident involving animal being ridden injuring other specified person
C0261219|ICD9CM|AB|E828.8|Ridden anim acc-pers NEC
C0261220|ICD9CM|PT|E828.9|Accident involving animal being ridden injuring unspecified person
C0261220|ICD9CM|AB|E828.9|Ridden anim acc-pers NOS
C0261221|ICD9CM|PT|E829.0|Other road vehicle accidents injuring pedestrian
C0261221|ICD9CM|AB|E829.0|Oth road veh acc-pedest
C0261222|ICD9CM|PT|E829.4|Other road vehicle accidents injuring occupant of streetcar
C0261222|ICD9CM|AB|E829.4|Oth rd veh acc-st car
C0261224|ICD9CM|PT|E829.9|Other road vehicle accidents injuring unspecified person
C0261224|ICD9CM|AB|E829.9|Oth rd veh acc-pers NOS
C0261225|ICD9CM|HT|E830|Accident to watercraft causing submersion
C0261226|ICD9CM|PT|E830.0|Accident to watercraft causing submersion injuring occupant of small boat, unpowered
C0261226|ICD9CM|AB|E830.0|Boat acc w submers-unpow
C0261227|ICD9CM|PT|E830.1|Accident to watercraft causing submersion injuring occupant of small boat, powered
C0261227|ICD9CM|AB|E830.1|Boat acc w submers-power
C0261228|ICD9CM|PT|E830.2|Accident to watercraft causing submersion injuring occupant of other watercraft -- crew
C0261228|ICD9CM|AB|E830.2|Boat acc w submers-crew
C0261229|ICD9CM|PT|E830.3|Accident to watercraft causing submersion injuring occupant of other watercraft -- other than crew
C0261229|ICD9CM|AB|E830.3|Boat acc w submers-psgr
C0261230|ICD9CM|PT|E830.4|Accident to watercraft causing submersion injuring water skier
C0261230|ICD9CM|AB|E830.4|Boat submers-water skier
C0261231|ICD9CM|PT|E830.5|Accident to watercraft causing submersion injuring swimmer
C0261231|ICD9CM|AB|E830.5|Boat submers-swimmer
C0261232|ICD9CM|PT|E830.6|Accident to watercraft causing submersion injuring dockers, stevedores
C0261232|ICD9CM|AB|E830.6|Boat submers-dockers
C0261233|ICD9CM|PT|E830.8|Accident to watercraft causing submersion injuring other specified person
C0261233|ICD9CM|AB|E830.8|Boat submers-pers NEC
C0261234|ICD9CM|PT|E830.9|Accident to watercraft causing submersion injuring unspecified person
C0261234|ICD9CM|AB|E830.9|Boat submers-pers NOS
C0261235|ICD9CM|HT|E831|Accident to watercraft causing other injury
C0261236|ICD9CM|PT|E831.0|Accident to watercraft causing other injury to occupant of small boat, unpowered
C0261236|ICD9CM|AB|E831.0|Boat acc inj NEC-unpower
C0261237|ICD9CM|PT|E831.1|Accident to watercraft causing other injury to occupant of small boat, powered
C0261237|ICD9CM|AB|E831.1|Boat acc inj NEC-power
C0261238|ICD9CM|PT|E831.2|Accident to watercraft causing other injury to occupant of other watercraft -- crew
C0261238|ICD9CM|AB|E831.2|Boat acc inj NEC-crew
C0261239|ICD9CM|PT|E831.3|Accident to watercraft causing other injury to occupant of other watercraft -- other than crew
C0261239|ICD9CM|AB|E831.3|Boat acc inj NEC-passeng
C0261240|ICD9CM|PT|E831.4|Accident to watercraft causing other injury to water skier
C0261240|ICD9CM|AB|E831.4|Boat acc inj NEC-skier
C0261241|ICD9CM|PT|E831.5|Accident to watercraft causing other injury to swimmer
C0261241|ICD9CM|AB|E831.5|Boat acc inj NEC-swim
C0261242|ICD9CM|PT|E831.6|Accident to watercraft causing other injury to dockers, stevedores
C0261242|ICD9CM|AB|E831.6|Boat acc inj NEC-docker
C0261243|ICD9CM|PT|E831.8|Accident to watercraft causing other injury to other specified person
C0261243|ICD9CM|AB|E831.8|Boat inj NEC-person NEC
C0261244|ICD9CM|PT|E831.9|Accident to watercraft causing other injury to unspecified person
C0261244|ICD9CM|AB|E831.9|Boat inj NEC-person NOS
C0261245|ICD9CM|HT|E832|Other accidental submersion or drowning in water transport accident
C0261246|ICD9CM|PT|E832.0|Other accidental submersion or drowning in water transport accident injuring occupant of small boat, unpowered
C0261246|ICD9CM|AB|E832.0|Submers NEC-unpow boat
C0261247|ICD9CM|PT|E832.1|Other accidental submersion or drowning in water transport accident injuring occupant of small boat, powered
C0261247|ICD9CM|AB|E832.1|Submers NEC-power boat
C0261248|ICD9CM|PT|E832.2|Other accidental submersion or drowning in water transport accident injuring occupant of other watercraft -- crew
C0261248|ICD9CM|AB|E832.2|Submers NEC-crew
C0261249|ICD9CM|PT|E832.3|Other accidental submersion or drowning in water transport accident injuring occupant of other watercraft -- other than crew
C0261249|ICD9CM|AB|E832.3|Submers NEC-passenger
C0261250|ICD9CM|PT|E832.4|Other accidental submersion or drowning in water transport accident injuring water skier
C0261250|ICD9CM|AB|E832.4|Submers NEC-water skier
C0261251|ICD9CM|PT|E832.5|Other accidental submersion or drowning in water transport accident injuring swimmer
C0261251|ICD9CM|AB|E832.5|Submers NEC-swimmer
C0261252|ICD9CM|PT|E832.6|Other accidental submersion or drowning in water transport accident injuring dockers, stevedores
C0261252|ICD9CM|AB|E832.6|Submers NEC-docker
C0261253|ICD9CM|PT|E832.8|Other accidental submersion or drowning in water transport accident injuring other specified person
C0261253|ICD9CM|AB|E832.8|Submers NEC-person NEC
C0261254|ICD9CM|PT|E832.9|Other accidental submersion or drowning in water transport accident injuring unspecified person
C0261254|ICD9CM|AB|E832.9|Submers NEC-person NOS
C0261255|ICD9CM|HT|E833|Fall on stairs or ladders in water transport
C0261256|ICD9CM|PT|E833.0|Fall on stairs or ladders in water transport injuring occupant of small boat, unpowered
C0261256|ICD9CM|AB|E833.0|W/craft stair fall-unpow
C0261257|ICD9CM|PT|E833.1|Fall on stairs or ladders in water transport injuring occupant of small boat, powered
C0261257|ICD9CM|AB|E833.1|W/craft stair fall-power
C0261258|ICD9CM|PT|E833.2|Fall on stairs or ladders in water transport injuring occupant of other watercraft -- crew
C0261258|ICD9CM|AB|E833.2|Wtrcraft stair fall-crew
C0261259|ICD9CM|PT|E833.3|Fall on stairs or ladders in water transport injuring occupant of other watercraft -- other than crew
C0261259|ICD9CM|AB|E833.3|Wtrcraft stair fall-psgr
C0261260|ICD9CM|PT|E833.4|Fall on stairs or ladders in water transport injuring water skier
C0261260|ICD9CM|AB|E833.4|W/craft stair fall-skier
C0261261|ICD9CM|PT|E833.5|Fall on stairs or ladders in water transport injuring swimmer
C0261261|ICD9CM|AB|E833.5|W/craft stair fall-swim
C0261262|ICD9CM|PT|E833.6|Fall on stairs or ladders in water transport injuring dockers, stevedores
C0261262|ICD9CM|AB|E833.6|W/crf stair fall-docker
C0261263|ICD9CM|PT|E833.8|Fall on stairs or ladders in water transport injuring other specified person
C0261263|ICD9CM|AB|E833.8|W/crf stair fall-per NEC
C0261264|ICD9CM|PT|E833.9|Fall on stairs or ladders in water transport injuring unspecified person
C0261264|ICD9CM|AB|E833.9|W/crf stair fall-per NOS
C0261265|ICD9CM|HT|E834|Other fall from one level to another in water transport
C0261266|ICD9CM|PT|E834.0|Other fall from one level to another in water transport injuring occupant of small boat, unpowered
C0261266|ICD9CM|AB|E834.0|W/craft fall NEC-unpow
C0261267|ICD9CM|PT|E834.1|Other fall from one level to another in water transport injuring occupant of small boat, powered
C0261267|ICD9CM|AB|E834.1|W/craft fall NEC-power
C0261268|ICD9CM|PT|E834.2|Other fall from one level to another in water transport injuring occupant of other watercraft -- crew
C0261268|ICD9CM|AB|E834.2|Watercraft fall NEC-crew
C0261269|ICD9CM|PT|E834.3|Other fall from one level to another in water transport injuring occupant of other watercraft -- other than crew
C0261269|ICD9CM|AB|E834.3|Wtrcraft fall NEC-pasngr
C0261270|ICD9CM|PT|E834.4|Other fall from one level to another in water transport injuring water skier
C0261270|ICD9CM|AB|E834.4|W/craft fall NEC-skier
C0261271|ICD9CM|PT|E834.5|Other fall from one level to another in water transport injuring swimmer
C0261271|ICD9CM|AB|E834.5|W/craft fall NEC-swim
C0261272|ICD9CM|PT|E834.6|Other fall from one level to another in water transport injuring dockers, stevedores
C0261272|ICD9CM|AB|E834.6|Wtrcraft fall NEC-docker
C0261273|ICD9CM|PT|E834.8|Other fall from one level to another in water transport injuring other specified person
C0261273|ICD9CM|AB|E834.8|W/crft fall NEC-pers NEC
C0261274|ICD9CM|PT|E834.9|Other fall from one level to another in water transport injuring unspecified person
C0261274|ICD9CM|AB|E834.9|W/crft fall NEC-pers NOS
C0261275|ICD9CM|HT|E835|Other and unspecified fall in water transport
C0261276|ICD9CM|PT|E835.0|Other and unspecified fall in water transport injuring occupant of small boat, unpowered
C0261276|ICD9CM|AB|E835.0|W/craft fall NOS-unpow
C0261277|ICD9CM|PT|E835.1|Other and unspecified fall in water transport injuring occupant of small boat, powered
C0261277|ICD9CM|AB|E835.1|W/craft fall NOS-power
C0261278|ICD9CM|PT|E835.2|Other and unspecified fall in water transport injuring occupant of other watercraft -- crew
C0261278|ICD9CM|AB|E835.2|Wtrcraft fall NOS-crew
C0261279|ICD9CM|PT|E835.3|Other and unspecified fall in water transport injuring occupant of other watercraft -- other than crew
C0261279|ICD9CM|AB|E835.3|Wtrcraft fall NOS-pasngr
C0261280|ICD9CM|PT|E835.4|Other and unspecified fall in water transport injuring water skier
C0261280|ICD9CM|AB|E835.4|W/craft fall NOS-skier
C0261281|ICD9CM|PT|E835.5|Other and unspecified fall in water transport injuring swimmer
C0261281|ICD9CM|AB|E835.5|W/craft fall NOS-swim
C0261282|ICD9CM|PT|E835.6|Other and unspecified fall in water transport injuring dockers, stevedores
C0261282|ICD9CM|AB|E835.6|Wtrcraft fall NOS-docker
C0261283|ICD9CM|PT|E835.8|Other and unspecified fall in water transport injuring other specified person
C0261283|ICD9CM|AB|E835.8|W/crft fall NOS-pers NEC
C0261284|ICD9CM|PT|E835.9|Other and unspecified fall in water transport injuring unspecified person
C0261284|ICD9CM|AB|E835.9|W/crft fall NOS-pers NOS
C0261285|ICD9CM|HT|E836|Machinery accident in water transport
C0261286|ICD9CM|PT|E836.0|Machinery accident in water transport injuring occupant of small boat, unpowered
C0261286|ICD9CM|AB|E836.0|Machine acc-unpow boat
C0261287|ICD9CM|PT|E836.1|Machinery accident in water transport injuring occupant of small boat, powered
C0261287|ICD9CM|AB|E836.1|Mach acc-occ power boat
C0261288|ICD9CM|PT|E836.2|Machinery accident in water transport injuring occupant of other watercraft -- crew
C0261288|ICD9CM|AB|E836.2|Machinery accident-crew
C0261289|ICD9CM|PT|E836.3|Machinery accident in water transport injuring occupant of other watercraft -- other than crew
C0261289|ICD9CM|AB|E836.3|Machinery acc-pasngr
C0261290|ICD9CM|PT|E836.4|Machinery accident in water transport injuring water skier
C0261290|ICD9CM|AB|E836.4|Machine accident-skier
C0261291|ICD9CM|PT|E836.5|Machinery accident in water transport injuring swimmer
C0261291|ICD9CM|AB|E836.5|Machine accident-swim
C0261292|ICD9CM|PT|E836.6|Machinery accident in water transport injuring dockers, stevedores
C0261292|ICD9CM|AB|E836.6|Machinery acc-docker
C0261293|ICD9CM|PT|E836.8|Machinery accident in water transport injuring other specified person
C0261293|ICD9CM|AB|E836.8|Machinery acc-pers NEC
C0261294|ICD9CM|PT|E836.9|Machinery accident in water transport injuring unspecified person
C0261294|ICD9CM|AB|E836.9|Machinery acc-pers NOS
C0261295|ICD9CM|HT|E837|Explosion, fire, or burning in watercraft
C0261296|ICD9CM|PT|E837.0|Explosion, fire, or burning in watercraft injuring occupant of small boat, unpowered
C0261296|ICD9CM|AB|E837.0|Explosion-occ unpow boat
C0261297|ICD9CM|PT|E837.1|Explosion, fire, or burning in watercraft injuring occupant of small boat, powered
C0261297|ICD9CM|AB|E837.1|Explosion-occ power boat
C0261298|ICD9CM|PT|E837.2|Explosion, fire, or burning in watercraft injuring occupant of other watercraft -- crew
C0261298|ICD9CM|AB|E837.2|Watercraft explos-crew
C0261299|ICD9CM|PT|E837.3|Explosion, fire, or burning in watercraft injuring occupant of other watercraft -- other than crew
C0261299|ICD9CM|AB|E837.3|Watercraft explos-pasngr
C0261300|ICD9CM|PT|E837.4|Explosion, fire, or burning in watercraft injuring water skier
C0261300|ICD9CM|AB|E837.4|Watercraft explos-skier
C0261301|ICD9CM|PT|E837.5|Explosion, fire, or burning in watercraft injuring swimmer
C0261301|ICD9CM|AB|E837.5|Watercraft explos-swim
C0261302|ICD9CM|PT|E837.6|Explosion, fire, or burning in watercraft injuring dockers, stevedores
C0261302|ICD9CM|AB|E837.6|Watercraft explos-docker
C0261303|ICD9CM|PT|E837.8|Explosion, fire, or burning in watercraft injuring other specified person
C0261303|ICD9CM|AB|E837.8|Watercraft expl-pers NEC
C0261304|ICD9CM|PT|E837.9|Explosion, fire, or burning in watercraft injuring unspecified person
C0261304|ICD9CM|AB|E837.9|Watercraft expl-pers NOS
C0261306|ICD9CM|PT|E838.0|Other and unspecified water transport accident injuring occupant of small boat, unpowered
C0261306|ICD9CM|AB|E838.0|Watercraft acc NEC-unpow
C0261307|ICD9CM|PT|E838.1|Other and unspecified water transport accident injuring occupant of small boat, powered
C0261307|ICD9CM|AB|E838.1|Watercraft acc NEC-power
C0261308|ICD9CM|PT|E838.2|Other and unspecified water transport accident injuring occupant of other watercraft -- crew
C0261308|ICD9CM|AB|E838.2|Watercraft acc NEC-crew
C0261309|ICD9CM|PT|E838.3|Other and unspecified water transport accident injuring occupant of other watercraft -- other than crew
C0261309|ICD9CM|AB|E838.3|Watercrft acc NEC-pasngr
C0261310|ICD9CM|PT|E838.4|Other and unspecified water transport accident injuring water skier
C0261310|ICD9CM|AB|E838.4|Watercraft acc NEC-skier
C0261311|ICD9CM|PT|E838.5|Other and unspecified water transport accident injuring swimmer
C0261311|ICD9CM|AB|E838.5|Watrcrft acc NEC-swimmer
C0261312|ICD9CM|PT|E838.6|Other and unspecified water transport accident injuring dockers, stevedores
C0261312|ICD9CM|AB|E838.6|Watercrft acc NEC-docker
C0261313|ICD9CM|PT|E838.8|Other and unspecified water transport accident injuring other specified person
C0261313|ICD9CM|AB|E838.8|Wtrcrft acc NEC-pers NEC
C0261314|ICD9CM|PT|E838.9|Other and unspecified water transport accident injuring unspecified person
C0261314|ICD9CM|HT|E838|Other and unspecified water transport accident
C0261314|ICD9CM|AB|E838.9|Wtrcrft acc NEC-pers NOS
C0261315|ICD9CM|HT|E840|Accident to powered aircraft at takeoff or landing
C0261316|ICD9CM|PT|E840.0|Accident to powered aircraft at takeoff or landing injuring occupant of spacecraft
C0261316|ICD9CM|AB|E840.0|Tk off/land-spcrft
C0261317|ICD9CM|PT|E840.1|Accident to powered aircraft at takeoff or landing injuring occupant of military aircraft, any
C0261317|ICD9CM|AB|E840.1|Tk off/land-milit craft
C0261318|ICD9CM|PT|E840.2|Accident to powered aircraft at takeoff or landing injuring crew of commercial aircraft (powered) in surface to surface transport
C0261318|ICD9CM|AB|E840.2|Tk off/land-crew aircrft
C0261319|ICD9CM|PT|E840.3|Accident to powered aircraft at takeoff or landing injuring other occupant of commercial aircraft (powered) in surface to surface transport
C0261319|ICD9CM|AB|E840.3|Tk off/land-psng aircrft
C0261320|ICD9CM|PT|E840.4|Accident to powered aircraft at takeoff or landing injuring occupant of commercial aircraft (powered) in surface to air transport
C0261320|ICD9CM|AB|E840.4|Tk off/land-comm crf NEC
C0261321|ICD9CM|PT|E840.5|Accident to powered aircraft at takeoff or landing injuring occupant of other powered aircraft
C0261321|ICD9CM|AB|E840.5|Tk off/land-aircraft NEC
C0261322|ICD9CM|PT|E840.6|Accident to powered aircraft at takeoff or landing injuring occupant of unpowered aircraft, except parachutist
C0261322|ICD9CM|AB|E840.6|Tk off/land-unp aircrft
C0261323|ICD9CM|PT|E840.7|Accident to powered aircraft at takeoff or landing injuring parachutist (military) (other)
C0261323|ICD9CM|AB|E840.7|Tk off/land-parachutist
C0261324|ICD9CM|PT|E840.8|Accident to powered aircraft at takeoff or landing injuring ground crew, airline employee
C0261324|ICD9CM|AB|E840.8|Tk off/land-ground crew
C0261325|ICD9CM|PT|E840.9|Accident to powered aircraft at takeoff or landing injuring other person
C0261325|ICD9CM|AB|E840.9|Tk off/land-pers NEC
C0261327|ICD9CM|PT|E841.0|Accident to powered aircraft, other and unspecified, injuring occupant of spacecraft
C0261327|ICD9CM|AB|E841.0|Pow aircraft acc-spcrft
C0261328|ICD9CM|PT|E841.1|Accident to powered aircraft, other and unspecified, injuring occupant of military aircraft, any
C0261328|ICD9CM|AB|E841.1|Power aircraft acc-milit
C0261329|ICD9CM|PT|E841.2|Accident to powered aircraft, other and unspecified, injuring crew of commercial aircraft (powered) in surface to surface transport
C0261329|ICD9CM|AB|E841.2|Power aircraft acc-crew
C0261330|ICD9CM|PT|E841.3|Accident to powered aircraft, other and unspecified, injuring other occupant of commercial aircraft (powered) in surface to surface transport
C0261330|ICD9CM|AB|E841.3|Power aircraft acc-psngr
C0261331|ICD9CM|PT|E841.4|Accident to powered aircraft, other and unspecified, injuring occupant of commercial aircraft (powered) in surface to air transport
C0261331|ICD9CM|AB|E841.4|Aircraf acc-occ comm NEC
C0261332|ICD9CM|PT|E841.5|Accident to powered aircraft, other and unspecified, injuring occupant of other powered aircraft
C0261332|ICD9CM|AB|E841.5|Oth powered aircraft acc
C0261333|ICD9CM|PT|E841.6|Accident to powered aircraft, other and unspecified, injuring occupant of unpowered aircraft, except parachutist
C0261333|ICD9CM|AB|E841.6|Pow airc acc-unp aircr
C0261334|ICD9CM|PT|E841.7|Accident to powered aircraft, other and unspecified, injuring parachutist (military) (other)
C0261334|ICD9CM|AB|E841.7|Aircraft acc-parachutist
C0261335|ICD9CM|PT|E841.8|Accident to powered aircraft, other and unspecified, injuring ground crew, airline employee
C0261335|ICD9CM|AB|E841.8|Aircraft acc-ground crew
C0261336|ICD9CM|PT|E841.9|Accident to powered aircraft, other and unspecified, injuring other person
C0261336|ICD9CM|AB|E841.9|Aircrft acc NOS-pers NEC
C0261337|ICD9CM|HT|E842|Accident to unpowered aircraft
C0261338|ICD9CM|PT|E842.6|Accident to unpowered aircraft injuring occupant of unpowered aircraft, except parachutist
C0261338|ICD9CM|AB|E842.6|Unpower aircraft acc-occ
C0261340|ICD9CM|PT|E842.8|Accident to unpowered aircraft injuring ground crew, airline employee
C0261340|ICD9CM|AB|E842.8|Unpow aircrf acc-gr crew
C0261341|ICD9CM|PT|E842.9|Accident to unpowered aircraft injuring other person
C0261341|ICD9CM|AB|E842.9|Unpow aircrf acc-per NEC
C0261342|ICD9CM|HT|E843|Fall in, on, or from aircraft
C0261343|ICD9CM|PT|E843.0|Fall in, on, or from aircraft injuring occupant of spacecraft
C0261343|ICD9CM|AB|E843.0|Fall-occ spacecraft
C0261344|ICD9CM|PT|E843.1|Fall in, on, or from aircraft injuring occupant of military aircraft, any
C0261344|ICD9CM|AB|E843.1|Fall-milit aircraft occp
C0261345|ICD9CM|PT|E843.2|Fall in, on, or from aircraft injuring crew of commercial aircraft (powered) in surface to surface transport
C0261345|ICD9CM|AB|E843.2|Fall-crew comm aircraft
C0261346|ICD9CM|PT|E843.3|Fall in, on, or from aircraft injuring other occupant of commercial aircraft (powered) in surface to surface transport
C0261346|ICD9CM|AB|E843.3|Fall-psng comm aircraft
C0261347|ICD9CM|PT|E843.4|Fall in, on, or from aircraft injuring occupant of commercial aircraft (powered) in surface to air transport
C0261347|ICD9CM|AB|E843.4|Fall-occ comm aircrf NEC
C0261348|ICD9CM|PT|E843.5|Fall in, on, or from aircraft injuring occupant of other powered aircraft
C0261348|ICD9CM|AB|E843.5|Fall-occup oth aircraft
C0261349|ICD9CM|PT|E843.6|Fall in, on, or from aircraft injuring occupant of unpowered aircraft, except parachutist
C0261349|ICD9CM|AB|E843.6|Fall-occ unpower aircraf
C0261350|ICD9CM|PT|E843.7|Fall in, on, or from aircraft injuring parachutist (military) (other)
C0261350|ICD9CM|AB|E843.7|Fall-parachutist
C0261351|ICD9CM|PT|E843.8|Fall in, on, or from aircraft injuring ground crew, airline employee
C0261351|ICD9CM|AB|E843.8|Aircrft fall-ground crew
C0261352|ICD9CM|PT|E843.9|Fall in, on, or from aircraft injuring other person
C0261352|ICD9CM|AB|E843.9|Aircraft fall-person NEC
C0261353|ICD9CM|HT|E844|Other specified air transport accidents
C0261354|ICD9CM|PT|E844.0|Other specified air transport accidents injuring occupant of spacecraft
C0261354|ICD9CM|AB|E844.0|Aircrft acc NEC-spcrft
C0261355|ICD9CM|PT|E844.1|Other specified air transport accidents injuring occupant of military aircraft, any
C0261355|ICD9CM|AB|E844.1|Aircrft acc NEC-military
C0261356|ICD9CM|PT|E844.2|Other specified air transport accidents injuring crew of commercial aircraft (powered) in surface to surface transport
C0261356|ICD9CM|AB|E844.2|Aircrft acc NEC-crew
C0261357|ICD9CM|PT|E844.3|Other specified air transport accidents injuring other occupant of commercial aircraft (powered) in surface to surface transport
C0261357|ICD9CM|AB|E844.3|Aircrft acc NEC-pasngr
C0261358|ICD9CM|PT|E844.4|Other specified air transport accidents injuring occupant of commercial aircraft (powered) in surface to air transport
C0261358|ICD9CM|AB|E844.4|Aircrft acc NEC-comm NEC
C0261359|ICD9CM|PT|E844.5|Other specified air transport accidents injuring occupant of other powered aircraft
C0261359|ICD9CM|AB|E844.5|Aircrft acc NEC-occp NEC
C0261360|ICD9CM|PT|E844.6|Other specified air transport accidents injuring occupant of unpowered aircraft, except parachutist
C0261360|ICD9CM|AB|E844.6|Aircr acc NEC-unp aircr
C0261361|ICD9CM|PT|E844.7|Other specified air transport accidents injuring parachutist (military) (other)
C0261361|ICD9CM|AB|E844.7|Aircrft acc-parachutist
C0261362|ICD9CM|PT|E844.8|Other specified air transport accidents injuring ground crew, airline employee
C0261362|ICD9CM|AB|E844.8|Aircrft acc NEC-grd crew
C0261363|ICD9CM|PT|E844.9|Other specified air transport accidents injuring other person
C0261363|ICD9CM|AB|E844.9|Aircrft acc NEC-pers NEC
C0261364|ICD9CM|HT|E845|Accident involving spacecraft
C0261365|ICD9CM|PT|E845.0|Accident involving spacecraft injuring occupant of spacecraft
C0261365|ICD9CM|AB|E845.0|Spacecraft acc-occupant
C0261366|ICD9CM|PT|E845.8|Accident involving spacecraft injuring ground crew, airline employee
C0261366|ICD9CM|AB|E845.8|Spacecraft acc-grnd crew
C0261367|ICD9CM|PT|E845.9|Accident involving spacecraft injuring other person
C0261367|ICD9CM|AB|E845.9|Spacecraft acc-pers NEC
C0261368|ICD9CM|PT|E846|Accidents involving powered vehicles used solely within the buildings and premises of industrial or commercial establishment
C0261368|ICD9CM|AB|E846|Indus veh acc on premise
C0261369|ICD9CM|PT|E847|Accidents involving cable cars not running on rails
C0261369|ICD9CM|AB|E847|Cabl car acc not on rail
C0261370|ICD9CM|PT|E848|Accidents involving other vehicles, not elsewhere classifiable
C0261370|ICD9CM|AB|E848|Oth vehicle acc NEC
C0261371|ICD9CM|HT|E849-E849.9|PLACE OF OCCURRENCE
C0261372|ICD9CM|PT|E849.1|Farm accidents
C0261372|ICD9CM|AB|E849.1|Accident on farm
C0261373|ICD9CM|PT|E849.2|Mine and quarry accidents
C0261373|ICD9CM|AB|E849.2|Accident in mine/quarry
C0261374|ICD9CM|PT|E849.3|Accidents occurring in industrial places and premises
C0261374|ICD9CM|AB|E849.3|Acc on industr premises
C0261375|ICD9CM|PT|E849.4|Accidents occurring in place for recreation and sport
C0261375|ICD9CM|AB|E849.4|Accid in recreation area
C0261376|ICD9CM|PT|E849.5|Street and highway accidents
C0261376|ICD9CM|AB|E849.5|Accid on street/highway
C0261377|ICD9CM|PT|E849.6|Accidents occurring in public building
C0261377|ICD9CM|AB|E849.6|Accident in public bldg
C0261378|ICD9CM|PT|E849.7|Accidents occurring in residential institution
C0261378|ICD9CM|AB|E849.7|Accid in resident instit
C0261379|ICD9CM|PT|E849.8|Accidents occurring in other specified places
C0261379|ICD9CM|AB|E849.8|Accident in place NEC
C0261380|ICD9CM|PT|E849.9|Accidents occurring in unspecified place
C0261380|ICD9CM|AB|E849.9|Accident in place NOS
C0261381|ICD9CM|HT|E850|Accidental poisoning by analgesics, antipyretics, and antirheumatics
C0261382|ICD9CM|PT|E850.0|Accidental poisoning by heroin
C0261382|ICD9CM|AB|E850.0|Acc poison-heroin
C0261383|ICD9CM|PT|E850.1|Accidental poisoning by methadone
C0261383|ICD9CM|AB|E850.1|Acc poison-methadone
C0261384|ICD9CM|PT|E850.2|Accidental poisoning by other opiates and related narcotics
C0261384|ICD9CM|AB|E850.2|Acc poison-opiates NEC
C0261385|ICD9CM|PT|E850.3|Accidental poisoning by salicylates
C0261385|ICD9CM|AB|E850.3|Acc poison-salicylates
C0261387|ICD9CM|PT|E850.5|Accidental poisoning by pyrazole derivatives
C0261387|ICD9CM|AB|E850.5|Acc poison-pyrazole derv
C0261389|ICD9CM|PT|E850.7|Accidental poisoning by other non-narcotic analgesics
C0261389|ICD9CM|AB|E850.7|Acc poison-nonnarc analg
C0261390|ICD9CM|PT|E850.8|Accidental poisoning by other specified analgesics and antipyretics
C0261390|ICD9CM|AB|E850.8|Acc poison-analgesic NEC
C0261391|ICD9CM|PT|E850.9|Accidental poisoning by unspecified analgesic or antipyretic
C0261391|ICD9CM|AB|E850.9|Acc poison-analgesic NOS
C0261392|ICD9CM|PT|E851|Accidental poisoning by barbiturates
C0261392|ICD9CM|AB|E851|Acc poison-barbiturates
C0261393|ICD9CM|HT|E852|Accidental poisoning by other sedatives and hypnotics
C0261394|ICD9CM|PT|E852.0|Accidental poisoning by chloral hydrate group
C0261394|ICD9CM|AB|E852.0|Acc poisn-chlorl hydrate
C0261395|ICD9CM|PT|E852.1|Accidental poisoning by paraldehyde
C0261395|ICD9CM|AB|E852.1|Acc poison-paraldehyde
C0261396|ICD9CM|PT|E852.2|Accidental poisoning by bromine compounds
C0261396|ICD9CM|AB|E852.2|Acc poison-bromine cmpnd
C0261397|ICD9CM|PT|E852.3|Accidental poisoning by methaqualone compounds
C0261397|ICD9CM|AB|E852.3|Acc poison-methaqualone
C0261398|ICD9CM|PT|E852.4|Accidental poisoning by glutethimide group
C0261398|ICD9CM|AB|E852.4|Acc poison-glutethimide
C0261400|ICD9CM|PT|E852.8|Accidental poisoning by other specified sedatives and hypnotics
C0261400|ICD9CM|AB|E852.8|Acc poison-sedatives NEC
C0261401|ICD9CM|PT|E852.9|Accidental poisoning by unspecified sedative or hypnotic
C0261401|ICD9CM|AB|E852.9|Acc poison-sedatives NOS
C0261402|ICD9CM|HT|E853|Accidental poisoning by tranquilizers
C0261403|ICD9CM|PT|E853.0|Accidental poisoning by phenothiazine-based tranquilizers
C0261403|ICD9CM|AB|E853.0|Acc pois-phenthiaz tranq
C0261404|ICD9CM|PT|E853.1|Accidental poisoning by butyrophenone-based tranquilizers
C0261404|ICD9CM|AB|E853.1|Acc pois-butyrphen tranq
C0261405|ICD9CM|PT|E853.2|Accidental poisoning by benzodiazepine-based tranquilizers
C0261405|ICD9CM|AB|E853.2|Acc poisn-benzdiaz tranq
C0261406|ICD9CM|PT|E853.8|Accidental poisoning by other specified tranquilizers
C0261406|ICD9CM|AB|E853.8|Acc poisn-tranquilzr NEC
C0261407|ICD9CM|PT|E853.9|Accidental poisoning by unspecified tranquilizer
C0261407|ICD9CM|AB|E853.9|Acc poisn-tranquilzr NOS
C0261408|ICD9CM|HT|E854|Accidental poisoning by other psychotropic agents
C0261408|ICD9CM|PT|E854.8|Accidental poisoning by other psychotropic agents
C0261408|ICD9CM|AB|E854.8|Acc poisn psychotrop NEC
C0261409|ICD9CM|PT|E854.0|Accidental poisoning by antidepressants
C0261409|ICD9CM|AB|E854.0|Acc poison-antidepressnt
C0261411|ICD9CM|PT|E854.2|Accidental poisoning by psychostimulants
C0261411|ICD9CM|AB|E854.2|Acc poisn-psychstimulant
C0261412|ICD9CM|PT|E854.3|Accidental poisoning by central nervous system stimulants
C0261412|ICD9CM|AB|E854.3|Acc poison-cns stimulant
C0261413|ICD9CM|HT|E855|Accidental poisoning by other drugs acting on central and autonomic nervous system
C0261414|ICD9CM|PT|E855.0|Accidental poisoning by anticonvulsant and anti-parkinsonism drugs
C0261414|ICD9CM|AB|E855.0|Acc poisn-anticonvulsant
C0261415|ICD9CM|PT|E855.1|Accidental poisoning by other central nervous system depressants
C0261415|ICD9CM|AB|E855.1|Acc poisn-cns depres NEC
C0261416|ICD9CM|PT|E855.2|Accidental poisoning by local anesthetics
C0261416|ICD9CM|AB|E855.2|Acc poisn-local anesthet
C0261418|ICD9CM|PT|E855.4|Accidental poisoning by parasympatholytics [anticholinergics and antimuscarinics] and spasmolytics
C0261418|ICD9CM|AB|E855.4|Acc poisn-anticholinerg
C0261421|ICD9CM|PT|E855.8|Accidental poisoning by other specified drugs acting on central and autonomic nervous systems
C0261421|ICD9CM|AB|E855.8|Acc poison-cns drug NEC
C0261422|ICD9CM|PT|E855.9|Accidental poisoning by unspecified drug acting on central and autonomic nervous systems
C0261422|ICD9CM|AB|E855.9|Acc poison-cns drug NOS
C0261423|ICD9CM|PT|E856|Accidental poisoning by antibiotics
C0261423|ICD9CM|AB|E856|Acc poison-antibiotics
C0261424|ICD9CM|PT|E857|Accidental poisoning by other anti-infectives
C0261424|ICD9CM|AB|E857|Acc pois-oth anti-infect
C0261425|ICD9CM|HT|E858|Accidental poisoning by other drugs
C0261426|ICD9CM|PT|E858.0|Accidental poisoning by hormones and synthetic substitutes
C0261426|ICD9CM|AB|E858.0|Acc poison-hormones
C0261427|ICD9CM|PT|E858.1|Accidental poisoning by primarily systemic agents
C0261427|ICD9CM|AB|E858.1|Acc poisn-systemic agent
C0261428|ICD9CM|PT|E858.2|Accidental poisoning by agents primarily affecting blood constituents
C0261428|ICD9CM|AB|E858.2|Acc poison-blood agent
C0261429|ICD9CM|PT|E858.3|Accidental poisoning by agents primarily affecting cardiovascular system
C0261429|ICD9CM|AB|E858.3|Acc poisn-cardiovasc agt
C0261430|ICD9CM|PT|E858.4|Accidental poisoning by agents primarily affecting gastrointestinal system
C0261430|ICD9CM|AB|E858.4|Acc poison-gi agent
C0261431|ICD9CM|PT|E858.5|Accidental poisoning by water, mineral, and uric acid metabolism drugs
C0261431|ICD9CM|AB|E858.5|Acc poisn-metabol agnt
C0261432|ICD9CM|PT|E858.6|Accidental poisoning by agents primarily acting on the smooth and skeletal muscles and respiratory system
C0261432|ICD9CM|AB|E858.6|Acc poisn-muscl/resp agt
C0261434|ICD9CM|PT|E858.8|Accidental poisoning by other specified drugs
C0261434|ICD9CM|AB|E858.8|Acc poisoning-drug NEC
C0261435|ICD9CM|PT|E858.9|Accidental poisoning by unspecified drug
C0261435|ICD9CM|AB|E858.9|Acc poisoning-drug NOS
C0261437|ICD9CM|PT|E860.0|Accidental poisoning by alcoholic beverages
C0261437|ICD9CM|AB|E860.0|Acc poisn-alcohol bevrag
C0261438|ICD9CM|PT|E860.1|Accidental poisoning by other and unspecified ethyl alcohol and its products
C0261438|ICD9CM|AB|E860.1|Acc poison-ethyl alcohol
C0261439|ICD9CM|PT|E860.2|Accidental poisoning by methyl alcohol
C0261439|ICD9CM|AB|E860.2|Acc poisn-methyl alcohol
C0261440|ICD9CM|PT|E860.3|Accidental poisoning by isopropyl alcohol
C0261440|ICD9CM|AB|E860.3|Acc poisn-isopropyl alc
C0261441|ICD9CM|PT|E860.4|Accidental poisoning by fusel oil
C0261441|ICD9CM|AB|E860.4|Acc poison-fusel oil
C0261442|ICD9CM|PT|E860.8|Accidental poisoning by other specified alcohols
C0261442|ICD9CM|AB|E860.8|Acc poison-alcohol NEC
C0261444|ICD9CM|HT|E861|Accidental poisoning by cleansing and polishing agents, disinfectants, paints, and varnishes
C0261445|ICD9CM|PT|E861.0|Accidental poisoning by synthetic detergents and shampoos
C0261445|ICD9CM|AB|E861.0|Acc pois-synth detergent
C0261446|ICD9CM|PT|E861.1|Accidental poisoning by soap products
C0261446|ICD9CM|AB|E861.1|Acc poison-soap products
C0261447|ICD9CM|PT|E861.2|Accidental poisoning by polishes
C0261447|ICD9CM|AB|E861.2|Acc poison-polishes
C0261449|ICD9CM|PT|E861.4|Accidental poisoning by disinfectants
C0261449|ICD9CM|AB|E861.4|Acc poison-disinfectants
C0261450|ICD9CM|PT|E861.5|Accidental poisoning by lead paints
C0261450|ICD9CM|AB|E861.5|Acc poison-lead paints
C0261451|ICD9CM|PT|E861.6|Accidental poisoning by other paints and varnishes
C0261451|ICD9CM|AB|E861.6|Acc poison-paints NEC
C0261452|ICD9CM|PT|E861.9|Accidental poisoning by unspecified cleansing and polishing agents, disinfectants, paints, and varnishes
C0261452|ICD9CM|AB|E861.9|Acc poison-cleanser NOS
C0261454|ICD9CM|PT|E862.0|Accidental poisoning by petroleum solvents
C0261454|ICD9CM|AB|E862.0|Acc poisn-petrol solvent
C0261456|ICD9CM|PT|E862.2|Accidental poisoning by lubricating oils
C0261456|ICD9CM|AB|E862.2|Acc pois-lubricating oil
C0261457|ICD9CM|PT|E862.3|Accidental poisoning by petroleum solids
C0261457|ICD9CM|AB|E862.3|Acc pois-petroleum solid
C0261460|ICD9CM|HT|E863|Accidental poisoning by agricultural and horticultural chemical and pharmaceutical preparations other than plant foods and fertilizers
C0261461|ICD9CM|PT|E863.0|Accidental poisoning by insecticides of organochlorine compounds
C0261461|ICD9CM|AB|E863.0|Acc pois-chlorine pestic
C0261462|ICD9CM|PT|E863.1|Accidental poisoning by insecticides of organophosphorus compounds
C0261462|ICD9CM|AB|E863.1|Acc pois-phosph pesticid
C0261463|ICD9CM|PT|E863.2|Accidental poisoning by carbamates
C0261463|ICD9CM|AB|E863.2|Acc poison-carbamates
C0261464|ICD9CM|PT|E863.3|Accidental poisoning by mixtures of insecticides
C0261464|ICD9CM|AB|E863.3|Acc poisn-mixed pesticid
C0261465|ICD9CM|PT|E863.4|Accidental poisoning by other and unspecified insecticides
C0261465|ICD9CM|AB|E863.4|Acc poison-pesticide NEC
C0261466|ICD9CM|PT|E863.5|Accidental poisoning by herbicides
C0261466|ICD9CM|AB|E863.5|Acc poison-herbicides
C0261467|ICD9CM|PT|E863.6|Accidental poisoning by fungicides
C0261467|ICD9CM|AB|E863.6|Acc poison-fungicides
C0261468|ICD9CM|PT|E863.7|Accidental poisoning by rodenticides
C0261468|ICD9CM|AB|E863.7|Acc poison-rodenticides
C0261469|ICD9CM|PT|E863.8|Accidental poisoning by fumigants
C0261469|ICD9CM|AB|E863.8|Acc poison-fumigants
C0261470|ICD9CM|PT|E863.9|Accidental poisoning by other and unspecified agricultural and horticultural chemical and pharmaceutical preparations other than plant foods and fertilizers
C0261470|ICD9CM|AB|E863.9|Acc pois-agrcult NEC/NOS
C0261479|ICD9CM|PT|E865.1|Accidental poisoning by shellfish
C0261479|ICD9CM|AB|E865.1|Acc poison-shellfish
C0261481|ICD9CM|PT|E865.4|Accidental poisoning from other specified plants
C0261481|ICD9CM|AB|E865.4|Acc poison-plants NEC
C0261482|ICD9CM|PT|E865.5|Accidental poisoning from mushrooms and other fungi
C0261482|ICD9CM|AB|E865.5|Acc poison-mushrooms
C0261483|ICD9CM|PT|E865.8|Accidental poisoning from other specified foods
C0261483|ICD9CM|AB|E865.8|Acc poison-food NEC
C0261484|ICD9CM|PT|E865.9|Accidental poisoning from unspecified foodstuff or poisonous plant
C0261484|ICD9CM|AB|E865.9|Acc poisn-food/plant NOS
C0261485|ICD9CM|HT|E866|Accidental poisoning by other and unspecified solid and liquid substances
C0261486|ICD9CM|PT|E866.0|Accidental poisoning by lead and its compounds and fumes
C0261486|ICD9CM|AB|E866.0|Acc poisoning-lead
C0261487|ICD9CM|PT|E866.1|Accidental poisoning by mercury and its compounds and fumes
C0261487|ICD9CM|AB|E866.1|Acc poisoning-mercury
C0261488|ICD9CM|PT|E866.2|Accidental poisoning by antimony and its compounds and fumes
C0261488|ICD9CM|AB|E866.2|Acc poisoning-antimony
C0261489|ICD9CM|PT|E866.3|Accidental poisoning by arsenic and its compounds and fumes
C0261489|ICD9CM|AB|E866.3|Acc poisoning-arsenic
C0261490|ICD9CM|PT|E866.4|Accidental poisoning by other metals and their compounds and fumes
C0261490|ICD9CM|AB|E866.4|Acc poison-metals NEC
C0261491|ICD9CM|PT|E866.5|Accidental poisoning by plant foods and fertilizers
C0261491|ICD9CM|AB|E866.5|Acc poison-plant food
C0261492|ICD9CM|PT|E866.6|Accidental poisoning by glues and adhesives
C0261492|ICD9CM|AB|E866.6|Acc poison-glues
C0261493|ICD9CM|PT|E866.7|Accidental poisoning by cosmetics
C0261493|ICD9CM|AB|E866.7|Acc poison-cosmetics
C0261494|ICD9CM|PT|E866.8|Accidental poisoning by other specified solid or liquid substances
C0261494|ICD9CM|AB|E866.8|Acc pois-solid/liq NEC
C0261495|ICD9CM|PT|E866.9|Accidental poisoning by unspecified solid or liquid substance
C0261495|ICD9CM|AB|E866.9|Acc pois-solid/liq NOS
C0261496|ICD9CM|PT|E867|Accidental poisoning by gas distributed by pipeline
C0261496|ICD9CM|AB|E867|Acc poison-piped gas
C0261497|ICD9CM|HT|E868|Accidental poisoning by other utility gas and other carbon monoxide
C0261498|ICD9CM|PT|E868.0|Accidental poisoning by liquefied petroleum gas distributed in mobile containers
C0261498|ICD9CM|AB|E868.0|Acc pois-liq petrol gas
C0261499|ICD9CM|PT|E868.1|Accidental poisoning by other and unspecified utility gas
C0261499|ICD9CM|AB|E868.1|Acc pois-utl gas NEC/NOS
C0261500|ICD9CM|PT|E868.2|Accidental poisoning by motor vehicle exhaust gas
C0261500|ICD9CM|AB|E868.2|Acc poison-exhaust gas
C0261501|ICD9CM|PT|E868.3|Accidental poisoning by carbon monoxide from incomplete combustion of other domestic fuels
C0261501|ICD9CM|AB|E868.3|Acc pois-co/domestc fuel
C0261502|ICD9CM|PT|E868.8|Accidental poisoning by carbon monoxide from other sources
C0261502|ICD9CM|AB|E868.8|Acc pois-carbn monox NEC
C0261503|ICD9CM|PT|E868.9|Accidental poisoning by unspecified carbon monoxide
C0261503|ICD9CM|AB|E868.9|Acc pois-carbn monox NOS
C0261504|ICD9CM|HT|E869|Accidental poisoning by other gases and vapors
C0261505|ICD9CM|PT|E869.0|Accidental poisoning by nitrogen oxides
C0261505|ICD9CM|AB|E869.0|Acc poisn-nitrogen oxide
C0261506|ICD9CM|PT|E869.1|Accidental poisoning by sulfur dioxide
C0261506|ICD9CM|AB|E869.1|Acc poisn-sulfur dioxide
C0261507|ICD9CM|PT|E869.2|Accidental poisoning by freon
C0261507|ICD9CM|AB|E869.2|Acc poison-freon
C0261509|ICD9CM|PT|E869.8|Accidental poisoning by other specified gases and vapors
C0261509|ICD9CM|AB|E869.8|Acc poison-gas/vapor NEC
C0261510|ICD9CM|PT|E869.9|Accidental poisoning by unspecified gases and vapors
C0261510|ICD9CM|AB|E869.9|Acc poison-gas/vapor NOS
C0261513|ICD9CM|HT|E870|Accidental cut, puncture, perforation, or hemorrhage during medical care
C0261513|ICD9CM|PT|E870.9|Accidental cut, puncture, perforation or hemorrhage during unspecified medical care
C0261513|ICD9CM|AB|E870.9|Acc cut in med care NOS
C0261514|ICD9CM|PT|E870.2|Accidental cut, puncture, perforation or hemorrhage during kidney dialysis or other perfusion
C0261514|ICD9CM|AB|E870.2|Acc cut/hem-perfusn NEC
C0261515|ICD9CM|PT|E870.3|Accidental cut, puncture, perforation or hemorrhage during injection or vaccination
C0261515|ICD9CM|AB|E870.3|Acc cut/hem in injection
C0261516|ICD9CM|PT|E870.4|Accidental cut, puncture, perforation or hemorrhage during endoscopic examination
C0261516|ICD9CM|AB|E870.4|Acc cut/hem w scope exam
C0261517|ICD9CM|PT|E870.5|Accidental cut, puncture, perforation or hemorrhage during aspiration of fluid or tissue, puncture, and catheterization
C0261517|ICD9CM|AB|E870.5|Acc cut/hem w catheteriz
C0261518|ICD9CM|PT|E870.6|Accidental cut, puncture, perforation or hemorrhage during heart catheterization
C0261518|ICD9CM|AB|E870.6|Acc cut/hem w heart cath
C0261519|ICD9CM|PT|E870.7|Accidental cut, puncture, perforation or hemorrhage during administration of enema
C0261519|ICD9CM|AB|E870.7|Acc cut/hem w enema
C0261520|ICD9CM|PT|E870.8|Accidental cut, puncture, perforation or hemorrhage during other specified medical care
C0261520|ICD9CM|AB|E870.8|Acc cut in med care NEC
C0261522|ICD9CM|HT|E871|Foreign object left in body during procedure
C0261531|ICD9CM|PT|E871.8|Foreign object left in body during other specified procedures
C0261531|ICD9CM|AB|E871.8|Post-op foreign body NEC
C0261532|ICD9CM|PT|E871.9|Foreign object left in body during unspecified procedure
C0261532|ICD9CM|AB|E871.9|Post-op foreign body NOS
C0261533|ICD9CM|PT|E872.0|Failure of sterile precautions during surgical operation
C0261533|ICD9CM|HT|E872|Failure of sterile precautions during procedure
C0261533|ICD9CM|AB|E872.0|Failure sterile surgery
C0261536|ICD9CM|PT|E872.2|Failure of sterile precautions during kidney dialysis and other perfusion
C0261536|ICD9CM|AB|E872.2|Fail sterile perfusn NEC
C0261539|ICD9CM|PT|E872.5|Failure of sterile precautions during aspiration of fluid or tissue, puncture, and catheterization
C0261539|ICD9CM|AB|E872.5|Fail sterile catheter
C0261541|ICD9CM|PT|E872.8|Failure of sterile precautions during other specified procedures
C0261541|ICD9CM|AB|E872.8|Fail sterile proced NEC
C0261542|ICD9CM|PT|E872.9|Failure of sterile precautions during unspecified procedure
C0261542|ICD9CM|AB|E872.9|Fail sterile proced NOS
C0261543|ICD9CM|HT|E873|Failure in dosage
C0261543|ICD9CM|AB|E873.9|Failure in dosage NOS
C0261543|ICD9CM|PT|E873.9|Unspecified failure in dosage
C0261547|ICD9CM|PT|E873.3|Inadvertent exposure of patient to radiation during medical care
C0261547|ICD9CM|AB|E873.3|Inadv radiat exp-medical
C0261548|ICD9CM|PT|E873.4|Failure in dosage in electroshock or insulin-shock therapy
C0261548|ICD9CM|AB|E873.4|Dosag fail-shock therapy
C0261551|ICD9CM|PT|E873.8|Other specified failure in dosage
C0261551|ICD9CM|AB|E873.8|Failure in dosage NEC
C0261553|ICD9CM|HT|E874|Mechanical failure of instrument or apparatus during procedure
C0261554|ICD9CM|PT|E874.0|Mechanical failure of instrument or apparatus during surgical operation
C0261554|ICD9CM|AB|E874.0|Instrmnt fail in surgery
C0261555|ICD9CM|PT|E874.1|Mechanical failure of instrument or apparatus during infusion and transfusion
C0261555|ICD9CM|AB|E874.1|Instrumnt fail-infusion
C0261556|ICD9CM|PT|E874.2|Mechanical failure of instrument or apparatus during kidney dialysis and other perfusion
C0261556|ICD9CM|AB|E874.2|Instrmnt fail-perfus NEC
C0261557|ICD9CM|PT|E874.3|Mechanical failure of instrument or apparatus during endoscopic examination
C0261557|ICD9CM|AB|E874.3|Instrumnt fail-endoscopy
C0261558|ICD9CM|PT|E874.4|Mechanical failure of instrument or apparatus during aspiration of fluid or tissue, puncture, and catheterization
C0261558|ICD9CM|AB|E874.4|Instrmnt fail-catheteriz
C0261559|ICD9CM|PT|E874.5|Mechanical failure of instrument or apparatus during heart catheterization
C0261559|ICD9CM|AB|E874.5|Instrmnt fail-heart cath
C0261560|ICD9CM|PT|E874.8|Mechanical failure of instrument or apparatus during other specified procedures
C0261560|ICD9CM|AB|E874.8|Instrmnt fail-proced NEC
C0261561|ICD9CM|PT|E874.9|Mechanical failure of instrument or apparatus during unspecified procedure
C0261561|ICD9CM|AB|E874.9|Instrmnt fail-proced NOS
C0261562|ICD9CM|HT|E875|Contaminated or infected blood, other fluid, drug, or biological substance
C0261565|ICD9CM|PT|E875.2|Contaminated drug or biological substance administered by other means
C0261565|ICD9CM|AB|E875.2|Contaminated drug NEC
C0261566|ICD9CM|PT|E875.8|Misadventure to patient from other contamination
C0261566|ICD9CM|AB|E875.8|Contamination NEC
C0261567|ICD9CM|PT|E875.9|Misadventure to patient from unspecified contamination
C0261567|ICD9CM|AB|E875.9|Contamination NOS
C0261568|ICD9CM|HT|E876|Other and unspecified misadventures during medical care
C0261570|ICD9CM|AB|E876.1|Wrong fluid in infusion
C0261570|ICD9CM|PT|E876.1|Wrong fluid in infusion
C0261572|ICD9CM|PT|E876.3|Endotracheal tube wrongly placed during anesthetic procedure
C0261572|ICD9CM|AB|E876.3|Misplaced endotrach tube
C0261573|ICD9CM|PT|E876.4|Failure to introduce or to remove other tube or instrument
C0261573|ICD9CM|AB|E876.4|Fail introd/remove tube
C0261575|ICD9CM|PT|E876.8|Other specified misadventures during medical care
C0261575|ICD9CM|AB|E876.8|Medical misadventure NEC
C0261577|ICD9CM|HT|E878|Surgical operation and other surgical procedures as the cause of abnormal reaction of patient, or of later complication, without mention of misadventure at the time of operation
C0261578|ICD9CM|PT|E878.0|Surgical operation with transplant of whole organ causing abnormal patient reaction, or later complication, without mention of misadventure at time of operation
C0261578|ICD9CM|AB|E878.0|Abn react-org transplant
C0261579|ICD9CM|PT|E878.1|Surgical operation with implant of artificial internal device causing abnormal patient reaction, or later complication,without mention of misadventure at time of operation
C0261579|ICD9CM|AB|E878.1|Abn react-artif implant
C0261580|ICD9CM|PT|E878.2|Surgical operation with anastomosis, bypass, or graft, with natural or artificial tissues used as implant causing abnormal patient reaction, or later complication, without mention of misadventure at time of operation
C0261580|ICD9CM|AB|E878.2|Abn react-anastom/graft
C0261584|ICD9CM|PT|E878.6|Removal of other organ (partial) (total) causing abnormal patient reaction, or later complication, without mention of misadventure at time of operation
C0261584|ICD9CM|AB|E878.6|Abn reac-organ rem NEC
C0261585|ICD9CM|PT|E878.8|Other specified surgical operations and procedures causing abnormal patient reaction, or later complication, without mention of misadventure at time of operation
C0261585|ICD9CM|AB|E878.8|Abn react-surg proc NEC
C0261586|ICD9CM|PT|E878.9|Unspecified surgical operations and procedures causing abnormal patient reaction, or later complication, without mention of misadventure at time of operation
C0261586|ICD9CM|AB|E878.9|Abn react-surg proc NOS
C0261587|ICD9CM|HT|E879|Other procedures, without mention of misadventure at the time of procedure, as the cause of abnormal reaction of patient, or of later complication
C0261588|ICD9CM|PT|E879.0|Cardiac catheterization as the cause of abnormal reaction of patient, or of later complication, without mention of misadventure at time of procedure
C0261588|ICD9CM|AB|E879.0|Abn react-cardiac cath
C0261589|ICD9CM|PT|E879.1|Kidney dialysis as the cause of abnormal reaction of patient, or of later complication, without mention of misadventure at time of procedure
C0261589|ICD9CM|AB|E879.1|Abn react-renal dialysis
C0261590|ICD9CM|PT|E879.2|Radiological procedure and radiotherapy as the cause of abnormal reaction of patient, or of later complication, without mention of misadventure at time of procedure
C0261590|ICD9CM|AB|E879.2|Abn react-radiotherapy
C0261591|ICD9CM|PT|E879.3|Shock therapy as the cause of abnormal reaction of patient, or of later complication, without mention of misadventure at time of procedure
C0261591|ICD9CM|AB|E879.3|Abn react-shock therapy
C0261592|ICD9CM|PT|E879.4|Aspiration of fluid as the cause of abnormal reaction of patient, or of later complication, without mention of misadventure at time of procedure
C0261592|ICD9CM|AB|E879.4|Abn react-fluid aspirat
C0261594|ICD9CM|PT|E879.6|Urinary catheterization as the cause of abnormal reaction of patient, or of later complication, without mention of misadventure at time of procedure
C0261594|ICD9CM|AB|E879.6|Abn react-urinary cath
C0261595|ICD9CM|PT|E879.7|Blood sampling as the cause of abnormal reaction of patient, or of later complication, without mention of misadventure at time of procedure
C0261595|ICD9CM|AB|E879.7|Abn react-blood sampling
C0261596|ICD9CM|PT|E879.8|Other specified procedures as the cause of abnormal reaction of patient, or of later complication, without mention of misadventure at time of procedure
C0261596|ICD9CM|AB|E879.8|Abn react-procedure NEC
C0261597|ICD9CM|PT|E879.9|Unspecified procedure as the cause of abnormal reaction of patient, or of later complication, without mention of misadventure at time of procedure
C0261597|ICD9CM|AB|E879.9|Abn react-procedure NOS
C0261598|ICD9CM|HT|E880|Accidental fall on or from stairs or steps
C0261599|ICD9CM|AB|E880.0|Fall on escalator
C0261599|ICD9CM|PT|E880.0|Accidental fall on or from escalator
C0261600|ICD9CM|PT|E880.9|Accidental fall on or from other stairs or steps
C0261600|ICD9CM|AB|E880.9|Fall on stair/step NEC
C0261601|ICD9CM|HT|E881|Accidental fall on or from ladders or scaffolding
C0261603|ICD9CM|PT|E881.1|Accidental fall from scaffolding
C0261603|ICD9CM|AB|E881.1|Fall from scaffolding
C0261604|ICD9CM|PT|E882|Accidental fall from or out of building or other structure
C0261604|ICD9CM|AB|E882|Fall from building
C0261605|ICD9CM|HT|E883|Accidental fall into hole or other opening in surface
C0261606|ICD9CM|PT|E883.0|Accident from diving or jumping into water [swimming pool]
C0261606|ICD9CM|AB|E883.0|Diving accident
C0261607|ICD9CM|PT|E883.1|Accidental fall into well
C0261607|ICD9CM|AB|E883.1|Fall into well
C0261608|ICD9CM|PT|E883.2|Accidental fall into storm drain or manhole
C0261608|ICD9CM|AB|E883.2|Fall into storm drain
C0261609|ICD9CM|PT|E883.9|Accidental fall into other hole or other opening in surface
C0261609|ICD9CM|AB|E883.9|Fall into other hole
C0261611|ICD9CM|PT|E884.0|Accidental fall from playground equipment
C0261611|ICD9CM|AB|E884.0|Fall from playgrnd equip
C0261612|ICD9CM|PT|E884.1|Accidental fall from cliff
C0261612|ICD9CM|AB|E884.1|Fall from cliff
C0261613|ICD9CM|AB|E884.2|Fall from chair
C0261613|ICD9CM|PT|E884.2|Accidental fall from chair
C0261615|ICD9CM|HT|E885|Fall on same level from slipping, tripping, or stumbling
C0261617|ICD9CM|PT|E886.0|Fall on same level from collision, pushing, or shoving, by or with other person in sports
C0261617|ICD9CM|AB|E886.0|Fall in sports
C0261618|ICD9CM|PT|E886.9|Other and unspecified falls on same level from collision, pushing, or shoving, by or with other person
C0261618|ICD9CM|AB|E886.9|Fall on level NEC/NOS
C0261619|ICD9CM|HT|E888|Other and unspecified accidental fall
C0261620|ICD9CM|HT|E890|Conflagration in private dwelling
C0261621|ICD9CM|PT|E890.0|Explosion caused by conflagration in private dwelling
C0261621|ICD9CM|AB|E890.0|Privat dwell fire-explos
C0261623|ICD9CM|PT|E890.2|Other smoke and fumes from conflagration in private dwelling
C0261623|ICD9CM|AB|E890.2|Priv dwel fire-fumes NOS
C0261624|ICD9CM|PT|E890.3|Burning caused by conflagration in private dwelling
C0261624|ICD9CM|AB|E890.3|Priv dwel fire-burning
C0261625|ICD9CM|PT|E890.8|Other accident resulting from conflagration in private dwelling
C0261625|ICD9CM|AB|E890.8|Priv dwel fire-accid NEC
C0261626|ICD9CM|PT|E890.9|Unspecified accident resulting from conflagration in private dwelling
C0261626|ICD9CM|AB|E890.9|Priv dwel fire-accid NOS
C0261627|ICD9CM|HT|E891|Conflagration in other and unspecified building or structure
C0261628|ICD9CM|PT|E891.0|Explosion caused by conflagration in other and unspecified building or structure
C0261628|ICD9CM|AB|E891.0|Fire in bldg-explosion
C0261629|ICD9CM|PT|E891.1|Fumes from combustion of polyvinylchloride [pvc] and similar material in conflagration in other and unspecified building or structure
C0261629|ICD9CM|AB|E891.1|Fire in bldg-pvc fumes
C0261630|ICD9CM|PT|E891.2|Other smoke and fumes from conflagration in other and unspecified building or structure
C0261630|ICD9CM|AB|E891.2|Fire in bldg-fumes NOS
C0261631|ICD9CM|PT|E891.3|Burning caused by conflagration in other and unspecified building or structure
C0261631|ICD9CM|AB|E891.3|Fire in bldg-burning
C0261633|ICD9CM|PT|E891.9|Unspecified accident resulting from conflagration of other and unspecified building or structure
C0261633|ICD9CM|AB|E891.9|Fire in bldg-accid NOS
C0261634|ICD9CM|PT|E892|Conflagration not in building or structure
C0261634|ICD9CM|AB|E892|Fire not in building
C0261635|ICD9CM|HT|E893|Accident caused by ignition of clothing
C0261637|ICD9CM|PT|E893.1|Accident caused by ignition of clothing from controlled fire in other building or structure
C0261637|ICD9CM|AB|E893.1|Clothing fire-bldg NEC
C0261638|ICD9CM|PT|E893.2|Accident caused by ignition of clothing from controlled fire not in building or structure
C0261638|ICD9CM|AB|E893.2|Clothing fire not in bld
C0261639|ICD9CM|PT|E893.8|Accident caused by ignition of clothing from other specified sources
C0261639|ICD9CM|AB|E893.8|Clothing fire NEC
C0261641|ICD9CM|PT|E894|Ignition of highly inflammable material
C0261641|ICD9CM|AB|E894|Fire-highly inflam mater
C0261642|ICD9CM|PT|E895|Accident caused by controlled fire in private dwelling
C0261642|ICD9CM|AB|E895|Burn acc in privat dwell
C0261644|ICD9CM|PT|E897|Accident caused by controlled fire not in building or structure
C0261644|ICD9CM|AB|E897|Burn acc not in bldg
C0261645|ICD9CM|HT|E898|Accident caused by other specified fire and flames
C0261647|ICD9CM|PT|E898.1|Accident caused by other burning materials
C0261647|ICD9CM|AB|E898.1|Fire accident NEC
C0261648|ICD9CM|HT|E900|Accident caused by excessive heat
C0261649|ICD9CM|PT|E900.1|Accidents due to excessive heat of man-made origin
C0261649|ICD9CM|AB|E900.1|Excessive heat, man-made
C0261650|ICD9CM|HT|E901|Accidents due to excessive cold
C0261651|ICD9CM|PT|E901.1|Accident due to excessive cold of man-made origin
C0261651|ICD9CM|AB|E901.1|Excessive cold, man-made
C0261652|ICD9CM|PT|E901.8|Accident due to excessive cold of other specified origin
C0261652|ICD9CM|AB|E901.8|Excessive cold NEC
C0261654|ICD9CM|HT|E902|Accident due to high and low air pressure and changes in air pressure
C0261655|ICD9CM|PT|E902.1|Accident due to changes in air pressure in aircraft
C0261655|ICD9CM|AB|E902.1|Air press chnge: aircrft
C0261656|ICD9CM|PT|E902.8|Accident due to changes in air pressure due to other specified causes
C0261656|ICD9CM|AB|E902.8|Air pressure change NEC
C0261657|ICD9CM|PT|E902.9|Accident due to changes in air pressure from unspecified cause
C0261657|ICD9CM|AB|E902.9|Air pressure change NOS
C0261658|ICD9CM|HT|E904|Hunger, thirst, exposure, and neglect
C0261659|ICD9CM|PT|E904.0|Accident due to abandonment or neglect of infants and helpless persons
C0261659|ICD9CM|AB|E904.0|Abandonment/lack of care
C0261662|ICD9CM|HT|E905|Venomous animals and plants as the cause of poisoning and toxic reactions
C0261663|ICD9CM|PT|E905.2|Scorpion sting causing poisoning and toxic reactions
C0261663|ICD9CM|AB|E905.2|Scorpion sting
C0261664|ICD9CM|PT|E905.3|Sting of hornets, wasps, and bees causing poisoning and toxic reactions
C0261664|ICD9CM|AB|E905.3|Hornet/wasp/bee sting
C0261665|ICD9CM|PT|E905.4|Centipede and venomous millipede (tropical) bite causing poisoning and toxic reactions
C0261665|ICD9CM|AB|E905.4|Centipede bite
C0261666|ICD9CM|PT|E905.5|Other venomous arthropods causing poisoning and toxic reactions
C0261666|ICD9CM|AB|E905.5|Venomous arthropods NEC
C0261667|ICD9CM|PT|E905.6|Venomous marine animals and plants causing poisoning and toxic reactions
C0261667|ICD9CM|AB|E905.6|Venom sea animals/plants
C0261668|ICD9CM|PT|E905.7|Poisoning and toxic reactions caused by other plants
C0261668|ICD9CM|AB|E905.7|Poisoning by other plant
C0261669|ICD9CM|PT|E905.8|Poisoning and toxic reactions caused by other specified animals and plants
C0261669|ICD9CM|AB|E905.8|Venomous bite/sting NEC
C0261670|ICD9CM|PT|E905.9|Poisoning and toxic reactions caused by unspecified animals and plants
C0261670|ICD9CM|AB|E905.9|Venomous bite/sting NOS
C0261674|ICD9CM|PT|E906.8|Other specified injury caused by animal
C0261674|ICD9CM|AB|E906.8|Inj NEC caused by animal
C0261675|ICD9CM|PT|E906.9|Unspecified injury caused by animal
C0261675|ICD9CM|AB|E906.9|Inj NOS caused by animal
C0261676|ICD9CM|HT|E908|Accident due to cataclysmic storms, and floods resulting from storms
C0261676|ICD9CM|PT|E908.9|Unspecified cataclysmic storms, and floods resulting from storms
C0261676|ICD9CM|AB|E908.9|Acc d/t storm/flood NOS
C0261677|ICD9CM|HT|E909|Accident due to cataclysmic earth surface movements and eruptions
C0261678|ICD9CM|HT|E910|Accidental drowning and submersion
C0261679|ICD9CM|PT|E910.0|Accidental drowning and submersion while water-skiing
C0261679|ICD9CM|AB|E910.0|Water-skiing accident
C0261681|ICD9CM|PT|E910.2|Accidental drowning and submersion while engaged in other sport or recreational activity without diving equipment
C0261681|ICD9CM|AB|E910.2|Swimming accident NOS
C0261682|ICD9CM|PT|E910.3|Accidental drowning and submersion while swimming or diving for purposes other than recreation or sport
C0261682|ICD9CM|AB|E910.3|Swimming/diving acc NEC
C0261683|ICD9CM|PT|E910.4|Accidental drowning and submersion in bathtub
C0261683|ICD9CM|AB|E910.4|Drowning in bathtub
C0261684|ICD9CM|PT|E910.9|Unspecified accidental drowning or submersion
C0261684|ICD9CM|AB|E910.9|Accidental drowning NOS
C0261685|ICD9CM|PT|E911|Inhalation and ingestion of food causing obstruction of respiratory tract or suffocation
C0261685|ICD9CM|AB|E911|Resp obstr-food inhal
C0261686|ICD9CM|PT|E912|Inhalation and ingestion of other object causing obstruction of respiratory tract or suffocation
C0261686|ICD9CM|AB|E912|Resp obstr-inhal obj NEC
C0261688|ICD9CM|PT|E913.0|Accidental mechanical suffocation in bed or cradle
C0261688|ICD9CM|AB|E913.0|Suffocat in bed/cradle
C0261689|ICD9CM|PT|E913.1|Accidental mechanical suffocation by plastic bag
C0261689|ICD9CM|AB|E913.1|Suffocation-plastic bag
C0261690|ICD9CM|PT|E913.2|Accidental mechanical suffocation due to lack of air (in closed place)
C0261690|ICD9CM|AB|E913.2|Suffocation-lack of air
C0261691|ICD9CM|PT|E913.3|Accidental mechanical suffocation by falling earth or other substance
C0261691|ICD9CM|AB|E913.3|Cave-in NOS
C0261692|ICD9CM|PT|E913.8|Accidental mechanical suffocation by other specified means
C0261692|ICD9CM|AB|E913.8|Suffocation NEC
C0261693|ICD9CM|PT|E914|Foreign body accidentally entering eye and adnexa
C0261693|ICD9CM|AB|E914|FB entering eye
C0261694|ICD9CM|PT|E915|Foreign body accidentally entering other orifice
C0261694|ICD9CM|AB|E915|FB entering oth orifice
C0261695|ICD9CM|PT|E916|Struck accidentally by falling object
C0261695|ICD9CM|AB|E916|Struck by falling object
C0261696|ICD9CM|HT|E917|Striking against or struck accidentally by objects or persons
C0261703|ICD9CM|PT|E919.0|Accidents caused by agricultural machines
C0261703|ICD9CM|AB|E919.0|Machine accid-agricult
C0261704|ICD9CM|PT|E919.1|Accidents caused by mining and earth-drilling machinery
C0261704|ICD9CM|AB|E919.1|Machine accid-mining
C0261705|ICD9CM|PT|E919.2|Accidents caused by lifting machines and appliances
C0261705|ICD9CM|AB|E919.2|Lifting machine accident
C0261706|ICD9CM|PT|E919.3|Accidents caused by metalworking machines
C0261706|ICD9CM|AB|E919.3|Metalworking machine acc
C0261707|ICD9CM|PT|E919.4|Accidents caused by woodworking and forming machines
C0261707|ICD9CM|AB|E919.4|Woodworking machine acc
C0261708|ICD9CM|PT|E919.5|Accidents caused by prime movers, except electrical motors
C0261708|ICD9CM|AB|E919.5|Prime mover machine acc
C0261709|ICD9CM|PT|E919.6|Accidents caused by transmission machinery
C0261709|ICD9CM|AB|E919.6|Transmission machine acc
C0261710|ICD9CM|PT|E919.7|Accidents caused by earth moving, scraping, and other excavating machines
C0261710|ICD9CM|AB|E919.7|Earth moving machine acc
C0261711|ICD9CM|PT|E919.8|Accidents caused by other specified machinery
C0261711|ICD9CM|AB|E919.8|Machinery accident NEC
C0261712|ICD9CM|HT|E919|Accidents caused by machinery
C0261712|ICD9CM|PT|E919.9|Accidents caused by unspecified machinery
C0261712|ICD9CM|AB|E919.9|Machinery accident NOS
C0261713|ICD9CM|PT|E920.9|Accidents caused by unspecified cutting and piercing instrument or object
C0261713|ICD9CM|HT|E920|Accidents caused by cutting and piercing instruments or objects
C0261713|ICD9CM|AB|E920.9|Acc-cutting instrum NOS
C0261714|ICD9CM|PT|E920.0|Accidents caused by powered lawn mower
C0261714|ICD9CM|AB|E920.0|Acc-powered lawn mower
C0261715|ICD9CM|PT|E920.1|Accidents caused by other powered hand tools
C0261715|ICD9CM|AB|E920.1|Acc-power hand tool NEC
C0261716|ICD9CM|PT|E920.2|Accidents caused by powered household appliances and implements
C0261716|ICD9CM|AB|E920.2|Acc-power house applianc
C0261717|ICD9CM|PT|E920.3|Accidents caused by knives, swords, and daggers
C0261717|ICD9CM|AB|E920.3|Knife/sword/dagger acc
C0261718|ICD9CM|PT|E920.4|Accidents caused by other hand tools and implements
C0261718|ICD9CM|AB|E920.4|Accid-other hand tools
C0261719|ICD9CM|PT|E920.8|Accidents caused by other specified cutting and piercing instruments or objects
C0261719|ICD9CM|AB|E920.8|Acc-cutting instrum NEC
C0261721|ICD9CM|PT|E921.0|Accident caused by explosion of boilers
C0261721|ICD9CM|AB|E921.0|Boiler explosion
C0261722|ICD9CM|PT|E921.1|Accident caused by explosion of gas cylinders
C0261722|ICD9CM|AB|E921.1|Gas cylinder explosion
C0261723|ICD9CM|PT|E921.8|Accident caused by explosion of other specified pressure vessels
C0261723|ICD9CM|AB|E921.8|Press vessel explos NEC
C0261724|ICD9CM|HT|E921|Accident caused by explosion of pressure vessel
C0261724|ICD9CM|PT|E921.9|Accident caused by explosion of unspecified pressure vessel
C0261724|ICD9CM|AB|E921.9|Press vessel explos NOS
C0261725|ICD9CM|PT|E922.9|Accident caused by unspecified firearm missile
C0261725|ICD9CM|AB|E922.9|Firearm accident NOS
C0261726|ICD9CM|PT|E922.0|Accident caused by handgun
C0261726|ICD9CM|AB|E922.0|Handgun accident
C0261728|ICD9CM|PT|E922.2|Accident caused by hunting rifle
C0261728|ICD9CM|AB|E922.2|Hunting rifle accident
C0261729|ICD9CM|PT|E922.3|Accident caused by military firearms
C0261729|ICD9CM|AB|E922.3|Military firearm accid
C0261730|ICD9CM|PT|E922.8|Accident caused by other specified firearm missile
C0261730|ICD9CM|AB|E922.8|Firearm accident NEC
C0261731|ICD9CM|HT|E923|Accident caused by explosive material
C0261731|ICD9CM|PT|E923.9|Accident caused by unspecified explosive material
C0261731|ICD9CM|AB|E923.9|Explosives accident NOS
C0261732|ICD9CM|PT|E923.0|Accident caused by fireworks
C0261732|ICD9CM|AB|E923.0|Fireworks accident
C0261733|ICD9CM|PT|E923.1|Accident caused by blasting materials
C0261733|ICD9CM|AB|E923.1|Blasting materials accid
C0261734|ICD9CM|PT|E923.2|Accident caused by explosive gases
C0261734|ICD9CM|AB|E923.2|Explosive gases accident
C0261735|ICD9CM|PT|E923.8|Accident caused by other explosive materials
C0261735|ICD9CM|AB|E923.8|Explosives accident NEC
C0261736|ICD9CM|HT|E924|Accident caused by hot substance or object, caustic or corrosive material, and steam
C0261737|ICD9CM|PT|E924.0|Accident caused by hot liquids and vapors, including steam
C0261737|ICD9CM|AB|E924.0|Acc-hot liquid & steam
C0261738|ICD9CM|PT|E924.8|Accident caused by other hot substance or object
C0261738|ICD9CM|AB|E924.8|Hot substance accid NEC
C0261739|ICD9CM|PT|E924.9|Accident caused by unspecified hot substance or object
C0261739|ICD9CM|AB|E924.9|Hot substance accid NOS
C0261740|ICD9CM|HT|E925|Accident caused by electric current
C0261740|ICD9CM|PT|E925.9|Accident caused by unspecified electric current
C0261740|ICD9CM|AB|E925.9|Electric current acc NOS
C0261741|ICD9CM|PT|E925.0|Accident caused by domestic wiring and appliances
C0261741|ICD9CM|AB|E925.0|Domestic wiring accident
C0261742|ICD9CM|PT|E925.1|Accident caused by electric current in electric power generating plants, distribution stations, transmission lines
C0261742|ICD9CM|AB|E925.1|Electr power generat acc
C0261743|ICD9CM|PT|E925.2|Accident caused by industrial wiring, appliances, and electrical machinery
C0261743|ICD9CM|AB|E925.2|Indust wiring/machin acc
C0261744|ICD9CM|PT|E925.8|Accident caused by other electric current
C0261744|ICD9CM|AB|E925.8|Electric current acc NEC
C0261746|ICD9CM|PT|E926.0|Exposure to radiofrequency radiation
C0261746|ICD9CM|AB|E926.0|Radiofreq radiat exposur
C0261747|ICD9CM|PT|E926.1|Exposure to infra-red radiation from heaters and lamps
C0261747|ICD9CM|AB|E926.1|Infra-red appl rad exos
C0261748|ICD9CM|PT|E926.3|Exposure to x-rays and other electromagnetic ionizing radiation
C0261748|ICD9CM|AB|E926.3|X-ray/gamma ray exposure
C0261749|ICD9CM|PT|E926.4|Exposure to lasers
C0261749|ICD9CM|AB|E926.4|Laser exposure
C0261750|ICD9CM|PT|E926.5|Exposure to radioactive isotopes
C0261750|ICD9CM|AB|E926.5|Radioact isotope exposur
C0261752|ICD9CM|PT|E928.0|Prolonged stay in weightless environment
C0261752|ICD9CM|AB|E928.0|Acc d/t weightless envir
C0261755|ICD9CM|PT|E929.2|Late effects of accidental poisoning
C0261755|ICD9CM|AB|E929.2|Late eff acc poisoning
C0261756|ICD9CM|PT|E929.3|Late effects of accidental fall
C0261756|ICD9CM|AB|E929.3|Late eff accidental fall
C0261757|ICD9CM|PT|E929.4|Late effects of accident caused by fire
C0261757|ICD9CM|AB|E929.4|Late eff fire acc
C0261758|ICD9CM|PT|E929.5|Late effects of accident due to natural and environmental factors
C0261758|ICD9CM|AB|E929.5|Late eff environment acc
C0261765|ICD9CM|PT|E930.3|Erythromycin and other macrolides causing adverse effects in therapeutic use
C0261765|ICD9CM|AB|E930.3|Adv eff erythromycin
C0261766|ICD9CM|PT|E930.4|Tetracycline group causing adverse effects in therapeutic use
C0261766|ICD9CM|AB|E930.4|Adv eff tetracycline
C0261767|ICD9CM|PT|E930.5|Cephalosporin group causing adverse effects in therapeutic use
C0261767|ICD9CM|AB|E930.5|Adv eff cephalosporin
C0261768|ICD9CM|PT|E930.6|Antimycobacterial antibiotics causing adverse effects in therapeutic use
C0261768|ICD9CM|AB|E930.6|Adv eff antmycob antbiot
C0261769|ICD9CM|PT|E930.7|Antineoplastic antibiotics causing adverse effects in therapeutic use
C0261769|ICD9CM|AB|E930.7|Adv eff antineop antbiot
C0261770|ICD9CM|PT|E930.8|Other specified antibiotics causing adverse effects in therapeutic use
C0261770|ICD9CM|AB|E930.8|Adv eff antibiotics NEC
C0261771|ICD9CM|PT|E930.9|Unspecified antibiotic causing adverse effects in therapeutic use
C0261771|ICD9CM|HT|E930|Antibiotics causing adverse effects in therapeutic use
C0261771|ICD9CM|AB|E930.9|Adv eff antibiotic NOS
C0261772|ICD9CM|HT|E931|Other anti-infectives causing adverse effects in therapeutic use
C0261773|ICD9CM|PT|E931.0|Sulfonamides causing adverse effects in therapeutic use
C0261773|ICD9CM|AB|E931.0|Adv eff sulfonamides
C0261774|ICD9CM|PT|E931.1|Arsenical anti-infectives causing adverse effects in therapeutic use
C0261774|ICD9CM|AB|E931.1|Adv eff arsenic anti-inf
C0261775|ICD9CM|PT|E931.2|Heavy metal anti-infectives causing adverse effects in therapeutic use
C0261775|ICD9CM|AB|E931.2|Adv eff metal anti-inf
C0261776|ICD9CM|PT|E931.3|Quinoline and hydroxyquinoline derivatives causing adverse effects in therapeutic use
C0261776|ICD9CM|AB|E931.3|Adv eff quinoline
C0261777|ICD9CM|PT|E931.4|Antimalarials and drugs acting on other blood protozoa causing adverse effects in therapeutic use
C0261777|ICD9CM|AB|E931.4|Adv eff antimalarials
C0261778|ICD9CM|PT|E931.5|Other antiprotozoal drugs causing adverse effects in therapeutic use
C0261778|ICD9CM|AB|E931.5|Adv eff antprotazoal NEC
C0261780|ICD9CM|PT|E931.7|Antiviral drugs causing adverse effects in therapeutic use
C0261780|ICD9CM|AB|E931.7|Adv eff antiviral drugs
C0261781|ICD9CM|PT|E931.8|Other antimycobacterial drugs causing adverse effects in therapeutic use
C0261781|ICD9CM|AB|E931.8|Adv eff antimycobac NEC
C0261782|ICD9CM|PT|E931.9|Other and unspecified anti-infectives causing adverse effects in therapeutic use
C0261782|ICD9CM|AB|E931.9|Adv eff antinfct NEC/NOS
C0261783|ICD9CM|HT|E932|Hormones and synthetic substitutes causing adverse effects in therapeutic use
C0261784|ICD9CM|PT|E932.0|Adrenal cortical steroids causing adverse effects in therapeutic use
C0261784|ICD9CM|AB|E932.0|Adv eff corticosteroids
C0261785|ICD9CM|PT|E932.1|Androgens and anabolic congeners causing adverse effects in therapeutic use
C0261785|ICD9CM|AB|E932.1|Adv eff androgens
C0261786|ICD9CM|PT|E932.2|Ovarian hormones and synthetic substitutes causing adverse effects in therapeutic use
C0261786|ICD9CM|AB|E932.2|Adv eff ovarian hormones
C0261787|ICD9CM|PT|E932.3|Insulins and antidiabetic agents causing adverse effects in therapeutic use
C0261787|ICD9CM|AB|E932.3|Adv eff insulin/antidiab
C0261788|ICD9CM|PT|E932.4|Anterior pituitary hormones causing adverse effects in therapeutic use
C0261788|ICD9CM|AB|E932.4|Adv eff ant pituitary
C0261789|ICD9CM|PT|E932.5|Posterior pituitary hormones causing adverse effects in therapeutic use
C0261789|ICD9CM|AB|E932.5|Adv eff post pituitary
C0261790|ICD9CM|PT|E932.6|Parathyroid and parathyroid derivatives causing adverse effects in therapeutic use
C0261790|ICD9CM|AB|E932.6|Adv eff parathyroid
C0261791|ICD9CM|PT|E932.7|Thyroid and thyroid derivatives causing adverse effects in therapeutic use
C0261791|ICD9CM|AB|E932.7|Adv eff thyroid & deriv
C0261793|ICD9CM|PT|E932.9|Other and unspecified hormones and synthetic substitutes causing adverse effects in therapeutic use
C0261793|ICD9CM|AB|E932.9|Adv eff hormones NEC/NOS
C0261794|ICD9CM|HT|E933|Primarily systemic agents causing adverse effects in therapeutic use
C0261795|ICD9CM|PT|E933.0|Antiallergic and antiemetic drugs causing adverse effects in therapeutic use
C0261795|ICD9CM|AB|E933.0|Adv eff anallrg/antemet
C0261796|ICD9CM|PT|E933.1|Antineoplastic and immunosuppressive drugs causing adverse effects in therapeutic use
C0261796|ICD9CM|AB|E933.1|Adv eff antineoplastic
C0261797|ICD9CM|PT|E933.2|Acidifying agents causing adverse effects in therapeutic use
C0261797|ICD9CM|AB|E933.2|Adv eff acidifying agent
C0261798|ICD9CM|PT|E933.3|Alkalizing agents causing adverse effects in therapeutic use
C0261798|ICD9CM|AB|E933.3|Adv eff alkalizing agent
C0261801|ICD9CM|PT|E933.8|Other systemic agents, not elsewhere classified, causing adverse effects in therapeutic use
C0261801|ICD9CM|AB|E933.8|Adv eff systemic agt NEC
C0261802|ICD9CM|PT|E933.9|Unspecified systemic agent causing adverse effects in therapeutic use
C0261802|ICD9CM|AB|E933.9|Adv eff systemic agt NOS
C0261803|ICD9CM|HT|E934|Agents primarily affecting blood constituents causing adverse effects in therapeutic use
C0261804|ICD9CM|PT|E934.0|Iron and its compounds causing adverse effects in therapeutic use
C0261804|ICD9CM|AB|E934.0|Adv eff iron & compounds
C0261805|ICD9CM|PT|E934.1|Liver preparations and other antianemic agents causing adverse effects in therapeutic use
C0261805|ICD9CM|AB|E934.1|Adv eff liver/antianemic
C0261806|ICD9CM|PT|E934.2|Anticoagulants causing adverse effects in therapeutic use
C0261806|ICD9CM|AB|E934.2|Adv eff anticoagulants
C0261807|ICD9CM|PT|E934.3|Vitamin k [phytonadione] causing adverse effects in therapeutic use
C0261807|ICD9CM|AB|E934.3|Adv eff vitamin k
C0261808|ICD9CM|PT|E934.4|Fibrinolysis-affecting drugs causing adverse effects in therapeutic use
C0261808|ICD9CM|AB|E934.4|Adv eff fibrinolysis agt
C0261809|ICD9CM|PT|E934.5|Anticoagulant antagonists and other coagulants causing adverse effects in therapeutic use
C0261809|ICD9CM|AB|E934.5|Adv eff coagulants
C0261810|ICD9CM|PT|E934.6|Gamma globulin causing adverse effects in therapeutic use
C0261810|ICD9CM|AB|E934.6|Adv eff gamma globulin
C0261811|ICD9CM|PT|E934.7|Natural blood and blood products causing adverse effects in therapeutic use
C0261811|ICD9CM|AB|E934.7|Adv eff blood products
C0261812|ICD9CM|PT|E934.8|Other agents affecting blood constituents causing adverse effects in therapeutic use
C0261812|ICD9CM|AB|E934.8|Adv eff blood agent NEC
C0261813|ICD9CM|PT|E934.9|Unspecified agent affecting blood constituents causing adverse effects in therapeutic use
C0261813|ICD9CM|AB|E934.9|Adv eff blood agent NOS
C0261814|ICD9CM|HT|E935|Analgesics, antipyretics, and antirheumatics causing adverse effects in therapeutic use
C0261815|ICD9CM|PT|E935.0|Heroin causing adverse effects in therapeutic use
C0261815|ICD9CM|AB|E935.0|Adv eff heroin
C0261816|ICD9CM|PT|E935.1|Methadone causing averse effects in therapeutic use
C0261816|ICD9CM|AB|E935.1|Adv eff methadone
C0261817|ICD9CM|PT|E935.2|Other opiates and related narcotics causing adverse effects in therapeutic use
C0261817|ICD9CM|AB|E935.2|Adv eff opiates
C0261819|ICD9CM|PT|E935.4|Aromatic analgesics, not elsewhere classified, causing adverse effects in therapeutic use
C0261819|ICD9CM|AB|E935.4|Adv eff arom analgsc NEC
C0261820|ICD9CM|PT|E935.5|Pyrazole derivatives causing adverse effects in therapeutic use
C0261820|ICD9CM|AB|E935.5|Adv eff pyrazole deriv
C0261822|ICD9CM|PT|E935.7|Other non-narcotic analgesics causing adverse effects in therapeutic use
C0261822|ICD9CM|AB|E935.7|Adv eff non-narc analgsc
C0261823|ICD9CM|PT|E935.8|Other specified analgesics and antipyretics causing adverse effects in therapeutic use
C0261823|ICD9CM|AB|E935.8|Adv eff analgesics NEC
C0261824|ICD9CM|PT|E935.9|Unspecified analgesic and antipyretic causing adverse effects in therapeutic use
C0261824|ICD9CM|AB|E935.9|Adv eff analgesic NOS
C0261826|ICD9CM|PT|E936.0|Oxazolidine derivatives causing adverse effects in therapeutic use
C0261826|ICD9CM|AB|E936.0|Adv eff oxazolidin deriv
C0261827|ICD9CM|PT|E936.1|Hydantoin derivatives causing adverse effects in therapeutic use
C0261827|ICD9CM|AB|E936.1|Adv eff hydantoin deriv
C0261829|ICD9CM|PT|E936.3|Other and unspecified anticonvulsants causing adverse effects in therapeutic use
C0261829|ICD9CM|AB|E936.3|Adv eff antconvl NEC/NOS
C0261831|ICD9CM|HT|E937|Sedatives and hypnotics causing adverse effects in therapeutic use
C0261832|ICD9CM|PT|E937.0|Barbiturates causing adverse effects in therapeutic use
C0261832|ICD9CM|AB|E937.0|Adv eff barbiturates
C0261833|ICD9CM|PT|E937.1|Chloral hydrate group causing adverse effects in therapeutic use
C0261833|ICD9CM|AB|E937.1|Adv eff chloral hydrate
C0261835|ICD9CM|PT|E937.3|Bromine compounds causing adverse effects in therapeutic use
C0261835|ICD9CM|AB|E937.3|Adv eff bromine compnds
C0261836|ICD9CM|PT|E937.4|Methaqualone compounds causing adverse effects in therapeutic use
C0261836|ICD9CM|AB|E937.4|Adv eff methaqualone
C0261837|ICD9CM|PT|E937.5|Glutethimide group causing adverse effects in therapeutic use
C0261837|ICD9CM|AB|E937.5|Adv eff glutethimide
C0261838|ICD9CM|PT|E937.6|Mixed sedatives, not elsewhere classified, causing adverse effects in therapeutic use
C0261838|ICD9CM|AB|E937.6|Adv eff mix sedative
C0261839|ICD9CM|PT|E937.8|Other sedatives and hypnotics causing adverse effects in therapeutic use
C0261839|ICD9CM|AB|E937.8|Adv eff sedat/hypnot NEC
C0261840|ICD9CM|PT|E937.9|Unspecified sedatives and hypnotics causing adverse effects in therapeutic use
C0261840|ICD9CM|AB|E937.9|Adv eff sedat/hypnot NOS
C0261841|ICD9CM|HT|E938|Other central nervous system depressants and anesthetics causing adverse effects in therapeutic use
C0261842|ICD9CM|PT|E938.0|Central nervous system muscle-tone depressants causing adverse effects in therapeutic use
C0261842|ICD9CM|AB|E938.0|Adv eff cns muscl depres
C0261843|ICD9CM|PT|E938.1|Halothane causing adverse effects in therapeutic use
C0261843|ICD9CM|AB|E938.1|Adv eff halothane
C0261844|ICD9CM|PT|E938.2|Other gaseous anesthetics causing adverse effects in therapeutic use
C0261844|ICD9CM|AB|E938.2|Adv eff gas anesthet NEC
C0261845|ICD9CM|PT|E938.3|Intravenous anesthetics causing adverse effects in therapeutic use
C0261845|ICD9CM|AB|E938.3|Adv eff intraven anesth
C0261846|ICD9CM|PT|E938.4|Other and unspecified general anesthetics causing adverse effects in therapeutic use
C0261846|ICD9CM|AB|E938.4|Adv eff gen anes NEC/NOS
C0261848|ICD9CM|PT|E938.6|Peripheral nerve- and plexus-blocking anesthetics causing adverse effects in therapeutic use
C0261848|ICD9CM|AB|E938.6|Adv eff nerve-block anes
C0261849|ICD9CM|PT|E938.7|Spinal anesthetics causing adverse effects in therapeutic use
C0261849|ICD9CM|AB|E938.7|Adv eff spinal anesthet
C0261850|ICD9CM|PT|E938.9|Other and unspecified local anesthetics causing adverse effects in therapeutic use
C0261850|ICD9CM|AB|E938.9|Adv eff loc anes NEC/NOS
C0261851|ICD9CM|HT|E939|Psychotropic agents causing adverse effects in therapeutic use
C0261852|ICD9CM|PT|E939.0|Antidepressants causing adverse effects in therapeutic use
C0261852|ICD9CM|AB|E939.0|Adv eff antidepressants
C0261853|ICD9CM|PT|E939.1|Phenothiazine-based tranquilizers causing adverse effects in therapeutic use
C0261853|ICD9CM|AB|E939.1|Adv eff phenothiaz tranq
C0261854|ICD9CM|PT|E939.2|Butyrophenone-based tranquilizers causing adverse effects in therapeutic use
C0261854|ICD9CM|AB|E939.2|Adv eff butyrophen tranq
C0261855|ICD9CM|PT|E939.3|Other antipsychotics, neuroleptics, and major tranquilizers causing adverse effects in therapeutic use
C0261855|ICD9CM|AB|E939.3|Adv eff antipsychotc NEC
C0261856|ICD9CM|PT|E939.4|Benzodiazepine-based tranquilizers causing adverse effects in therapeutic use
C0261856|ICD9CM|AB|E939.4|Adv eff benzodiaz tranq
C0261857|ICD9CM|PT|E939.5|Other tranquilizers causing adverse effects in therapeutic use
C0261857|ICD9CM|AB|E939.5|Adv eff tranquilizer NEC
C0261858|ICD9CM|PT|E939.6|Psychodysleptics [hallucinogens] causing adverse effects in therapeutic use
C0261858|ICD9CM|AB|E939.6|Adv eff hallucinogens
C0261859|ICD9CM|PT|E939.7|Psychostimulants causing adverse effects in therapeutic use
C0261859|ICD9CM|AB|E939.7|Adv eff psychostimulants
C0261860|ICD9CM|PT|E939.8|Other psychotropic agents causing adverse effects in therapeutic use
C0261860|ICD9CM|AB|E939.8|Adv eff psychotropic NEC
C0261861|ICD9CM|PT|E939.9|Unspecified psychotropic agent causing adverse effects in therapeutic use
C0261861|ICD9CM|AB|E939.9|Adv eff psychotropic NOS
C0261863|ICD9CM|PT|E940.0|Analeptics causing adverse effects in therapeutic use
C0261863|ICD9CM|AB|E940.0|Adv eff analeptics
C0261864|ICD9CM|PT|E940.1|Opiate antagonists causing adverse effects in therapeutic use
C0261864|ICD9CM|AB|E940.1|Adv eff opiat antagonist
C0261865|ICD9CM|PT|E940.8|Other specified central nervous system stimulants causing adverse effects in therapeutic use
C0261865|ICD9CM|AB|E940.8|Adv eff cns stimulnt NEC
C0261868|ICD9CM|PT|E941.0|Parasympathomimetics [cholinergics] causing adverse effects in therapeutic use
C0261868|ICD9CM|AB|E941.0|Adv eff cholinergics
C0261869|ICD9CM|PT|E941.1|Parasympatholytics [anticholinergics and antimuscarinics] and spasmolytics causing adverse effects in therapeutic use
C0261869|ICD9CM|AB|E941.1|Adv eff parasympatholytc
C0261870|ICD9CM|PT|E941.2|Sympathomimetics [adrenergics] causing adverse effects in therapeutic use
C0261870|ICD9CM|AB|E941.2|Adv eff sympathomimetics
C0261871|ICD9CM|PT|E941.3|Sympatholytics [antiadrenergics] causing adverse effects in therapeutic use
C0261871|ICD9CM|AB|E941.3|Adv eff sympatholytics
C0261872|ICD9CM|PT|E941.9|Unspecified drug primarily affecting the autonomic nervous system causing adverse effects in therapeutic use
C0261872|ICD9CM|AB|E941.9|Adv eff autonom agnt NOS
C0261874|ICD9CM|PT|E942.0|Cardiac rhythm regulators causing adverse effects in therapeutic use
C0261874|ICD9CM|AB|E942.0|Adv eff card rhyth regul
C0261875|ICD9CM|PT|E942.1|Cardiotonic glycosides and drugs of similar action causing adverse effects in therapeutic use
C0261875|ICD9CM|AB|E942.1|Adv eff cardiotonics
C0261877|ICD9CM|PT|E942.3|Ganglion-blocking agents causing adverse effects in therapeutic use
C0261877|ICD9CM|AB|E942.3|Adv eff ganglion-block
C0261878|ICD9CM|PT|E942.4|Coronary vasodilators causing adverse effects in therapeutic use
C0261878|ICD9CM|AB|E942.4|Adv eff coronary vasodil
C0261879|ICD9CM|PT|E942.5|Other vasodilators causing adverse effects in therapeutic use
C0261879|ICD9CM|AB|E942.5|Adv eff vasodilators NEC
C0261880|ICD9CM|PT|E942.6|Other antihypertensive agents causing adverse effects in therapeutic use
C0261880|ICD9CM|AB|E942.6|Adv eff antihyperten agt
C0261882|ICD9CM|PT|E942.8|Capillary-active drugs causing adverse effects in therapeutic use
C0261882|ICD9CM|AB|E942.8|Adv eff capillary-act
C0261885|ICD9CM|PT|E943.0|Antacids and antigastric secretion drugs causing adverse effects in therapeutic use
C0261885|ICD9CM|AB|E943.0|Adv eff antacids
C0261886|ICD9CM|PT|E943.1|Irritant cathartics causing adverse effects in therapeutic use
C0261886|ICD9CM|AB|E943.1|Adv eff irrit cathartic
C0261887|ICD9CM|PT|E943.2|Emollient cathartics causing adverse effects in therapeutic use
C0261887|ICD9CM|AB|E943.2|Adv eff emoll cathartics
C0261888|ICD9CM|PT|E943.3|Other cathartics, including intestinal atonia drugs, causing adverse effects in therapeutic use
C0261888|ICD9CM|AB|E943.3|Adv eff cathartics NEC
C0261889|ICD9CM|PT|E943.4|Digestants causing adverse effects in therapeutic use
C0261889|ICD9CM|AB|E943.4|Adv eff digestants
C0261891|ICD9CM|PT|E943.6|Emetics causing adverse effects in therapeutic use
C0261891|ICD9CM|AB|E943.6|Adv eff emetics
C0261892|ICD9CM|PT|E943.8|Other specified agents primarily affecting the gastro-intestinal system causing adverse effects in therapeutic use
C0261892|ICD9CM|AB|E943.8|Adv eff GI agent NEC
C0261894|ICD9CM|HT|E944|Water, mineral, and uric acid metabolism drugs causing adverse effects in therapeutic use
C0261895|ICD9CM|PT|E944.0|Mercurial diuretics causing adverse effects in therapeutic use
C0261895|ICD9CM|AB|E944.0|Adv eff mercury diuretic
C0261896|ICD9CM|PT|E944.1|Purine derivative diuretics causing adverse effects in therapeutic use
C0261896|ICD9CM|AB|E944.1|Adv eff purine diuretics
C0261898|ICD9CM|PT|E944.3|Saluretics causing adverse effects in therapeutic use
C0261898|ICD9CM|AB|E944.3|Adv eff saluretics
C0261899|ICD9CM|PT|E944.4|Other diuretics causing adverse effects in therapeutic use
C0261899|ICD9CM|AB|E944.4|Adv eff diuretics NEC
C0261901|ICD9CM|PT|E944.6|Other mineral salts, not elsewhere classified, causing adverse effects in therapeutic use
C0261901|ICD9CM|AB|E944.6|Adv eff mineral salt NEC
C0261902|ICD9CM|PT|E944.7|Uric acid metabolism drugs causing adverse effects in therapeutic use
C0261902|ICD9CM|AB|E944.7|Adv eff uric acid metab
C0261903|ICD9CM|HT|E945|Agents primarily acting on the smooth and skeletal muscles and respiratory system causing adverse effects in therapeutic use
C0261905|ICD9CM|PT|E945.1|Smooth muscle relaxants causing adverse effects in therapeutic use
C0261905|ICD9CM|AB|E945.1|Adv eff smooth musc relx
C0261907|ICD9CM|PT|E945.3|Other and unspecified drugs acting on muscles causing adverse effects in therapeutic use
C0261907|ICD9CM|AB|E945.3|Adv eff musc agt NEC/NOS
C0261908|ICD9CM|PT|E945.4|Antitussives causing adverse effects in therapeutic use
C0261908|ICD9CM|AB|E945.4|Adv eff antitussives
C0261911|ICD9CM|PT|E945.7|Antiasthmatics causing adverse effects in therapeutic use
C0261911|ICD9CM|AB|E945.7|Adv eff antiasthmatics
C0261912|ICD9CM|PT|E945.8|Other and unspecified respiratory drugs causing adverse effects in therapeutic use
C0261912|ICD9CM|AB|E945.8|Adv eff resp drg NEC/NOS
C0261913|ICD9CM|HT|E946|Agents primarily affecting skin and mucous membrane, ophthalmological, otorhinolaryngological, and dental drugs causing adverse effects in therapeutic use
C0261914|ICD9CM|PT|E946.0|Local anti-infectives and anti-inflammatory drugs causing adverse effects in therapeutic use
C0261914|ICD9CM|AB|E946.0|Adv eff loc anti-infectv
C0261915|ICD9CM|PT|E946.1|Antipruritics causing adverse effects in therapeutic use
C0261915|ICD9CM|AB|E946.1|Adv eff antipruritics
C0261919|ICD9CM|PT|E946.5|Eye anti-infectives and other eye drugs causing adverse effects in therapeutic use
C0261919|ICD9CM|AB|E946.5|Adv eff eye anti-inf/drg
C0261920|ICD9CM|PT|E946.6|Anti-infectives and other drugs and preparations for ear, nose, and throat causing adverse effects in therapeutic use
C0261920|ICD9CM|AB|E946.6|Adv eff ent anti-inf/drg
C0261921|ICD9CM|PT|E946.7|Dental drugs topically applied causing adverse effects in therapeutic use
C0261921|ICD9CM|AB|E946.7|Adv eff topic dental drg
C0261922|ICD9CM|PT|E946.8|Other agents primarily affecting skin and mucous membrane causing adverse effects in therapeutic use
C0261922|ICD9CM|AB|E946.8|Adv eff skin agent NEC
C0261923|ICD9CM|PT|E946.9|Unspecified agent primarily affecting skin and mucous membrane causing adverse effects in therapeutic use
C0261923|ICD9CM|AB|E946.9|Adv eff skin agent NOS
C0261925|ICD9CM|PT|E947.0|Dietetics causing adverse effects in therapeutic use
C0261925|ICD9CM|AB|E947.0|Adv eff dietetics
C0261926|ICD9CM|PT|E947.1|Lipotropic drugs causing adverse effects in therapeutic use
C0261926|ICD9CM|AB|E947.1|Adv eff lipotropic drugs
C0261928|ICD9CM|PT|E947.3|Alcohol deterrents causing adverse effects in therapeutic use
C0261928|ICD9CM|AB|E947.3|Adv eff alcohol deter
C0261929|ICD9CM|PT|E947.4|Pharmaceutical excipients causing adverse effects in therapeutic use
C0261929|ICD9CM|AB|E947.4|Adv eff pharmaceut excip
C0261930|ICD9CM|PT|E947.8|Other drugs and medicinal substances causing adverse effects in therapeutic use
C0261930|ICD9CM|HT|E947|Other and unspecified drugs and medicinal substances causing adverse effects in therapeutic use
C0261930|ICD9CM|AB|E947.8|Adv eff medicinal NEC
C0261933|ICD9CM|PT|E948.1|Typhoid and paratyphoid vaccines causing adverse effects in therapeutic use
C0261933|ICD9CM|AB|E948.1|Adv eff typhoid vaccine
C0261934|ICD9CM|PT|E948.2|Cholera vaccine causing adverse effects in therapeutic use
C0261934|ICD9CM|AB|E948.2|Adv eff cholera vaccine
C0261936|ICD9CM|PT|E948.4|Tetanus vaccine causing adverse effects in therapeutic use
C0261936|ICD9CM|AB|E948.4|Adv eff tetanus vaccine
C0261937|ICD9CM|PT|E948.5|Diphtheria vaccine causing adverse effects in therapeutic use
C0261937|ICD9CM|AB|E948.5|Adv eff diphther vaccine
C0261938|ICD9CM|PT|E948.6|Pertussis vaccine, including combinations with a pertussis component, causing adverse effects in therapeutic use
C0261938|ICD9CM|AB|E948.6|Adv eff pertussis vaccin
C0261939|ICD9CM|PT|E948.8|Other and unspecified bacterial vaccines causing adverse effects in therapeutic use
C0261939|ICD9CM|AB|E948.8|Adv eff bact vac NEC/NOS
C0261940|ICD9CM|PT|E948.9|Mixed bacterial vaccines, except combinations with a pertussis component, causing adverse effects in therapeutic use
C0261940|ICD9CM|AB|E948.9|Adv eff mix bact vaccine
C0261942|ICD9CM|PT|E949.0|Smallpox vaccine causing adverse effects in therapeutic use
C0261942|ICD9CM|AB|E949.0|Adv eff smallpox vaccine
C0261943|ICD9CM|PT|E949.1|Rabies vaccine causing adverse effects in therapeutic use
C0261943|ICD9CM|AB|E949.1|Adv eff rabies vaccine
C0261944|ICD9CM|PT|E949.2|Typhus vaccine causing adverse effects in therapeutic use
C0261944|ICD9CM|AB|E949.2|Adv eff typhus vaccine
C0261945|ICD9CM|PT|E949.3|Yellow fever vaccine causing adverse effects in therapeutic use
C0261945|ICD9CM|AB|E949.3|Adv eff yellow fever vac
C0261946|ICD9CM|PT|E949.4|Measles vaccine causing adverse effects in therapeutic use
C0261946|ICD9CM|AB|E949.4|Adv eff measles vaccine
C0261947|ICD9CM|PT|E949.5|Poliomyelitis vaccine causing adverse effects in therapeutic use
C0261947|ICD9CM|AB|E949.5|Adv eff polio vaccine
C0261948|ICD9CM|PT|E949.6|Other and unspecified viral and rickettsial vaccines causing adverse effects in therapeutic use
C0261948|ICD9CM|AB|E949.6|Adv eff viral vacc NEC
C0261949|ICD9CM|PT|E949.7|Mixed viral-rickettsial and bacterial vaccines, except combinations with a pertussis component, causing adverse effects in therapeutic use
C0261949|ICD9CM|AB|E949.7|Adv eff mixed viral-bact
C0261950|ICD9CM|PT|E949.9|Other and unspecified vaccines and biological substances causing adverse effects in therapeutic use
C0261950|ICD9CM|HT|E949|Other vaccines and biological substances causing adverse effects in therapeutic use
C0261950|ICD9CM|AB|E949.9|Adv eff biologic NEC/NOS
C0261951|ICD9CM|HT|E950|Suicide and self-inflicted poisoning by solid or liquid substances
C0261952|ICD9CM|PT|E950.0|Suicide and self-inflicted poisoning by analgesics, antipyretics, and antirheumatics
C0261952|ICD9CM|AB|E950.0|Poison-analgesics
C0261953|ICD9CM|PT|E950.1|Suicide and self-inflicted poisoning by barbiturates
C0261953|ICD9CM|AB|E950.1|Poison-barbiturates
C0261954|ICD9CM|PT|E950.2|Suicide and self-inflicted poisoning by other sedatives and hypnotics
C0261954|ICD9CM|AB|E950.2|Poison-sedat/hypnotic
C0261955|ICD9CM|PT|E950.3|Suicide and self-inflicted poisoning by tranquilizers and other psychotropic agents
C0261955|ICD9CM|AB|E950.3|Poison-psychotropic agt
C0261956|ICD9CM|PT|E950.4|Suicide and self-inflicted poisoning by other specified drugs and medicinal substances
C0261956|ICD9CM|AB|E950.4|Poison-drug/medicin NEC
C0261957|ICD9CM|PT|E950.5|Suicide and self-inflicted poisoning by unspecified drug or medicinal substance
C0261957|ICD9CM|AB|E950.5|Poison-drug/medicin NOS
C0261958|ICD9CM|PT|E950.6|Suicide and self-inflicted poisoning by agricultural and horticultural chemical and pharmaceutical preparations other than plant foods and fertilizers
C0261958|ICD9CM|AB|E950.6|Poison-agricult agent
C0261959|ICD9CM|PT|E950.7|Suicide and self-inflicted poisoning by corrosive and caustic substances
C0261959|ICD9CM|AB|E950.7|Poison-corrosiv/caustic
C0261960|ICD9CM|PT|E950.8|Suicide and self-inflicted poisoning by arsenic and its compounds
C0261960|ICD9CM|AB|E950.8|Poison-arsenic
C0261961|ICD9CM|PT|E950.9|Suicide and self-inflicted poisoning by other and unspecified solid and liquid substances
C0261961|ICD9CM|AB|E950.9|Poison-solid/liquid NEC
C0261962|ICD9CM|HT|E951|Suicide and self-inflicted poisoning by gases in domestic use
C0261963|ICD9CM|PT|E951.0|Suicide and self-inflicted poisoning by gas distributed by pipeline
C0261963|ICD9CM|AB|E951.0|Poison-piped gas
C0261964|ICD9CM|PT|E951.1|Suicide and self-inflicted poisoning by liquefied petroleum gas distributed in mobile containers
C0261964|ICD9CM|AB|E951.1|Poison-gas in container
C0261965|ICD9CM|PT|E951.8|Suicide and self-inflicted poisoning by other utility gas
C0261965|ICD9CM|AB|E951.8|Poison-utility gas NEC
C0261966|ICD9CM|HT|E952|Suicide and self-inflicted poisoning by other gases and vapors
C0261967|ICD9CM|PT|E952.0|Suicide and self-inflicted poisoning by motor vehicle exhaust gas
C0261967|ICD9CM|AB|E952.0|Poison-exhaust gas
C0261968|ICD9CM|PT|E952.1|Suicide and self-inflicted poisoning by other carbon monoxide
C0261968|ICD9CM|AB|E952.1|Poison-co NEC
C0261969|ICD9CM|PT|E952.8|Suicide and self-inflicted poisoning by other specified gases and vapors
C0261969|ICD9CM|AB|E952.8|Poison-gas/vapor NEC
C0261970|ICD9CM|PT|E952.9|Suicide and self-inflicted poisoning by unspecified gases and vapors
C0261970|ICD9CM|AB|E952.9|Poison-gas/vapor NOS
C0261971|ICD9CM|HT|E953|Suicide and self-inflicted injury by hanging, strangulation, and suffocation
C0261972|ICD9CM|PT|E953.0|Suicide and self-inflicted injury by hanging
C0261972|ICD9CM|AB|E953.0|Injury-hanging
C0261973|ICD9CM|PT|E953.1|Suicide and self-inflicted injury by suffocation by plastic bag
C0261973|ICD9CM|AB|E953.1|Injury-suff w plas bag
C0261974|ICD9CM|PT|E953.8|Suicide and self-inflicted injury by other specified means
C0261974|ICD9CM|PT|E958.8|Suicide and self-inflicted injury by other specified means
C0261974|ICD9CM|AB|E958.8|Injury-NEC
C0261974|ICD9CM|AB|E953.8|Injury-strang/suff NEC
C0261977|ICD9CM|PT|E955.0|Suicide and self-inflicted injury by handgun
C0261977|ICD9CM|AB|E955.0|Injury-handgun
C0261978|ICD9CM|PT|E955.1|Suicide and self-inflicted injury by shotgun
C0261978|ICD9CM|AB|E955.1|Injury-shotgun
C0261979|ICD9CM|PT|E955.2|Suicide and self-inflicted injury by hunting rifle
C0261979|ICD9CM|AB|E955.2|Injury-hunting rifle
C0261980|ICD9CM|PT|E955.3|Suicide and self-inflicted injury by military firearms
C0261980|ICD9CM|AB|E955.3|Injury-military firearm
C0261981|ICD9CM|PT|E955.4|Suicide and self-inflicted injury by other and unspecified firearm
C0261981|ICD9CM|AB|E955.4|Injury-firearm NEC
C0261982|ICD9CM|PT|E955.5|Suicide and self-inflicted injury by explosives
C0261982|ICD9CM|AB|E955.5|Injury-explosives
C0261983|ICD9CM|PT|E956|Suicide and self-inflicted injury by cutting and piercing instrument
C0261983|ICD9CM|AB|E956|Injury-cut instrument
C0261984|ICD9CM|HT|E957|Suicide and self-inflicted injuries by jumping from high place
C0261985|ICD9CM|PT|E957.0|Suicide and self-inflicted injuries by jumping from residential premises
C0261985|ICD9CM|AB|E957.0|Injury-jump fm residence
C0261987|ICD9CM|PT|E957.2|Suicide and self-inflicted injuries by jumping from natural sites
C0261987|ICD9CM|AB|E957.2|Injury-jump fm natur sit
C0261988|ICD9CM|PT|E957.9|Suicide and self-inflicted injuries by jumping from unspecified site
C0261988|ICD9CM|AB|E957.9|Injury-jump NEC
C0261989|ICD9CM|HT|E958|Suicide and self-inflicted injury by other and unspecified means
C0261990|ICD9CM|PT|E958.0|Suicide and self-inflicted injury by jumping or lying before moving object
C0261990|ICD9CM|AB|E958.0|Injury-moving object
C0261991|ICD9CM|PT|E958.1|Suicide and self-inflicted injury by burns, fire
C0261991|ICD9CM|AB|E958.1|Injury-burn, fire
C0261992|ICD9CM|PT|E958.2|Suicide and self-inflicted injury by scald
C0261992|ICD9CM|AB|E958.2|Injury-scald
C0261993|ICD9CM|PT|E958.3|Suicide and self-inflicted injury by extremes of cold
C0261993|ICD9CM|AB|E958.3|Injury-extreme cold
C0261994|ICD9CM|PT|E958.4|Suicide and self-inflicted injury by electrocution
C0261994|ICD9CM|AB|E958.4|Injury-electrocution
C0261995|ICD9CM|PT|E958.5|Suicide and self-inflicted injury by crashing of motor vehicle
C0261995|ICD9CM|AB|E958.5|Injury-motor veh crash
C0261996|ICD9CM|PT|E958.6|Suicide and self-inflicted injury by crashing of aircraft
C0261996|ICD9CM|AB|E958.6|Injury-aircraft crash
C0261997|ICD9CM|PT|E958.7|Suicide and self-inflicted injury by caustic substances, except poisoning
C0261997|ICD9CM|AB|E958.7|Injury-caustic substance
C0261999|ICD9CM|HT|E960|Fight, brawl, rape
C0262000|ICD9CM|AB|E960.0|Unarmed fight or brawl
C0262000|ICD9CM|PT|E960.0|Unarmed fight or brawl
C0262001|ICD9CM|PT|E961|Assault by corrosive or caustic substance, except poisoning
C0262001|ICD9CM|AB|E961|Assault-corrosiv/caust
C0262002|ICD9CM|HT|E962|Assault by poisoning
C0262002|ICD9CM|AB|E962.9|Assault-poisoning NOS
C0262002|ICD9CM|PT|E962.9|Assault by unspecified poisoning
C0262003|ICD9CM|PT|E962.0|Assault by drugs and medicinal substances
C0262003|ICD9CM|AB|E962.0|Assault-pois w medic agt
C0262004|ICD9CM|PT|E962.1|Assault by other solid and liquid substances
C0262004|ICD9CM|AB|E962.1|Assault-pois w solid/liq
C0262005|ICD9CM|PT|E962.2|Assault by other gases and vapors
C0262005|ICD9CM|AB|E962.2|Assault-pois w gas/vapor
C0262007|ICD9CM|PT|E963|Assault by hanging and strangulation
C0262007|ICD9CM|AB|E963|Assault-hanging/strangul
C0262008|ICD9CM|PT|E964|Assault by submersion [drowning]
C0262008|ICD9CM|AB|E964|Assault-submersion
C0262009|ICD9CM|HT|E965|Assault by firearms and explosives
C0262010|ICD9CM|PT|E965.0|Assault by handgun
C0262010|ICD9CM|AB|E965.0|Assault-handgun
C0262011|ICD9CM|PT|E965.1|Assault by shotgun
C0262011|ICD9CM|AB|E965.1|Assault-shotgun
C0262012|ICD9CM|PT|E965.2|Assault by hunting rifle
C0262012|ICD9CM|AB|E965.2|Assault-hunting rifle
C0262013|ICD9CM|PT|E965.3|Assault by military firearms
C0262013|ICD9CM|AB|E965.3|Assault-military weapon
C0262015|ICD9CM|PT|E965.5|Assault by antipersonnel bomb
C0262015|ICD9CM|AB|E965.5|Assault-antiperson bomb
C0262017|ICD9CM|PT|E965.7|Assault by letter bomb
C0262017|ICD9CM|AB|E965.7|Assault-letter bomb
C0262018|ICD9CM|PT|E965.8|Assault by other specified explosive
C0262018|ICD9CM|AB|E965.8|Assault-explosive NEC
C0262019|ICD9CM|PT|E965.9|Assault by unspecified explosive
C0262019|ICD9CM|AB|E965.9|Assault-explosive NOS
C0262023|ICD9CM|PT|E967.1|Perpetrator of child and adult abuse, by other specified person
C0262023|ICD9CM|AB|E967.1|Child abuse by pers NEC
C0262024|ICD9CM|HT|E968|Assault by other and unspecified means
C0262025|ICD9CM|PT|E968.0|Assault by fire
C0262025|ICD9CM|AB|E968.0|Assault-fire
C0262027|ICD9CM|PT|E968.2|Assault by striking by blunt or thrown object
C0262027|ICD9CM|AB|E968.2|Assault-striking w obj
C0262028|ICD9CM|PT|E968.3|Assault by hot liquid
C0262028|ICD9CM|AB|E968.3|Assault-hot liquid
C0262030|ICD9CM|PT|E968.8|Assault by other specified means
C0262030|ICD9CM|AB|E968.8|Assault NEC
C0262032|ICD9CM|PT|E970|Injury due to legal intervention by firearms
C0262032|ICD9CM|AB|E970|Legal intervent-firearm
C0262033|ICD9CM|PT|E971|Injury due to legal intervention by explosives
C0262033|ICD9CM|AB|E971|Legal intervent-explosiv
C0262034|ICD9CM|PT|E972|Injury due to legal intervention by gas
C0262034|ICD9CM|AB|E972|Legal intervent-gas
C0262035|ICD9CM|PT|E973|Injury due to legal intervention by blunt object
C0262035|ICD9CM|AB|E973|Legal interven-blunt obj
C0262037|ICD9CM|PT|E975|Injury due to legal intervention by other specified means
C0262037|ICD9CM|AB|E975|Legal intervention NEC
C0262038|ICD9CM|PT|E976|Injury due to legal intervention by unspecified means
C0262038|ICD9CM|AB|E976|Legal intervention NOS
C0262040|ICD9CM|HT|E980|Poisoning by solid or liquid substances, undetermined whether accidentally or purposely inflicted
C0262041|ICD9CM|PT|E980.0|Poisoning by analgesics, antipyretics, and antirheumatics, undetermined whether accidentally or purposely inflicted
C0262041|ICD9CM|AB|E980.0|Undeterm pois-analgesics
C0262042|ICD9CM|PT|E980.1|Poisoning by barbiturates, undetermined whether accidentally or purposely inflicted
C0262042|ICD9CM|AB|E980.1|Undeterm pois-barbiturat
C0262043|ICD9CM|PT|E980.2|Poisoning by other sedatives and hypnotics, undetermined whether accidentally or purposely inflicted
C0262043|ICD9CM|AB|E980.2|Undet pois-sed/hypn NEC
C0262044|ICD9CM|PT|E980.3|Poisoning by tranquilizers and other psychotropic agents, undetermined whether accidentally or purposely inflicted
C0262044|ICD9CM|AB|E980.3|Undeterm pois-psychotrop
C0262045|ICD9CM|PT|E980.4|Poisoning by other specified drugs and medicinal substances, undetermined whether accidentally or purposely inflicted
C0262045|ICD9CM|AB|E980.4|Undet pois-med agnt NEC
C0262046|ICD9CM|PT|E980.5|Poisoning by unspecified drug or medicinal substance, undetermined whether accidentally or purposely inflicted
C0262046|ICD9CM|AB|E980.5|Undet pois-med agnt NOS
C0262047|ICD9CM|PT|E980.6|Poisoning by corrosive and caustic substances, undetermined whether accidentally or purposely inflicted
C0262047|ICD9CM|AB|E980.6|Undet pois-corros/caust
C0262048|ICD9CM|PT|E980.7|Poisoning by agricultural and horticultural chemical and pharmaceutical preparations other than plant foods and fertilizers, undetermined whether accidentally or purposely inflicted
C0262048|ICD9CM|AB|E980.7|Undet pois-agricult agnt
C0262049|ICD9CM|PT|E980.8|Poisoning by arsenic and its compounds, undetermined whether accidentally or purposely inflicted
C0262049|ICD9CM|AB|E980.8|Undeter pois-arsenic
C0262050|ICD9CM|PT|E980.9|Poisoning by other and unspecified solid and liquid substances, undetermined whether accidentally or purposely inflicted
C0262050|ICD9CM|AB|E980.9|Undeter pois-sol/liq NEC
C0262051|ICD9CM|HT|E981|Poisoning by gases in domestic use, undetermined whether accidentally or purposely inflicted
C0262052|ICD9CM|PT|E981.0|Poisoning by gas distributed by pipeline, undetermined whether accidentally or purposely inflicted
C0262052|ICD9CM|AB|E981.0|Undeter pois-piped gas
C0262053|ICD9CM|PT|E981.1|Poisoning by liquefied petroleum gas distributed in mobile containers, undetermined whether accidentally or purposely inflicted
C0262053|ICD9CM|AB|E981.1|Undet pois-container gas
C0262054|ICD9CM|PT|E981.8|Poisoning by other utility gas, undetermined whether accidentally or purposely inflicted
C0262054|ICD9CM|AB|E981.8|Undet pois-util gas NEC
C0262055|ICD9CM|HT|E982|Poisoning by other gases, undetermined whether accidentally or purposely inflicted
C0262056|ICD9CM|PT|E982.0|Poisoning by motor vehicle exhaust gas, undetermined whether accidentally or purposely inflicted
C0262056|ICD9CM|AB|E982.0|Undeter pois-exhaust gas
C0262057|ICD9CM|PT|E982.1|Poisoning by other carbon monoxide, undetermined whether accidentally or purposely inflicted
C0262057|ICD9CM|AB|E982.1|Undetermin poison-co NEC
C0262058|ICD9CM|PT|E982.8|Poisoning by other specified gases and vapors, undetermined whether accidentally or purposely inflicted
C0262058|ICD9CM|AB|E982.8|Undet pois-gas/vapor NEC
C0262059|ICD9CM|PT|E982.9|Poisoning by unspecified gases and vapors, undetermined whether accidentally or purposely inflicted
C0262059|ICD9CM|AB|E982.9|Undet pois-gas/vapor NOS
C0262060|ICD9CM|HT|E983|Hanging, strangulation, or suffocation, undetermined whether accidentally or purposely inflicted
C0262061|ICD9CM|PT|E983.0|Hanging, undetermined whether accidentally or purposely inflicted
C0262061|ICD9CM|AB|E983.0|Undetermin circ-hanging
C0262062|ICD9CM|PT|E983.1|Suffocation by plastic bag, undetermined whether accidentally or purposely inflicted
C0262062|ICD9CM|AB|E983.1|Undet circ-suf plast bag
C0262063|ICD9CM|PT|E983.8|Strangulation or suffocation by other specified means, undetermined whether accidentally or purposely inflicted
C0262063|ICD9CM|AB|E983.8|Undet circ-suffocate NEC
C0262064|ICD9CM|PT|E983.9|Strangulation or suffocation by unspecified means, undetermined whether accidentally or purposely inflicted
C0262064|ICD9CM|AB|E983.9|Undet circ-suffocate NOS
C0262065|ICD9CM|PT|E984|Submersion (drowning), undetermined whether accidentally or purposely inflicted
C0262065|ICD9CM|AB|E984|Undeterm circ-submersion
C0262067|ICD9CM|PT|E985.0|Injury by handgun, undetermined whether accidentally or purposely inflicted
C0262067|ICD9CM|AB|E985.0|Undetermin circ-handgun
C0262068|ICD9CM|PT|E985.1|Injury by shotgun, undetermined whether accidentally or purposely inflicted
C0262068|ICD9CM|AB|E985.1|Undetermin circ-shotgun
C0262069|ICD9CM|PT|E985.2|Injury by hunting rifle, undetermined whether accidentally or purposely inflicted
C0262069|ICD9CM|AB|E985.2|Undet circ-hunting rifle
C0262070|ICD9CM|PT|E985.3|Injury by military firearms, undetermined whether accidentally or purposely inflicted
C0262070|ICD9CM|AB|E985.3|Undet circ-military arms
C0262071|ICD9CM|PT|E985.4|Injury by other and unspecified firearm, undetermined whether accidentally or purposely inflicted
C0262071|ICD9CM|AB|E985.4|Undeter circ-firearm NEC
C0262072|ICD9CM|PT|E985.5|Injury by explosives, undetermined whether accidentally or purposely inflicted
C0262072|ICD9CM|AB|E985.5|Undeterm circ-explosive
C0262073|ICD9CM|PT|E986|Injury by cutting and piercing instruments, undetermined whether accidentally or purposely inflicted
C0262073|ICD9CM|AB|E986|Undet circ-cut instrumnt
C0262074|ICD9CM|HT|E987|Falling from high place, undetermined whether accidentally or purposely inflicted
C0262075|ICD9CM|PT|E987.0|Falling from residential premises, undetermined whether accidentally or purposely inflicted
C0262075|ICD9CM|AB|E987.0|Undet circ-fall residenc
C0262076|ICD9CM|PT|E987.1|Falling from other man-made structures, undetermined whether accidentally or purposely inflicted
C0262076|ICD9CM|AB|E987.1|Undet fall structure NEC
C0262077|ICD9CM|PT|E987.2|Falling from natural sites, undetermined whether accidentally or purposely inflicted
C0262077|ICD9CM|AB|E987.2|Undet fall natural site
C0262078|ICD9CM|PT|E987.9|Falling from unspecified site, undetermined whether accidentally or purposely inflicted
C0262078|ICD9CM|AB|E987.9|Undet circ-fall site NOS
C0262080|ICD9CM|PT|E988.0|Injury by jumping or lying before moving object, undetermined whether accidentally or purposely inflicted
C0262080|ICD9CM|AB|E988.0|Undeterm circ-moving obj
C0262081|ICD9CM|PT|E988.1|Injury by burns or fire, undetermined whether accidentally or purposely inflicted
C0262081|ICD9CM|AB|E988.1|Undeterm circ-burn, fire
C0262083|ICD9CM|PT|E988.3|Injury by extremes of cold, undetermined whether accidentally or purposely inflicted
C0262083|ICD9CM|AB|E988.3|Undeterm circ-extrm cold
C0262084|ICD9CM|PT|E988.4|Injury by electrocution, undetermined whether accidentally or purposely inflicted
C0262084|ICD9CM|AB|E988.4|Undeterm circ-electrocut
C0262085|ICD9CM|PT|E988.5|Injury by crashing of motor vehicle, undetermined whether accidentally or purposely inflicted
C0262085|ICD9CM|AB|E988.5|Undet circ-mot veh crash
C0262086|ICD9CM|PT|E988.6|Injury by crashing of aircraft, undetermined whether accidentally or purposely inflicted
C0262086|ICD9CM|AB|E988.6|Undet circ-aircrft crash
C0262087|ICD9CM|PT|E988.7|Injury by caustic substances, except poisoning, undetermined whether accidentally or purposely inflicted
C0262087|ICD9CM|AB|E988.7|Undet circ-caustic subst
C0262088|ICD9CM|PT|E988.8|Injury by other specified means, undetermined whether accidentally or purposely inflicted
C0262088|ICD9CM|HT|E988|Injury by other and unspecified means, undetermined whether accidentally or purposely inflicted
C0262088|ICD9CM|AB|E988.8|Undetermin circumst NEC
C0262089|ICD9CM|PT|E988.9|Injury by unspecified means, undetermined whether accidentally or purposely inflicted
C0262089|ICD9CM|AB|E988.9|Undetermin circumst NOS
C0262091|ICD9CM|HT|E990|Injury due to war operations by fires and conflagrations
C0262092|ICD9CM|PT|E990.0|Injury due to war operations from gasoline bomb
C0262092|ICD9CM|AB|E990.0|War inj:gasoline bomb
C0262093|ICD9CM|PT|E990.9|Injury due to war operations from other and unspecified source
C0262093|ICD9CM|AB|E990.9|War injury:fire NEC
C0262094|ICD9CM|HT|E991|Injury due to war operations by bullets and fragments
C0262095|ICD9CM|PT|E991.0|Injury due to war operations from rubber bullets (rifle)
C0262095|ICD9CM|AB|E991.0|War inj:rubber bullet
C0262096|ICD9CM|PT|E991.1|Injury due to war operations from pellets (rifle)
C0262096|ICD9CM|AB|E991.1|War injury:pellets
C0262097|ICD9CM|PT|E991.2|Injury due to war operations from other bullets
C0262097|ICD9CM|AB|E991.2|War injury:bullet NEC
C0262098|ICD9CM|PT|E991.3|Injury due to war operations from antipersonnel bomb (fragments)
C0262098|ICD9CM|AB|E991.3|War inj:antiperson bomb
C0262099|ICD9CM|PT|E991.9|Injury due to war operations from other and unspecified fragments
C0262099|ICD9CM|AB|E991.9|War inj:fragments NEC
C0262100|ICD9CM|HT|E992|Injury due to war operations by explosion of marine weapons
C0262101|ICD9CM|HT|E993|Injury due to war operations by other explosion
C0262102|ICD9CM|HT|E994|Injury due to war operations by destruction of aircraft
C0262103|ICD9CM|HT|E995|Injury due to war operations by other and unspecified forms of conventional warfare
C0262105|ICD9CM|HT|E997|Injury due to war operations by other forms of unconventional warfare
C0262106|ICD9CM|PT|E997.0|Injury due to war operations by lasers
C0262106|ICD9CM|AB|E997.0|War injury:lasers
C0262107|ICD9CM|PT|E997.1|Injury due to war operations by biological warfare
C0262107|ICD9CM|AB|E997.1|War injury:biol warfare
C0262108|ICD9CM|PT|E997.2|Injury due to war operations by gases, fumes, and chemicals
C0262108|ICD9CM|AB|E997.2|War injury:gas/fum/chem
C0262109|ICD9CM|PT|E997.8|Injury due to other specified forms of unconventional warfare
C0262109|ICD9CM|AB|E997.8|War inj-unconven war NEC
C0262110|ICD9CM|PT|E997.9|Injury due to unspecified form of unconventional warfare
C0262110|ICD9CM|AB|E997.9|War inj-unconven war NOS
C0262111|ICD9CM|HT|E998|Injury due to war operations but occurring after cessation of hostilities
C0262113|ICD9CM|PT|85.21|Local excision of lesion of breast
C0262113|ICD9CM|AB|85.21|Local excis breast les
C0262671|ICD9CM|AB|75.37|Amnioinfusion
C0262671|ICD9CM|PT|75.37|Amnioinfusion
C0263013|ICD9CM|AB|723.6|Panniculitis of neck
C0263013|ICD9CM|PT|723.6|Panniculitis specified as affecting neck
C0263292|ICD9CM|PT|692.70|Unspecified dermatitis due to sun
C0263292|ICD9CM|AB|692.70|Solar dermatitis NOS
C0263296|ICD9CM|PT|692.81|Dermatitis due to cosmetics
C0263296|ICD9CM|AB|692.81|Cosmetic dermatitis
C0263304|ICD9CM|PT|692.83|Dermatitis due to metals
C0263304|ICD9CM|AB|692.83|Dermatitis metals
C0263518|ICD9CM|AB|704.02|Telogen effluvium
C0263518|ICD9CM|PT|704.02|Telogen effluvium
C0263660|ICD9CM|HT|710-739.99|DISEASES OF THE MUSCULOSKELETAL SYSTEM AND CONNECTIVE TISSUE
C0263681|ICD9CM|PT|711.01|Pyogenic arthritis, shoulder region
C0263681|ICD9CM|AB|711.01|Pyogen arthritis-shlder
C0263682|ICD9CM|PT|711.02|Pyogenic arthritis, upper arm
C0263682|ICD9CM|AB|711.02|Pyogen arthritis-up/arm
C0263683|ICD9CM|PT|711.03|Pyogenic arthritis, forearm
C0263683|ICD9CM|AB|711.03|Pyogen arthritis-forearm
C0263684|ICD9CM|PT|711.04|Pyogenic arthritis, hand
C0263684|ICD9CM|AB|711.04|Pyogen arthritis-hand
C0263687|ICD9CM|PT|711.06|Pyogenic arthritis, lower leg
C0263687|ICD9CM|AB|711.06|Pyogen arthritis-l/leg
C0263690|ICD9CM|PT|711.09|Pyogenic arthritis, multiple sites
C0263690|ICD9CM|AB|711.09|Pyogen arthritis-mult
C0263708|ICD9CM|PT|712.91|Unspecified crystal arthropathy, shoulder region
C0263708|ICD9CM|AB|712.91|Cryst arthrop NOS-shldr
C0263709|ICD9CM|PT|712.92|Unspecified crystal arthropathy, upper arm
C0263709|ICD9CM|AB|712.92|Cryst arthrop NOS-up/arm
C0263710|ICD9CM|PT|712.93|Unspecified crystal arthropathy, forearm
C0263710|ICD9CM|AB|712.93|Crys arthrop NOS-forearm
C0263711|ICD9CM|PT|712.94|Unspecified crystal arthropathy, hand
C0263711|ICD9CM|AB|712.94|Cryst arthrop NOS-hand
C0263714|ICD9CM|PT|712.96|Unspecified crystal arthropathy, lower leg
C0263714|ICD9CM|AB|712.96|Cryst arthrop NOS-l/leg
C0263715|ICD9CM|PT|712.97|Unspecified crystal arthropathy, ankle and foot
C0263715|ICD9CM|AB|712.97|Cryst arthrop NOS-ankle
C0263716|ICD9CM|PT|712.98|Unspecified crystal arthropathy, other specified sites
C0263716|ICD9CM|AB|712.98|Cry arthrop NOS-oth site
C0263717|ICD9CM|PT|712.99|Unspecified crystal arthropathy, multiple sites
C0263717|ICD9CM|AB|712.99|Cryst arthrop NOS-mult
C0263723|ICD9CM|PT|713.1|Arthropathy associated with gastrointestinal conditions other than infections
C0263723|ICD9CM|AB|713.1|Arthrop w noninf GI dis
C0263724|ICD9CM|PT|713.2|Arthropathy associated with hematological disorders
C0263724|ICD9CM|AB|713.2|Arthropath w hematol dis
C0263726|ICD9CM|PT|713.3|Arthropathy associated with dermatological disorders
C0263726|ICD9CM|AB|713.3|Arthropathy w skin dis
C0263727|ICD9CM|PT|713.4|Arthropathy associated with respiratory disorders
C0263727|ICD9CM|AB|713.4|Arthropathy w resp dis
C0263730|ICD9CM|PT|713.6|Arthropathy associated with hypersensitivity reaction
C0263730|ICD9CM|AB|713.6|Arthrop w hypersen react
C0263732|ICD9CM|PT|713.8|Arthropathy associated with other conditions classifiable elsewhere
C0263732|ICD9CM|AB|713.8|Arthrop w oth dis NEC
C0263742|ICD9CM|HT|715|Osteoarthrosis and allied disorders
C0263752|ICD9CM|PT|715.11|Osteoarthrosis, localized, primary, shoulder region
C0263752|ICD9CM|AB|715.11|Loc prim osteoart-shlder
C0263753|ICD9CM|PT|715.12|Osteoarthrosis, localized, primary, upper arm
C0263753|ICD9CM|AB|715.12|Loc prim osteoart-up/arm
C0263754|ICD9CM|PT|715.13|Osteoarthrosis, localized, primary, forearm
C0263754|ICD9CM|AB|715.13|Loc prim osteoart-forarm
C0263755|ICD9CM|PT|715.14|Osteoarthrosis, localized, primary, hand
C0263755|ICD9CM|AB|715.14|Loc prim osteoarth-hand
C0263758|ICD9CM|PT|715.16|Osteoarthrosis, localized, primary, lower leg
C0263758|ICD9CM|AB|715.16|Loc prim osteoart-l/leg
C0263759|ICD9CM|PT|715.17|Osteoarthrosis, localized, primary, ankle and foot
C0263759|ICD9CM|AB|715.17|Loc prim osteoarth-ankle
C0263774|ICD9CM|HT|715.8|Osteoarthrosis involving or with mention of more than one site, but not specified as generalized
C0263793|ICD9CM|PT|718.01|Articular cartilage disorder, shoulder region
C0263793|ICD9CM|AB|718.01|Artic cartil dis-shlder
C0263794|ICD9CM|PT|718.02|Articular cartilage disorder, upper arm
C0263794|ICD9CM|AB|718.02|Artic cartil dis-up/arm
C0263795|ICD9CM|PT|718.03|Articular cartilage disorder, forearm
C0263795|ICD9CM|AB|718.03|Artic cartil dis-forearm
C0263799|ICD9CM|PT|718.07|Articular cartilage disorder, ankle and foot
C0263799|ICD9CM|AB|718.07|Artic cartil dis-ankle
C0263801|ICD9CM|PT|718.09|Articular cartilage disorder, multiple sites
C0263801|ICD9CM|AB|718.09|Artic cartil dis-mult jt
C0263805|ICD9CM|PT|718.22|Pathological dislocation of joint, upper arm
C0263805|ICD9CM|AB|718.22|Pathol dislocat-up/arm
C0263806|ICD9CM|PT|718.23|Pathological dislocation of joint, forearm
C0263806|ICD9CM|AB|718.23|Pathol dislocat-forearm
C0263809|ICD9CM|PT|718.26|Pathological dislocation of joint, lower leg
C0263809|ICD9CM|AB|718.26|Pathol dislocat-l/leg
C0263810|ICD9CM|PT|718.27|Pathological dislocation of joint, ankle and foot
C0263810|ICD9CM|AB|718.27|Pathol dislocat-ankle
C0263812|ICD9CM|PT|718.29|Pathological dislocation of joint, multiple sites
C0263812|ICD9CM|AB|718.29|Pathol dislocat-mult jts
C0263814|ICD9CM|PT|718.32|Recurrent dislocation of joint, upper arm
C0263814|ICD9CM|AB|718.32|Recur dislocat-up/arm
C0263815|ICD9CM|PT|718.33|Recurrent dislocation of joint, forearm
C0263815|ICD9CM|AB|718.33|Recur dislocat-forearm
C0263816|ICD9CM|PT|718.34|Recurrent dislocation of joint, hand
C0263816|ICD9CM|AB|718.34|Recur dislocat-hand
C0263819|ICD9CM|PT|718.36|Recurrent dislocation of joint, lower leg
C0263819|ICD9CM|AB|718.36|Recur dislocat-l/leg
C0263820|ICD9CM|PT|718.37|Recurrent dislocation of joint, ankle and foot
C0263820|ICD9CM|AB|718.37|Recur dislocat-ankle
C0263822|ICD9CM|PT|718.39|Recurrent dislocation of joint, multiple sites
C0263822|ICD9CM|AB|718.39|Recur dislocat-mult jts
C0263836|ICD9CM|PT|719.12|Hemarthrosis, upper arm
C0263836|ICD9CM|AB|719.12|Hemarthrosis-up/arm
C0263837|ICD9CM|AB|719.13|Hemarthrosis-forearm
C0263837|ICD9CM|PT|719.13|Hemarthrosis, forearm
C0263838|ICD9CM|PT|719.15|Hemarthrosis, pelvic region and thigh
C0263838|ICD9CM|AB|719.15|Hemarthrosis-pelvis
C0263840|ICD9CM|PT|719.16|Hemarthrosis, lower leg
C0263840|ICD9CM|AB|719.16|Hemarthrosis-l/leg
C0263841|ICD9CM|PT|719.17|Hemarthrosis, ankle and foot
C0263841|ICD9CM|AB|719.17|Hemarthrosis-ankle
C0263851|ICD9CM|PT|721.90|Spondylosis of unspecified site, without mention of myelopathy
C0263851|ICD9CM|AB|721.90|Spondylos NOS w/o myelop
C0263853|ICD9CM|PT|721.91|Spondylosis of unspecified site, with myelopathy
C0263853|ICD9CM|AB|721.91|Spondylosis NOS w myelop
C0263933|ICD9CM|AB|726.71|Achilles tendinitis
C0263933|ICD9CM|PT|726.71|Achilles bursitis or tendinitis
C0263962|ICD9CM|AB|726.33|Olecranon bursitis
C0263962|ICD9CM|PT|726.33|Olecranon bursitis
C0263978|ICD9CM|PT|729.90|Disorders of soft tissue, unspecified
C0263978|ICD9CM|AB|729.90|Soft tissue disord NOS
C0264022|ICD9CM|PT|730.91|Unspecified infection of bone, shoulder region
C0264022|ICD9CM|PT|730.21|Unspecified osteomyelitis, shoulder region
C0264022|ICD9CM|AB|730.21|Osteomyelitis NOS-shlder
C0264022|ICD9CM|AB|730.91|Bone infect NOS-shlder
C0264023|ICD9CM|PT|730.92|Unspecified infection of bone, upper arm
C0264023|ICD9CM|PT|730.22|Unspecified osteomyelitis, upper arm
C0264023|ICD9CM|AB|730.92|Bone infect NOS-up/arm
C0264023|ICD9CM|AB|730.22|Osteomyelitis NOS-up/arm
C0264024|ICD9CM|PT|730.93|Unspecified infection of bone, forearm
C0264024|ICD9CM|PT|730.23|Unspecified osteomyelitis, forearm
C0264024|ICD9CM|AB|730.23|Osteomyelit NOS-forearm
C0264024|ICD9CM|AB|730.93|Bone infect NOS-forearm
C0264025|ICD9CM|AB|730.24|Osteomyelitis NOS-hand
C0264025|ICD9CM|PT|730.24|Unspecified osteomyelitis, hand
C0264028|ICD9CM|PT|730.96|Unspecified infection of bone, lower leg
C0264028|ICD9CM|AB|730.96|Bone infect NOS-l/leg
C0264029|ICD9CM|PT|730.97|Unspecified infection of bone, ankle and foot
C0264029|ICD9CM|AB|730.97|Bone infect NOS-ankle
C0264031|ICD9CM|PT|730.29|Unspecified osteomyelitis, multiple sites
C0264031|ICD9CM|AB|730.29|Osteomyelitis NOS-mult
C0264039|ICD9CM|PT|730.07|Acute osteomyelitis, ankle and foot
C0264039|ICD9CM|AB|730.07|Ac osteomyelitis-ankle
C0264049|ICD9CM|PT|730.17|Chronic osteomyelitis, ankle and foot
C0264049|ICD9CM|AB|730.17|Chr osteomyelit-ankle
C0264051|ICD9CM|PT|730.19|Chronic osteomyelitis, multiple sites
C0264051|ICD9CM|AB|730.19|Chr osteomyelit-mult
C0264069|ICD9CM|HT|730.3|Periostitis without mention of osteomyelitis
C0264070|ICD9CM|PT|730.80|Other infections involving bone in diseases classified elsewhere, site unspecified
C0264070|ICD9CM|HT|730.8|Other infections involving bone in disease classified elsewhere
C0264070|ICD9CM|AB|730.80|Bone infect NEC-unspec
C0264132|ICD9CM|PT|738.9|Acquired deformity of unspecified site
C0264132|ICD9CM|AB|738.9|Acq deformity NOS
C0264133|ICD9CM|AB|734|Flat foot
C0264133|ICD9CM|PT|734|Flat foot
C0264134|ICD9CM|AB|735.2|Hallux rigidus
C0264134|ICD9CM|PT|735.2|Hallux rigidus
C0264150|ICD9CM|PT|736.70|Unspecified deformity of ankle and foot, acquired
C0264150|ICD9CM|AB|736.70|Acq ankle-foot def NOS
C0264155|ICD9CM|PT|736.9|Acquired deformity of limb, site unspecified
C0264155|ICD9CM|AB|736.9|Acq limb deformity NOS
C0264156|ICD9CM|PT|736.81|Unequal leg length (acquired)
C0264156|ICD9CM|AB|736.81|Unequal leg length
C0264222|ICD9CM|PT|465.9|Acute upper respiratory infections of unspecified site
C0264222|ICD9CM|AB|465.9|Acute uri NOS
C0264490|ICD9CM|PT|518.81|Acute respiratory failure
C0264490|ICD9CM|AB|518.81|Acute respiratry failure
C0264491|ICD9CM|PT|518.84|Acute and chronic respiratory failure
C0264491|ICD9CM|AB|518.84|Acute & chronc resp fail
C0264492|ICD9CM|PT|518.83|Chronic respiratory failure
C0264492|ICD9CM|AB|518.83|Chronic respiratory fail
C0264557|ICD9CM|AB|512.83|Chronic pneumothorax
C0264557|ICD9CM|PT|512.83|Chronic pneumothorax
C0264614|ICD9CM|PT|784.43|Hypernasality
C0264614|ICD9CM|AB|784.43|Hypernasality
C0264618|ICD9CM|AB|784.44|Hyponasality
C0264618|ICD9CM|PT|784.44|Hyponasality
C0264643|ICD9CM|PT|405.01|Malignant renovascular hypertension
C0264643|ICD9CM|AB|405.01|Mal renovasc hypertens
C0264694|ICD9CM|PT|414.9|Chronic ischemic heart disease, unspecified
C0264694|ICD9CM|AB|414.9|Chr ischemic hrt dis NOS
C0264706|ICD9CM|HT|410.6|Acute myocardial infarction, true posterior wall infarction
C0264743|ICD9CM|PT|390|Rheumatic fever without mention of heart involvement
C0264743|ICD9CM|AB|390|Rheum fev w/o hrt involv
C0264764|ICD9CM|PT|397.9|Rheumatic diseases of endocardium, valve unspecified
C0264764|ICD9CM|AB|397.9|Rheum endocarditis NOS
C0264765|ICD9CM|HT|394|Diseases of mitral valve
C0264766|ICD9CM|AB|394.0|Mitral stenosis
C0264766|ICD9CM|PT|394.0|Mitral stenosis
C0264767|ICD9CM|PT|394.2|Mitral stenosis with insufficiency
C0264767|ICD9CM|AB|394.2|Mitral stenosis w insuff
C0264772|ICD9CM|PT|396.1|Mitral valve stenosis and aortic valve insufficiency
C0264772|ICD9CM|AB|396.1|Mitral stenos/aort insuf
C0264774|ICD9CM|PT|396.3|Mitral valve insufficiency and aortic valve insufficiency
C0264774|ICD9CM|AB|396.3|Mitral/aortic val insuff
C0264776|ICD9CM|AB|397.0|Tricuspid valve disease
C0264776|ICD9CM|PT|397.0|Diseases of tricuspid valve
C0264865|ICD9CM|AB|424.90|Endocarditis NOS
C0264865|ICD9CM|HT|424.9|Endocarditis, valve unspecified
C0264865|ICD9CM|PT|424.90|Endocarditis, valve unspecified, unspecified cause
C0264886|ICD9CM|HT|426|Conduction disorders
C0264886|ICD9CM|AB|426.9|Conduction disorder NOS
C0264886|ICD9CM|PT|426.9|Conduction disorder, unspecified
C0265004|ICD9CM|HT|447.7|Aortic ectasia
C0265010|ICD9CM|PT|441.1|Thoracic aneurysm, ruptured
C0265010|ICD9CM|AB|441.1|Ruptur thoracic aneurysm
C0265011|ICD9CM|PT|441.4|Abdominal aneurysm without mention of rupture
C0265011|ICD9CM|AB|441.4|Abdom aortic aneurysm
C0265012|ICD9CM|PT|441.3|Abdominal aneurysm, ruptured
C0265012|ICD9CM|AB|441.3|Rupt abd aortic aneurysm
C0265027|ICD9CM|AB|448.1|Nevus, non-neoplastic
C0265027|ICD9CM|PT|448.1|Nevus, non-neoplastic
C0265035|ICD9CM|PT|455.0|Internal hemorrhoids without mention of complication
C0265035|ICD9CM|AB|455.0|Int hemorrhoid w/o compl
C0265041|ICD9CM|PT|455.3|External hemorrhoids without mention of complication
C0265041|ICD9CM|AB|455.3|Ext hemorrhoid w/o compl
C0265057|ICD9CM|PT|451.0|Phlebitis and thrombophlebitis of superficial vessels of lower extremities
C0265057|ICD9CM|AB|451.0|Superfic phlebitis-leg
C0265066|ICD9CM|PT|451.11|Phlebitis and thrombophlebitis of femoral vein (deep) (superficial)
C0265066|ICD9CM|AB|451.11|Femoral vein phlebitis
C0265098|ICD9CM|HT|433.0|Occlusion and stenosis of basilar artery
C0265122|ICD9CM|PT|423.9|Unspecified disease of pericardium
C0265122|ICD9CM|AB|423.9|Pericardial disease NOS
C0265547|ICD9CM|PT|755.4|Reduction deformities, unspecified limb
C0265547|ICD9CM|AB|755.4|Reduct deform limb NOS
C0265553|ICD9CM|PT|755.10|Syndactyly of multiple and unspecified sites
C0265553|ICD9CM|AB|755.10|Syndactyly, multiple/NOS
C0265566|ICD9CM|HT|755.2|Reduction deformities of upper limb, congenital
C0265566|ICD9CM|PT|755.20|Unspecified reduction deformity of upper limb
C0265566|ICD9CM|AB|755.20|Reduc deform up limb NOS
C0265609|ICD9CM|AB|755.56|Accessory carpal bones
C0265609|ICD9CM|PT|755.56|Accessory carpal bones
C0265618|ICD9CM|HT|755.3|Reduction deformities of lower limb, congenital
C0265618|ICD9CM|PT|755.30|Unspecified reduction deformity of lower limb
C0265618|ICD9CM|AB|755.30|Reduction deform leg NOS
C0265647|ICD9CM|AB|754.53|Metatarsus varus
C0265647|ICD9CM|PT|754.53|Metatarsus varus
C0265649|ICD9CM|AB|754.52|Metatarsus primus varus
C0265649|ICD9CM|PT|754.52|Metatarsus primus varus
C0265677|ICD9CM|AB|756.14|Hemivertebra
C0265677|ICD9CM|PT|756.14|Hemivertebra
C0265678|ICD9CM|PT|756.15|Fusion of spine (vertebra), congenital
C0265678|ICD9CM|AB|756.15|Congen fusion of spine
C0265706|ICD9CM|AB|756.73|Gastroschisis
C0265706|ICD9CM|PT|756.73|Gastroschisis
C0265830|ICD9CM|HT|746.0|Anomalies of pulmonary valve, congenital
C0265830|ICD9CM|PT|746.00|Congenital pulmonary valve anomaly, unspecified
C0265830|ICD9CM|AB|746.00|Pulmonary valve anom NOS
C0265970|ICD9CM|PT|692.75|Disseminated superficial actinic porokeratosis (DSAP)
C0265970|ICD9CM|AB|692.75|Dis sup actnc porokrtsis
C0265973|ICD9CM|AB|757.32|Vascular hamartomas
C0265973|ICD9CM|PT|757.32|Vascular hamartomas
C0266013|ICD9CM|PT|611.82|Hypoplasia of breast
C0266013|ICD9CM|AB|611.82|Hypoplasia of breast
C0266015|ICD9CM|PT|751.9|Unspecified anomaly of digestive system
C0266015|ICD9CM|AB|751.9|Anom digestive syst NOS
C0266021|ICD9CM|PT|750.8|Other specified anomalies of upper alimentary tract
C0266021|ICD9CM|AB|750.8|Upper GI anomaly NEC
C0266060|ICD9CM|PT|524.24|Open anterior occlusal relationship
C0266060|ICD9CM|AB|524.24|Open anterior occlusion
C0266071|ICD9CM|AB|524.35|Rotation of teeth
C0266071|ICD9CM|PT|524.35|Rotation of tooth/teeth
C0266094|ICD9CM|AB|744.81|Macrocheilia
C0266094|ICD9CM|PT|744.81|Macrocheilia
C0266095|ICD9CM|AB|744.82|Microcheilia
C0266095|ICD9CM|PT|744.82|Microcheilia
C0266118|ICD9CM|PT|750.23|Atresia, salivary duct
C0266118|ICD9CM|AB|750.23|Cong atresia, saliv duct
C0266384|ICD9CM|AB|752.31|Agenesis of uterus
C0266384|ICD9CM|PT|752.31|Agenesis of uterus
C0266385|ICD9CM|AB|752.36|Arcuate uterus
C0266385|ICD9CM|PT|752.36|Arcuate uterus
C0266387|ICD9CM|PT|752.34|Bicornuate uterus
C0266387|ICD9CM|AB|752.34|Bicornuate uterus
C0266389|ICD9CM|PT|752.33|Unicornuate uterus
C0266389|ICD9CM|AB|752.33|Unicornuate uterus
C0266399|ICD9CM|PT|752.32|Hypoplasia of uterus
C0266399|ICD9CM|AB|752.32|Hypoplasia of uterus
C0266404|ICD9CM|PT|752.43|Cervical agenesis
C0266404|ICD9CM|AB|752.43|Cervical agenesis
C0266436|ICD9CM|AB|752.63|Congenital chordee
C0266436|ICD9CM|PT|752.63|Congenital chordee
C0266521|ICD9CM|PT|374.43|Abnormal innervation syndrome of eyelid
C0266521|ICD9CM|AB|374.43|Abnorm innervation synd
C0266572|ICD9CM|PT|743.62|Congenital deformities of eyelids
C0266572|ICD9CM|AB|743.62|Congenital eyelid deform
C0266573|ICD9CM|AB|743.61|Congenital ptosis
C0266573|ICD9CM|PT|743.61|Congenital ptosis
C0266587|ICD9CM|PT|743.66|Specified congenital anomalies of orbit
C0266587|ICD9CM|AB|743.66|Spec anomaly of orbit
C0266589|ICD9CM|PT|744.3|Unspecified anomaly of ear
C0266589|ICD9CM|AB|744.3|Ear anomaly NOS
C0266592|ICD9CM|HT|744.0|Congenital anomalies of ear causing impairment of hearing
C0266592|ICD9CM|AB|744.00|Ear anom NOS/impair hear
C0266592|ICD9CM|PT|744.00|Unspecified anomaly of ear with impairment of hearing
C0266611|ICD9CM|AB|744.1|Accessory auricle
C0266611|ICD9CM|PT|744.1|Accessory auricle
C0266781|ICD9CM|PT|792.3|Nonspecific abnormal findings in amniotic fluid
C0266781|ICD9CM|AB|792.3|Abn find-amniotic fluid
C0266846|ICD9CM|PT|521.02|Dental caries extending into dentine
C0266846|ICD9CM|AB|521.02|Dental caries - dentine
C0266848|ICD9CM|PT|521.04|Arrested dental caries
C0266848|ICD9CM|AB|521.04|Dental caries - arrested
C0266853|ICD9CM|AB|521.01|Dental caries - enamel
C0266853|ICD9CM|PT|521.01|Dental caries limited to enamel
C0266878|ICD9CM|PT|521.42|Pathological resorption, external
C0266878|ICD9CM|AB|521.42|Path resorption-external
C0266909|ICD9CM|PT|522.7|Periapical abscess with sinus
C0266909|ICD9CM|AB|522.7|Periapical absc w sinus
C0266915|ICD9CM|PT|523.25|Gingival recession, generalized
C0266915|ICD9CM|AB|523.25|Gingival recess-general
C0266916|ICD9CM|PT|523.24|Gingival recession, localized
C0266916|ICD9CM|AB|523.24|Gingival recession-local
C0266929|ICD9CM|HT|523.4|Chronic periodontitis
C0266929|ICD9CM|PT|523.40|Chronic periodontitis, unspecified
C0266929|ICD9CM|AB|523.40|Chronc periodontitis NOS
C0266932|ICD9CM|HT|524.5|Dentofacial functional abnormalities
C0266932|ICD9CM|PT|524.50|Dentofacial functional abnormality, unspecified
C0266932|ICD9CM|AB|524.50|Dentofac funct abnor NOS
C0266933|ICD9CM|AB|524.51|Abnormal jaw closure
C0266933|ICD9CM|PT|524.51|Abnormal jaw closure
C0267071|ICD9CM|AB|787.22|Dysphagia, oropharyngeal
C0267071|ICD9CM|PT|787.22|Dysphagia, oropharyngeal phase
C0267092|ICD9CM|PT|456.1|Esophageal varices without mention of bleeding
C0267092|ICD9CM|AB|456.1|Esoph varices w/o bleed
C0267095|ICD9CM|AB|530.83|Esophageal leukoplakia
C0267095|ICD9CM|PT|530.83|Esophageal leukoplakia
C0267123|ICD9CM|PT|531.20|Acute gastric ulcer with hemorrhage and perforation, without mention of obstruction
C0267123|ICD9CM|AB|531.20|Ac stomac ulc w hem/perf
C0267124|ICD9CM|HT|531.3|Acute gastric ulcer without mention of hemorrhage or perforation
C0267125|ICD9CM|PT|531.30|Acute gastric ulcer without mention of hemorrhage or perforation, without mention of obstruction
C0267125|ICD9CM|AB|531.30|Acute stomach ulcer NOS
C0267136|ICD9CM|HT|531.7|Chronic gastric ulcer without mention of hemorrhage or perforation
C0267138|ICD9CM|PT|531.71|Chronic gastric ulcer without mention of hemorrhage or perforation, with obstruction
C0267138|ICD9CM|AB|531.71|Chr stomach ulc NOS-obst
C0267154|ICD9CM|HT|535.7|Eosinophilic gastritis
C0267166|ICD9CM|HT|535|Gastritis and duodenitis
C0267180|ICD9CM|PT|537.4|Fistula of stomach or duodenum
C0267180|ICD9CM|AB|537.4|Gastric/duodenal fistula
C0267183|ICD9CM|PT|537.6|Hourglass stricture or stenosis of stomach
C0267183|ICD9CM|AB|537.6|Hourglass stricture stom
C0267262|ICD9CM|PT|532.10|Acute duodenal ulcer with perforation, without mention of obstruction
C0267262|ICD9CM|AB|532.10|Ac duodenal ulcer w perf
C0267282|ICD9CM|HT|532.7|Chronic duodenal ulcer without mention of hemorrhage or perforation
C0267288|ICD9CM|PT|533.00|Acute peptic ulcer of unspecified site with hemorrhage, without mention of obstruction
C0267288|ICD9CM|HT|533.0|Acute peptic ulcer of unspecified site with hemorrhage
C0267288|ICD9CM|AB|533.00|Ac peptic ulcer w hemorr
C0267291|ICD9CM|HT|533.1|Acute peptic ulcer of unspecified site with perforation
C0267294|ICD9CM|HT|533.2|Acute peptic ulcer of unspecified site with hemorrhage and perforation
C0267298|ICD9CM|PT|533.30|Acute peptic ulcer of unspecified site without mention of hemorrhage and perforation, without mention of obstruction
C0267298|ICD9CM|AB|533.30|Acute peptic ulcer NOS
C0267326|ICD9CM|PT|534.30|Acute gastrojejunal ulcer without mention of hemorrhage or perforation, without mention of obstruction
C0267326|ICD9CM|AB|534.30|Ac marginal ulcer NOS
C0267347|ICD9CM|PT|534.70|Chronic gastrojejunal ulcer without mention of hemorrhage or perforation, without mention of obstruction
C0267347|ICD9CM|AB|534.70|Chr marginal ulcer NOS
C0267367|ICD9CM|PT|569.84|Angiodysplasia of intestine (without mention of hemorrhage)
C0267367|ICD9CM|AB|569.84|Angio intes w/o hmrhg
C0267383|ICD9CM|PT|555.2|Regional enteritis of small intestine with large intestine
C0267383|ICD9CM|AB|555.2|Reg enterit sm/lg intest
C0267388|ICD9CM|PT|556.0|Ulcerative (chronic) enterocolitis
C0267388|ICD9CM|AB|556.0|Ulcerative enterocolitis
C0267389|ICD9CM|PT|556.1|Ulcerative (chronic) ileocolitis
C0267389|ICD9CM|AB|556.1|Ulcerative ileocolitis
C0267390|ICD9CM|PT|556.3|Ulcerative (chronic) proctosigmoiditis
C0267390|ICD9CM|AB|556.3|Ulcertve prctosigmoidtis
C0267392|ICD9CM|PT|556.4|Pseudopolyposis of colon
C0267392|ICD9CM|AB|556.4|Pseudopolyposis colon
C0267448|ICD9CM|PT|558.42|Eosinophilic colitis
C0267448|ICD9CM|AB|558.42|Eosinophilic colitis
C0267498|ICD9CM|HT|562.0|Diverticula of small intestine
C0267567|ICD9CM|PT|566|Abscess of anal and rectal regions
C0267567|ICD9CM|AB|566|Anal & rectal abscess
C0267667|ICD9CM|PT|551.9|Hernia of unspecified site, with gangrene
C0267667|ICD9CM|AB|551.9|Hernia, site NOS w gangr
C0267751|ICD9CM|PT|567.21|Peritonitis (acute) generalized
C0267751|ICD9CM|AB|567.21|Peritonitis (acute) gen
C0267756|ICD9CM|AB|567.22|Peritoneal abscess
C0267756|ICD9CM|PT|567.22|Peritoneal abscess
C0267768|ICD9CM|AB|567.81|Choleperitonitis
C0267768|ICD9CM|PT|567.81|Choleperitonitis
C0267770|ICD9CM|AB|567.82|Sclerosing mesenteritis
C0267770|ICD9CM|PT|567.82|Sclerosing mesenteritis
C0267981|ICD9CM|PT|262|Other severe protein-calorie malnutrition
C0267981|ICD9CM|AB|262|Oth severe malnutrition
C0267994|ICD9CM|HT|276|Disorders of fluid, electrolyte, and acid-base balance
C0268301|ICD9CM|PT|259.52|Partial androgen insensitivity
C0268301|ICD9CM|AB|259.52|Part androgen insnsitvty
C0268329|ICD9CM|HT|277|Other and unspecified disorders of metabolism
C0268512|ICD9CM|PT|270.5|Disturbances of histidine metabolism
C0268512|ICD9CM|AB|270.5|Dis histidine metabolism
C0268613|ICD9CM|PT|270.4|Disturbances of sulphur-bearing amino-acid metabolism
C0268613|ICD9CM|AB|270.4|Sulph amino-acid met dis
C0268641|ICD9CM|PT|270.0|Disturbances of amino-acid transport
C0268641|ICD9CM|AB|270.0|Amino-acid transport dis
C0268701|ICD9CM|PT|593.9|Unspecified disorder of kidney and ureter
C0268701|ICD9CM|AB|593.9|Renal & ureteral dis NOS
C0268790|ICD9CM|AB|593.81|Renal vascular disorder
C0268790|ICD9CM|PT|593.81|Vascular disorders of kidney
C0268792|ICD9CM|PT|445.81|Atheroembolism of kidney
C0268792|ICD9CM|AB|445.81|Atheroembolism, kidney
C0268799|ICD9CM|AB|593.2|Cyst of kidney, acquired
C0268799|ICD9CM|PT|593.2|Cyst of kidney, acquired
C0268882|ICD9CM|PT|601.8|Other specified inflammatory diseases of prostate
C0268882|ICD9CM|AB|601.8|Prostatic inflam dis NEC
C0269032|ICD9CM|PT|614.5|Acute or unspecified pelvic peritonitis, female
C0269032|ICD9CM|AB|614.5|Ac pelv peritonitis-fem
C0269047|ICD9CM|PT|615.9|Unspecified inflammatory disease of uterus
C0269047|ICD9CM|AB|615.9|Uterine inflam dis NOS
C0269084|ICD9CM|PT|625.71|Vulvar vestibulitis
C0269084|ICD9CM|AB|625.71|Vulvar vestibulitis
C0269131|ICD9CM|PT|619.9|Unspecified fistula involving female genital tract
C0269131|ICD9CM|AB|619.9|Fem genital fistula NOS
C0269194|ICD9CM|AB|622.2|Leukoplakia of cervix
C0269194|ICD9CM|PT|622.2|Leukoplakia of cervix (uteri)
C0269223|ICD9CM|PT|624.4|Old laceration or scarring of vulva
C0269223|ICD9CM|AB|624.4|Old laceration of vulva
C0269226|ICD9CM|HT|346.4|Menstrual migraine
C0269294|ICD9CM|PT|639.0|Genital tract and pelvic infection following abortion or ectopic and molar pregnancies
C0269294|ICD9CM|AB|639.0|Postabortion gu infect
C0269403|ICD9CM|HT|634.2|Spontaneous abortion complicated by damage to pelvic organs or tissues
C0269403|ICD9CM|PT|634.20|Spontaneous abortion, complicated by damage to pelvic organs or tissues, unspecified
C0269403|ICD9CM|AB|634.20|Spon ab w pel damag-unsp
C0269441|ICD9CM|HT|635.8|Legally induced abortion with unspecified complication
C0269441|ICD9CM|PT|635.80|Legally induced abortion, with unspecified complication, unspecified
C0269441|ICD9CM|AB|635.80|Leg ab w compl NOS-unsp
C0269450|ICD9CM|PT|635.10|Legally induced abortion, complicated by delayed or excessive hemorrhage, unspecified
C0269450|ICD9CM|HT|635.1|Legally induced abortion complicated by delayed or excessive hemorrhage
C0269450|ICD9CM|AB|635.10|Legal abor w hemorr-unsp
C0269469|ICD9CM|HT|635.3|Legally induced abortion complicated by renal failure
C0269469|ICD9CM|PT|635.30|Legally induced abortion, complicated by renal failure,unspecified
C0269469|ICD9CM|AB|635.30|Leg abor w ren fail-unsp
C0269474|ICD9CM|HT|635.4|Legally induced abortion complicated by metabolic disorder
C0269474|ICD9CM|PT|635.40|Legally induced abortion, complicated by metabolic disorder, unspecified
C0269474|ICD9CM|AB|635.40|Leg ab w metab dis-unsp
C0269476|ICD9CM|HT|635.5|Legally induced abortion complicated by shock
C0269476|ICD9CM|PT|635.50|Legally induced abortion, complicated by shock, unspecified
C0269476|ICD9CM|AB|635.50|Legal abort w shock-unsp
C0269479|ICD9CM|HT|635.6|Legally induced abortion complicated by embolism
C0269479|ICD9CM|PT|635.60|Legally induced abortion, complicated by embolism, unspecified
C0269479|ICD9CM|AB|635.60|Legal abort w embol-unsp
C0269496|ICD9CM|HT|636.8|Illegally induced abortion with unspecified complication
C0269496|ICD9CM|PT|636.80|Illegally induced abortion, with unspecified complication, unspecified
C0269496|ICD9CM|AB|636.80|Illg ab w compl NOS-unsp
C0269505|ICD9CM|PT|636.10|Illegally induced abortion, complicated by delayed or excessive hemorrhage, unspecified
C0269505|ICD9CM|HT|636.1|Illegally induced abortion complicated by delayed or excessive hemorrhage
C0269505|ICD9CM|AB|636.10|Illeg ab w hemorr-unspec
C0269509|ICD9CM|HT|636.2|Illegally induced abortion complicated by damage to pelvic organs or tissue
C0269509|ICD9CM|PT|636.20|Illegally induced abortion, complicated by damage to pelvic organs or tissues, unspecified
C0269509|ICD9CM|AB|636.20|Illeg ab w pel damg-unsp
C0269524|ICD9CM|HT|636.3|Illegally induced abortion complicated by renal failure
C0269524|ICD9CM|PT|636.30|Illegally induced abortion, complicated by renal failure, unspecified
C0269524|ICD9CM|AB|636.30|Illeg ab w ren fail-unsp
C0269529|ICD9CM|HT|636.4|Illegally induced abortion complicated by metabolic disorder
C0269529|ICD9CM|PT|636.40|Illegally induced abortion, complicated by metabolic disorder, unspecified
C0269529|ICD9CM|AB|636.40|Illeg ab w met dis-unsp
C0269531|ICD9CM|HT|636.5|Illegally induced abortion complicated by shock
C0269531|ICD9CM|PT|636.50|Illegally induced abortion, complicated by shock, unspecified
C0269531|ICD9CM|AB|636.50|Illeg abort w shock-unsp
C0269534|ICD9CM|HT|636.6|Illegally induced abortion complicated by embolism
C0269534|ICD9CM|PT|636.60|Illegally induced abortion, complicated by embolism, unspecified
C0269534|ICD9CM|AB|636.60|Illeg ab w embolism-unsp
C0269549|ICD9CM|PT|638.9|Failed attempted abortion without mention of complication
C0269549|ICD9CM|AB|638.9|Attempted abort uncompl
C0269561|ICD9CM|PT|638.2|Failed attempted abortion complicated by damage to pelvic organs or tissues
C0269561|ICD9CM|AB|638.2|Attem abort w pelv damag
C0269599|ICD9CM|PT|640.93|Unspecified hemorrhage in early pregnancy, antepartum condition or complication
C0269599|ICD9CM|AB|640.93|Hem early preg-antepart
C0269607|ICD9CM|PT|640.83|Other specified hemorrhage in early pregnancy, antepartum condition or complication
C0269607|ICD9CM|AB|640.83|Hem early pg NEC-antepar
C0269608|ICD9CM|HT|641.9|Unspecified antepartum hemorrhage
C0269608|ICD9CM|PT|641.93|Unspecified antepartum hemorrhage, antepartum condition or complication
C0269608|ICD9CM|AB|641.93|Antepart hem NOS-antepar
C0269658|ICD9CM|HT|642.4|Mild or unspecified pre-eclampsia
C0269661|ICD9CM|HT|643.9|Unspecified vomiting of pregnancy
C0269673|ICD9CM|HT|646.2|Unspecified renal disease in pregnancy, without mention of hypertension
C0269683|ICD9CM|HT|648.1|Thyroid dysfunction complicating pregnancy, childbirth, or the puerperium
C0269684|ICD9CM|PT|648.20|Anemia of mother, unspecified as to episode of care or not applicable
C0269684|ICD9CM|HT|648.2|Anemia complicating pregnancy, childbirth, or the puerperium
C0269684|ICD9CM|AB|648.20|Anemia in preg-unspec
C0269685|ICD9CM|HT|648.3|Drug dependence complicating pregnancy, childbirth, or the puerperium
C0269685|ICD9CM|PT|648.30|Drug dependence of mother, unspecified as to episode of care or not applicable
C0269685|ICD9CM|AB|648.30|Drug depend preg-unspec
C0269709|ICD9CM|HT|652.7|Prolapsed arm of fetus
C0269713|ICD9CM|HT|653.0|Major abnormality of bony pelvis, not further specified, in pregnancy, labor, and delivery
C0269792|ICD9CM|HT|656.4|Intrauterine death affecting management of mother
C0269807|ICD9CM|HT|659.0|Failed mechanical induction of labor
C0269815|ICD9CM|HT|669.9|Unspecified complication of labor and delivery
C0269825|ICD9CM|HT|660.4|Shoulder (girdle) dystocia during labor and delivery
C0269852|ICD9CM|PT|663.53|Vasa previa complicating labor and delivery, antepartum condition or complication
C0269852|ICD9CM|AB|663.53|Vasa previa-antepartum
C0269858|ICD9CM|HT|665.9|Unspecified obstetrical trauma
C0269859|ICD9CM|HT|664.4|Unspecified perineal laceration during delivery
C0269859|ICD9CM|PT|664.41|Unspecified perineal laceration, delivered, with or without mention of antepartum condition
C0269859|ICD9CM|AB|664.41|Ob perineal lac NOS-del
C0269863|ICD9CM|HT|664.0|First-degree perineal laceration during delivery
C0269870|ICD9CM|HT|664.1|Second-degree perineal laceration during delivery
C0269870|ICD9CM|PT|664.11|Second-degree perineal laceration, delivered, with or without mention of antepartum condition
C0269870|ICD9CM|AB|664.11|Del w 2 deg lacerat-del
C0269874|ICD9CM|HT|664.2|Third-degree perineal laceration during delivery
C0269874|ICD9CM|PT|664.21|Third-degree perineal laceration, delivered, with or without mention of antepartum condition
C0269874|ICD9CM|AB|664.21|Del w 3 deg lacerat-del
C0269891|ICD9CM|HT|665.6|Obstetrical damage to pelvic joints and ligaments
C0269891|ICD9CM|PT|665.61|Damage to pelvic joints and ligaments, delivered, with or without mention of antepartum condition
C0269891|ICD9CM|AB|665.61|Damage to pelvic jt-del
C0269895|ICD9CM|PT|665.71|Pelvic hematoma, delivered, with or without mention of antepartum condition
C0269895|ICD9CM|HT|665.7|Obstetrical pelvic hematoma
C0269895|ICD9CM|AB|665.71|Ob pelvic hematoma-deliv
C0269898|ICD9CM|HT|666.0|Third-stage postpartum hemorrhage
C0269898|ICD9CM|PT|666.04|Third-stage postpartum hemorrhage, postpartum condition or complication
C0269898|ICD9CM|AB|666.04|Third-stage hem-postpart
C0269905|ICD9CM|HT|667.0|Retained placenta without hemorrhage
C0269916|ICD9CM|HT|668.1|Cardiac complications of anesthesia or other sedation in labor and delivery
C0269930|ICD9CM|HT|669.7|Cesarean delivery, without mention of indication
C0269932|ICD9CM|HT|670.1|Puerperal endometritis
C0269936|ICD9CM|HT|670.2|Puerperal sepsis
C0269945|ICD9CM|HT|671|Venous complications in pregnancy and the puerperium
C0269945|ICD9CM|HT|671.9|Unspecified venous complication in pregnancy and the puerperium
C0269945|ICD9CM|PT|671.90|Unspecified venous complication of pregnancy and the puerperium, unspecified as to episode of care or not applicable
C0269945|ICD9CM|AB|671.90|Ven compl preg NOS-unsp
C0269951|ICD9CM|HT|671.2|Superficial thrombophlebitis in pregnancy and the puerperium
C0269951|ICD9CM|PT|671.20|Superficial thrombophlebitis complicating pregnancy and the puerperium, unspecified as to episode of care or not applicable
C0269951|ICD9CM|AB|671.20|Thrombophleb preg-unspec
C0269959|ICD9CM|HT|673.3|Obstetrical pyemic and septic embolism
C0269959|ICD9CM|PT|673.30|Obstetrical pyemic and septic embolism, unspecified as to episode of care or not applicable
C0269959|ICD9CM|AB|673.30|Ob pyemic embol-unspec
C0269979|ICD9CM|HT|675.0|Infections of nipple associated with childbirth
C0269981|ICD9CM|HT|675.1|Abscess of breast associated with childbirth
C0269993|ICD9CM|HT|676.5|Suppressed lactation
C0269993|ICD9CM|PT|676.50|Suppressed lactation, unspecified as to episode of care or not applicable
C0269993|ICD9CM|AB|676.50|Suppr lactation-unspec
C0269995|ICD9CM|HT|676.6|Galactorrhea
C0269995|ICD9CM|PT|676.60|Galactorrhea associated with childbirth, unspecified as to episode of care or not applicable
C0269995|ICD9CM|AB|676.60|Galactorrhea preg-unspec
C0270025|ICD9CM|HT|762|Fetus or newborn affected by complications of placenta, cord, and membranes
C0270067|ICD9CM|HT|763.8|Other specified complications of labor and delivery affecting fetus or newborn
C0270067|ICD9CM|PT|763.89|Other specified complications of labor and delivery affecting fetus or newborn
C0270067|ICD9CM|AB|763.89|Compl del NEC aff NB
C0270075|ICD9CM|PT|779.9|Unspecified condition originating in the perinatal period
C0270075|ICD9CM|AB|779.9|Perinatal condition NOS
C0270078|ICD9CM|HT|765.0|Extreme immaturity
C0270089|ICD9CM|HT|767.1|Injuries to scalp due to birth trauma
C0270092|ICD9CM|PT|767.11|Epicranial subaponeurotic hemorrhage (massive)
C0270092|ICD9CM|AB|767.11|Epicranial subapo hemorr
C0270094|ICD9CM|PT|767.2|Fracture of clavicle due to birth trauma
C0270094|ICD9CM|AB|767.2|Clavicle fx at birth
C0270103|ICD9CM|PT|767.5|Facial nerve injury due to birth trauma
C0270103|ICD9CM|AB|767.5|Facial nerve inj-birth
C0270105|ICD9CM|PT|767.6|Injury to brachial plexus due to birth trauma
C0270105|ICD9CM|AB|767.6|Brach plexus inj-birth
C0270124|ICD9CM|AB|768.4|Fetal distress NOS
C0270124|ICD9CM|PT|768.4|Fetal distress, unspecified as to time of onset, in liveborn infant
C0270131|ICD9CM|PT|768.0|Fetal death from asphyxia or anoxia before onset of labor or at unspecified time
C0270131|ICD9CM|AB|768.0|Fetal death-anoxia NOS
C0270146|ICD9CM|PT|770.9|Unspecified respiratory condition of fetus and newborn
C0270146|ICD9CM|AB|770.9|NB respiratory cond NOS
C0270148|ICD9CM|PT|770.83|Cyanotic attacks of newborn
C0270148|ICD9CM|AB|770.83|Cyanotic attack, newborn
C0270163|ICD9CM|AB|770.4|Primary atelectasis
C0270163|ICD9CM|PT|770.4|Primary atelectasis
C0270183|ICD9CM|PT|772.9|Unspecified hemorrhage of newborn
C0270183|ICD9CM|AB|772.9|Neonatal hemorrhage NOS
C0270191|ICD9CM|HT|772.1|Intraventricular hemorrhage of fetus or newborn
C0270202|ICD9CM|PT|773.1|Hemolytic disease of fetus or newborn due to ABO isoimmunization
C0270202|ICD9CM|AB|773.1|NB hemolyt dis-abo isoim
C0270204|ICD9CM|PT|773.4|Kernicterus of fetus or newborn due to isoimmunization
C0270204|ICD9CM|AB|773.4|NB kernicterus:isoimmun
C0270206|ICD9CM|PT|774.6|Unspecified fetal and neonatal jaundice
C0270206|ICD9CM|AB|774.6|Fetal/neonatal jaund NOS
C0270221|ICD9CM|PT|775.0|Syndrome of "infant of a diabetic mother"
C0270221|ICD9CM|AB|775.0|Infant diabet mother syn
C0270246|ICD9CM|PT|777.1|Meconium obstruction in fetus or newborn
C0270246|ICD9CM|AB|777.1|Meconium obstruction
C0270249|ICD9CM|PT|777.3|Hematemesis and melena of newborn due to swallowed maternal blood
C0270249|ICD9CM|AB|777.3|Swallowed blood syndrome
C0270275|ICD9CM|PT|779.4|Drug reactions and intoxications specific to newborn
C0270275|ICD9CM|AB|779.4|NB drug reaction/intoxic
C0270307|ICD9CM|AB|313.0|Overanxious disorder
C0270307|ICD9CM|PT|313.0|Overanxious disorder specific to childhood and adolescence
C0270327|ICD9CM|AB|788.36|Nocturnal enuresis
C0270327|ICD9CM|PT|788.36|Nocturnal enuresis
C0270381|ICD9CM|PT|295.91|Unspecified schizophrenia, subchronic
C0270381|ICD9CM|AB|295.91|Schizophrenia NOS-subchr
C0270384|ICD9CM|PT|295.95|Unspecified schizophrenia, in remission
C0270384|ICD9CM|AB|295.95|Schizophrenia NOS-remiss
C0270390|ICD9CM|PT|295.25|Catatonic type schizophrenia, in remission
C0270390|ICD9CM|AB|295.25|Catatonia-remission
C0270395|ICD9CM|PT|295.15|Disorganized type schizophrenia, in remission
C0270395|ICD9CM|AB|295.15|Hebephrenia-remission
C0270398|ICD9CM|PT|295.32|Paranoid type schizophrenia, chronic
C0270398|ICD9CM|AB|295.32|Paranoid schizo-chronic
C0270403|ICD9CM|PT|295.92|Unspecified schizophrenia, chronic
C0270403|ICD9CM|AB|295.92|Schizophrenia NOS-chr
C0270406|ICD9CM|PT|295.61|Schizophrenic disorders, residual type, subchronic
C0270406|ICD9CM|AB|295.61|Schizoph dis resid-subch
C0270408|ICD9CM|PT|295.62|Schizophrenic disorders, residual type, chronic
C0270408|ICD9CM|AB|295.62|Schizophr dis resid-chr
C0270434|ICD9CM|PT|296.66|Bipolar I disorder, most recent episode (or current) mixed, in full remission
C0270434|ICD9CM|AB|296.66|Bipol I cur mixed remiss
C0270543|ICD9CM|PT|327.10|Organic hypersomnia, unspecified
C0270543|ICD9CM|AB|327.10|Organic hypersomnia NOS
C0270549|ICD9CM|PT|300.02|Generalized anxiety disorder
C0270549|ICD9CM|AB|300.02|Generalized anxiety dis
C0270627|ICD9CM|HT|341.2|Acute (transverse) myelitis
C0270627|ICD9CM|PT|341.20|Acute (transverse) myelitis NOS
C0270627|ICD9CM|AB|341.20|Acute myelitis NOS
C0270742|ICD9CM|PT|333.71|Athetoid cerebral palsy
C0270742|ICD9CM|AB|333.71|Athetoid cerebral palsy
C0270799|ICD9CM|PT|344.60|Cauda equina syndrome without mention of neurogenic bladder
C0270799|ICD9CM|AB|344.60|Cauda equina synd NOS
C0270805|ICD9CM|AB|343.1|Congenital hemiplegia
C0270805|ICD9CM|PT|343.1|Congenital hemiplegia
C0270823|ICD9CM|AB|345.2|Petit mal status
C0270823|ICD9CM|PT|345.2|Petit mal status
C0270862|ICD9CM|HT|346.3|Hemiplegic migraine
C0270890|ICD9CM|HT|353|Nerve root and plexus disorders
C0270890|ICD9CM|PT|353.9|Unspecified nerve root and plexus disorder
C0270890|ICD9CM|AB|353.9|Nerv root/plexus dis NOS
C0270909|ICD9CM|PT|355.3|Lesion of lateral popliteal nerve
C0270909|ICD9CM|AB|355.3|Lat popliteal nerve les
C0270932|ICD9CM|PT|357.3|Polyneuropathy in malignant disease
C0270932|ICD9CM|AB|357.3|Neuropathy in malig dis
C0270942|ICD9CM|PT|358.01|Myasthenia gravis with (acute) exacerbation
C0270942|ICD9CM|AB|358.01|Myasthna gravs w ac exac
C0271001|ICD9CM|AB|360.23|Siderosis
C0271001|ICD9CM|PT|360.23|Siderosis of globe
C0271008|ICD9CM|HT|360.5|Retained (old) intraocular foreign body, magnetic
C0271008|ICD9CM|PT|360.50|Foreign body, magnetic, intraocular, unspecified
C0271008|ICD9CM|AB|360.50|Old magnet fb, eye NOS
C0271015|ICD9CM|HT|360.6|Retained (old) intraocular foreign body, nonmagnetic
C0271083|ICD9CM|PT|362.51|Nonexudative senile macular degeneration
C0271083|ICD9CM|AB|362.51|Nonexudat macular degen
C0271084|ICD9CM|PT|362.52|Exudative senile macular degeneration
C0271084|ICD9CM|AB|362.52|Exudative macular degen
C0271086|ICD9CM|AB|362.55|Toxic maculopathy
C0271086|ICD9CM|PT|362.55|Toxic maculopathy
C0271111|ICD9CM|AB|364.51|Progressive iris atrophy
C0271111|ICD9CM|PT|364.51|Essential or progressive iris atrophy
C0271128|ICD9CM|PT|364.61|Implantation cysts of iris, ciliary body, and anterior chamber
C0271128|ICD9CM|AB|364.61|Implantation cysts
C0271142|ICD9CM|HT|365.5|Glaucoma associated with disorders of the lens
C0271166|ICD9CM|AB|366.16|Senile nuclear cataract
C0271166|ICD9CM|PT|366.16|Senile nuclear sclerosis
C0271172|ICD9CM|PT|366.33|Cataract with neovascularization
C0271172|ICD9CM|AB|366.33|Cataract w neovasculizat
C0271202|ICD9CM|AB|368.46|Homonymous hemianopsia
C0271202|ICD9CM|PT|368.46|Homonymous bilateral field defects
C0271207|ICD9CM|AB|368.47|Heteronymous hemianopsia
C0271207|ICD9CM|PT|368.47|Heteronymous bilateral field defects
C0271220|ICD9CM|PT|369.04|Better eye: near-total vision impairment; lesser eye: near-total vision impairment
C0271220|ICD9CM|AB|369.04|Near-tot impair-both eye
C0271224|ICD9CM|PT|369.08|Better eye: profound vision impairment; lesser eye: profound vision impairment
C0271224|ICD9CM|AB|369.08|Profound impair both eye
C0271225|ICD9CM|AB|369.10|Blindness/low vision
C0271225|ICD9CM|PT|369.10|Moderate or severe impairment, better eye, impairment level not further specified
C0271234|ICD9CM|PT|369.20|Moderate or severe impairment, both eyes, impairment level not further specified
C0271234|ICD9CM|AB|369.20|Low vision, 2 eyes NOS
C0271236|ICD9CM|PT|369.22|Better eye: severe vision impairment; lesser eye: severe vision impairment
C0271236|ICD9CM|AB|369.22|Severe impair-both eyes
C0271239|ICD9CM|PT|369.25|Better eye: moderate vision impairment; lesser eye: moderate vision impairment
C0271239|ICD9CM|AB|369.25|Moderate impair-both eye
C0271275|ICD9CM|AB|371.04|Adherent leucoma
C0271275|ICD9CM|PT|371.04|Adherent leucoma
C0271311|ICD9CM|PT|374.05|Trichiasis of eyelid without entropion
C0271311|ICD9CM|AB|374.05|Trichiasis w/o entropion
C0271342|ICD9CM|PT|377.14|Glaucomatous atrophy [cupping] of optic disc
C0271342|ICD9CM|AB|377.14|Cupping of optic disc
C0271370|ICD9CM|PT|378.51|Third or oculomotor nerve palsy, partial
C0271370|ICD9CM|AB|378.51|Partial third nerv palsy
C0271371|ICD9CM|AB|378.52|Total third nerve palsy
C0271371|ICD9CM|PT|378.52|Third or oculomotor nerve palsy, total
C0271375|ICD9CM|PT|378.53|Fourth or trochlear nerve palsy
C0271375|ICD9CM|AB|378.53|Fourth nerve palsy
C0271384|ICD9CM|PT|379.53|Visual deprivation nystagmus
C0271384|ICD9CM|AB|379.53|Visual deprivatn nystagm
C0271411|ICD9CM|PT|388.72|Referred otogenic pain
C0271411|ICD9CM|AB|388.72|Referred pain of ear
C0271413|ICD9CM|PT|380.31|Hematoma of auricle or pinna
C0271413|ICD9CM|AB|380.31|Hematoma auricle/pinna
C0271431|ICD9CM|HT|382.0|Acute suppurative otitis media
C0271432|ICD9CM|HT|381.0|Acute nonsuppurative otitis media
C0271432|ICD9CM|PT|381.00|Acute nonsuppurative otitis media, unspecified
C0271432|ICD9CM|AB|381.00|Ac nonsup otitis med NOS
C0271446|ICD9CM|AB|381.4|Nonsupp otitis media NOS
C0271446|ICD9CM|PT|381.4|Nonsuppurative otitis media, not specified as acute or chronic
C0271454|ICD9CM|PT|382.3|Unspecified chronic suppurative otitis media
C0271454|ICD9CM|AB|382.3|Chr sup otitis media NOS
C0271468|ICD9CM|PT|381.81|Dysfunction of Eustachian tube
C0271468|ICD9CM|PT|381.9|Unspecified Eustachian tube disorder
C0271468|ICD9CM|AB|381.9|Eustachian tube dis NOS
C0271468|ICD9CM|AB|381.81|Dysfunct eustachian tube
C0271471|ICD9CM|PT|381.62|Intrinsic cartilagenous obstruction of Eustachian tube
C0271471|ICD9CM|AB|381.62|Intrinsic eustach obstr
C0271510|ICD9CM|AB|388.44|Auditory recruitment
C0271510|ICD9CM|PT|388.44|Auditory recruitment
C0271635|ICD9CM|HT|250.0|Diabetes mellitus without mention of complication
C0271640|ICD9CM|HT|249|Secondary diabetes mellitus
C0271680|ICD9CM|PT|357.2|Polyneuropathy in diabetes
C0271680|ICD9CM|AB|357.2|Neuropathy in diabetes
C0271761|ICD9CM|PT|241.1|Nontoxic multinodular goiter
C0271761|ICD9CM|AB|241.1|Nontox multinodul goiter
C0271763|ICD9CM|HT|242.9|Thyrotoxicosis without mention of goiter or other cause
C0271847|ICD9CM|PT|588.81|Secondary hyperparathyroidism (of renal origin)
C0271847|ICD9CM|AB|588.81|Sec hyperparathyrd-renal
C0271930|ICD9CM|AB|648.23|Anemia-antepartum
C0271930|ICD9CM|PT|648.23|Anemia of mother, antepartum condition or complication
C0271985|ICD9CM|AB|282.45|Delta-beta thalassemia
C0271985|ICD9CM|PT|282.45|Delta-beta thalassemia
C0272078|ICD9CM|PT|282.61|Hb-SS disease without crisis
C0272078|ICD9CM|AB|282.61|Hb-SS disease w/o crisis
C0272126|ICD9CM|AB|287.32|Evans' syndrome
C0272126|ICD9CM|PT|287.32|Evans' syndrome
C0272153|ICD9CM|AB|776.4|Polycythemia neonatorum
C0272153|ICD9CM|PT|776.4|Polycythemia neonatorum
C0272178|ICD9CM|PT|288.03|Drug induced neutropenia
C0272178|ICD9CM|AB|288.03|Drug induced neutropenia
C0272181|ICD9CM|PT|288.04|Neutropenia due to infection
C0272181|ICD9CM|AB|288.04|Neutropenia d/t infectn
C0272285|ICD9CM|PT|289.84|Heparin-induced thrombocytopenia (HIT)
C0272285|ICD9CM|AB|289.84|Heparin-indu thrombocyto
C0272422|ICD9CM|PT|959.09|Injury of face and neck
C0272422|ICD9CM|AB|959.09|Face & neck injury
C0272443|ICD9CM|PT|959.3|Elbow, forearm, and wrist injury
C0272443|ICD9CM|AB|959.3|Elb/forearm/wrst inj NOS
C0272468|ICD9CM|PT|802.22|Closed fracture of mandible, subcondylar
C0272468|ICD9CM|AB|802.22|Subcondylar fx mandib-cl
C0272469|ICD9CM|PT|802.24|Closed fracture of mandible, ramus, unspecified
C0272469|ICD9CM|AB|802.24|Fx ramus NOS-closed
C0272471|ICD9CM|PT|802.32|Open fracture of mandible, subcondylar
C0272471|ICD9CM|AB|802.32|Subcondyl fx mandib-open
C0272472|ICD9CM|PT|802.34|Open fracture of mandible, ramus, unspecified
C0272472|ICD9CM|AB|802.34|Fx ramus NOS-open
C0272576|ICD9CM|PT|808.8|Closed unspecified fracture of pelvis
C0272576|ICD9CM|AB|808.8|Pelvic fracture NOS-clos
C0272577|ICD9CM|PT|808.9|Open unspecified fracture of pelvis
C0272577|ICD9CM|AB|808.9|Pelvic fracture NOS-open
C0272580|ICD9CM|PT|808.43|Multiple closed pelvic fractures with disruption of pelvic circle
C0272580|ICD9CM|AB|808.43|Pelv fx-clos/pelv disrup
C0272582|ICD9CM|PT|808.53|Multiple open pelvic fractures with disruption of pelvic circle
C0272582|ICD9CM|AB|808.53|Pelv fx-open/pelv disrup
C0272609|ICD9CM|PT|812.20|Closed fracture of unspecified part of humerus
C0272609|ICD9CM|AB|812.20|Fx humerus NOS-closed
C0272610|ICD9CM|PT|812.30|Open fracture of unspecified part of humerus
C0272610|ICD9CM|AB|812.30|Fx humerus NOS-open
C0272638|ICD9CM|PT|813.21|Closed fracture of shaft of radius (alone)
C0272638|ICD9CM|AB|813.21|Fx radius shaft-closed
C0272641|ICD9CM|PT|813.31|Open fracture of shaft of radius (alone)
C0272641|ICD9CM|AB|813.31|Fx radius shaft-open
C0272647|ICD9CM|PT|813.43|Closed fracture of distal end of ulna (alone)
C0272647|ICD9CM|AB|813.43|Fx distal ulna-closed
C0272665|ICD9CM|PT|814.03|Closed fracture of triquetral [cuneiform] bone of wrist
C0272665|ICD9CM|AB|814.03|Fx triquetral, wrist-cl
C0272666|ICD9CM|PT|814.05|Closed fracture of trapezium bone [larger multangular] of wrist
C0272666|ICD9CM|AB|814.05|Fx trapezium bone-closed
C0272668|ICD9CM|PT|814.07|Closed fracture of capitate bone [os magnum] of wrist
C0272668|ICD9CM|AB|814.07|Fx capitate bone-closed
C0272669|ICD9CM|PT|814.08|Closed fracture of hamate [unciform] bone of wrist
C0272669|ICD9CM|AB|814.08|Fx hamate bone-closed
C0272672|ICD9CM|PT|814.13|Open fracture of triquetral [cuneiform] bone of wrist
C0272672|ICD9CM|AB|814.13|Fx triquetral, wrist-opn
C0272673|ICD9CM|PT|814.15|Open fracture of trapezium bone [larger multangular] of wrist
C0272673|ICD9CM|AB|814.15|Fx trapezium bone-open
C0272675|ICD9CM|PT|814.17|Open fracture of capitate bone [os magnum] of wrist
C0272675|ICD9CM|AB|814.17|Fx capitate bone-open
C0272676|ICD9CM|PT|814.18|Open fracture of hamate [unciform] bone of wrist
C0272676|ICD9CM|AB|814.18|Fx hamate bone-open
C0272677|ICD9CM|HT|815|Fracture of metacarpal bone(s)
C0272684|ICD9CM|PT|815.01|Closed fracture of base of thumb [first] metacarpal
C0272684|ICD9CM|AB|815.01|Fx 1st metacarp base-cl
C0272686|ICD9CM|PT|815.02|Closed fracture of base of other metacarpal bone(s)
C0272686|ICD9CM|AB|815.02|Fx metacarp base NEC-cl
C0272687|ICD9CM|PT|815.03|Closed fracture of shaft of metacarpal bone(s)
C0272687|ICD9CM|AB|815.03|Fx metacarpal shaft-clos
C0272688|ICD9CM|PT|815.04|Closed fracture of neck of metacarpal bone(s)
C0272688|ICD9CM|AB|815.04|Fx metacarpal neck-close
C0272689|ICD9CM|PT|815.11|Open fracture of base of thumb [first] metacarpal
C0272689|ICD9CM|AB|815.11|Fx 1st metacarp base-opn
C0272691|ICD9CM|PT|815.12|Open fracture of base of other metacarpal bone(s)
C0272691|ICD9CM|AB|815.12|Fx metacarp base NEC-opn
C0272692|ICD9CM|PT|815.13|Open fracture of shaft of metacarpal bone(s)
C0272692|ICD9CM|AB|815.13|Fx metacarpal shaft-open
C0272693|ICD9CM|PT|815.14|Open fracture of neck of metacarpal bone(s)
C0272693|ICD9CM|AB|815.14|Fx metacarpal neck-open
C0272729|ICD9CM|PT|821.00|Closed fracture of unspecified part of femur
C0272729|ICD9CM|AB|821.00|Fx femur NOS-closed
C0272751|ICD9CM|PT|820.8|Closed fracture of unspecified part of neck of femur
C0272751|ICD9CM|AB|820.8|Fx neck of femur NOS-cl
C0272752|ICD9CM|PT|820.9|Open fracture of unspecified part of neck of femur
C0272752|ICD9CM|AB|820.9|Fx neck of femur NOS-opn
C0272754|ICD9CM|PT|821.21|Closed fracture of condyle, femoral
C0272754|ICD9CM|AB|821.21|Fx femoral condyle-close
C0272757|ICD9CM|PT|821.31|Open fracture of condyle, femoral
C0272757|ICD9CM|AB|821.31|Fx femoral condyle-open
C0272769|ICD9CM|PT|824.8|Unspecified fracture of ankle, closed
C0272769|ICD9CM|AB|824.8|Fx ankle NOS-closed
C0272770|ICD9CM|PT|824.9|Unspecified fracture of ankle, open
C0272770|ICD9CM|AB|824.9|Fx ankle NOS-open
C0272776|ICD9CM|PT|825.20|Closed fracture of unspecified bone(s) of foot [except toes]
C0272776|ICD9CM|AB|825.20|Fx foot bone NOS-closed
C0272778|ICD9CM|PT|825.30|Open fracture of unspecified bone(s) of foot [except toes]
C0272778|ICD9CM|AB|825.30|Fx foot bone NOS-open
C0272826|ICD9CM|PT|833.15|Open dislocation of metacarpal (bone), proximal end
C0272826|ICD9CM|AB|833.15|Dislocat metacarpal-open
C0272828|ICD9CM|PT|834.01|Closed dislocation of metacarpophalangeal (joint)
C0272828|ICD9CM|AB|834.01|Disloc metacarpophaln-cl
C0272842|ICD9CM|PT|836.60|Dislocation of knee, unspecified, open
C0272842|ICD9CM|AB|836.60|Dislocat knee NOS-open
C0272870|ICD9CM|PT|840.0|Acromioclavicular (joint) (ligament) sprain
C0272870|ICD9CM|AB|840.0|Sprain acromioclavicular
C0272880|ICD9CM|PT|842.01|Sprain of carpal (joint) of wrist
C0272880|ICD9CM|AB|842.01|Sprain carpal
C0272881|ICD9CM|PT|842.02|Sprain of radiocarpal (joint) (ligament) of wrist
C0272881|ICD9CM|AB|842.02|Sprain radiocarpal
C0272905|ICD9CM|PT|845.11|Sprain of tarsometatarsal (joint) (ligament) of foot
C0272905|ICD9CM|AB|845.11|Sprain tarsometatarsal
C0272914|ICD9CM|PT|846.0|Sprain of lumbosacral (joint) (ligament)
C0272914|ICD9CM|AB|846.0|Sprain lumbosacral
C0272920|ICD9CM|AB|848.41|Sprain sternoclavicular
C0272920|ICD9CM|PT|848.41|Sprain of sternoclavicular (joint) (ligament)
C0272955|ICD9CM|PT|851.03|Cortex (cerebral) contusion without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0272955|ICD9CM|AB|851.03|Cortex contus-mod coma
C0272961|ICD9CM|PT|851.11|Cortex (cerebral) contusion with open intracranial wound, with no loss of consciousness
C0272961|ICD9CM|AB|851.11|Opn cortx contus-no coma
C0272966|ICD9CM|PT|851.16|Cortex (cerebral) contusion with open intracranial wound, with loss of consciousness of unspecified duration
C0272966|ICD9CM|AB|851.16|Opn cort contus-coma NOS
C0272967|ICD9CM|PT|851.19|Cortex (cerebral) contusion with open intracranial wound, with concussion, unspecified
C0272967|ICD9CM|AB|851.19|Opn cortx contus-concuss
C0272977|ICD9CM|HT|851.3|Cortex (cerebral) laceration with open intracranial wound
C0272978|ICD9CM|PT|851.30|Cortex (cerebral) laceration with open intracranial wound, unspecified state of consciousness
C0272978|ICD9CM|AB|851.30|Cortex lacer w opn wound
C0272979|ICD9CM|PT|851.31|Cortex (cerebral) laceration with open intracranial wound, with no loss of consciousness
C0272979|ICD9CM|AB|851.31|Opn cortex lacer-no coma
C0272984|ICD9CM|PT|851.36|Cortex (cerebral) laceration with open intracranial wound, with loss of consciousness of unspecified duration
C0272984|ICD9CM|AB|851.36|Opn cortx lacer-coma NOS
C0272985|ICD9CM|PT|851.39|Cortex (cerebral) laceration with open intracranial wound, with concussion, unspecified
C0272985|ICD9CM|AB|851.39|Opn cortx lacer-concuss
C0273088|ICD9CM|PT|852.19|Subarachnoid hemorrhage following injury with open intracranial wound, with concussion, unspecified
C0273088|ICD9CM|AB|852.19|Opn subarach hem-concuss
C0273097|ICD9CM|PT|852.39|Subdural hemorrhage following injury with open intracranial wound, with concussion, unspecified
C0273097|ICD9CM|AB|852.39|Opn subdur hem-concuss
C0273099|ICD9CM|PT|852.40|Extradural hemorrhage following injury without mention of open intracranial wound, unspecified state of consciousness
C0273099|ICD9CM|AB|852.40|Traumatic extradural hem
C0273100|ICD9CM|PT|852.41|Extradural hemorrhage following injury without mention of open intracranial wound, with no loss of consciousness
C0273100|ICD9CM|AB|852.41|Extradural hem w/o coma
C0273104|ICD9CM|PT|852.46|Extradural hemorrhage following injury without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0273104|ICD9CM|PT|852.45|Extradural hemorrhage following injury without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0273104|ICD9CM|AB|852.46|Extradural hem-coma NOS
C0273104|ICD9CM|AB|852.45|Extradural hem-deep coma
C0273106|ICD9CM|PT|852.59|Extradural hemorrhage following injury with open intracranial wound, with concussion, unspecified
C0273106|ICD9CM|AB|852.59|Extradural hem-concuss
C0273127|ICD9CM|PT|862.9|Injury to multiple and unspecified intrathoracic organs, with open wound into cavity
C0273127|ICD9CM|AB|862.9|Intrathorac inj NOS-open
C0273164|ICD9CM|PT|863.81|Injury to pancreas, head, without mention of open wound into cavity
C0273164|ICD9CM|AB|863.81|Pancreas, head inj-close
C0273175|ICD9CM|PT|864.03|Injury to liver without mention of open wound into cavity, laceration, moderate
C0273175|ICD9CM|AB|864.03|Liver laceration, mod
C0273182|ICD9CM|PT|864.14|Injury to liver with open wound into cavity, laceration, major
C0273182|ICD9CM|AB|864.14|Liver lacerat, major-opn
C0273197|ICD9CM|PT|866.03|Injury to kidney without mention of open wound into cavity, complete disruption of kidney parenchyma
C0273197|ICD9CM|AB|866.03|Kidney disruption-closed
C0273236|ICD9CM|PT|879.8|Open wound(s) (multiple) of unspecified site(s), without mention of complication
C0273236|ICD9CM|AB|879.8|Open wound site NOS
C0273237|ICD9CM|PT|879.9|Open wound(s) (multiple) of unspecified site(s), complicated
C0273237|ICD9CM|PT|873.39|Open wound of multiple sites of nose, complicated
C0273237|ICD9CM|AB|879.9|Opn wound site NOS-compl
C0273237|ICD9CM|AB|873.39|Mult open wnd nose-compl
C0273244|ICD9CM|PT|870.3|Penetrating wound of orbit, without mention of foreign body
C0273244|ICD9CM|AB|870.3|Penetr wnd orbit w/o FB
C0273248|ICD9CM|AB|872.01|Open wound of auricle
C0273248|ICD9CM|PT|872.01|Open wound of auricle, ear, without mention of complication
C0273250|ICD9CM|PT|872.9|Open wound of ear, part unspecified, complicated
C0273250|ICD9CM|AB|872.9|Open wound ear NOS-compl
C0273251|ICD9CM|HT|872.1|Open wound of external ear, complicated
C0273253|ICD9CM|PT|872.61|Open wound of ear drum, without mention of complication
C0273253|ICD9CM|AB|872.61|Open wound of ear drum
C0273254|ICD9CM|AB|872.62|Open wound of ossicles
C0273254|ICD9CM|PT|872.62|Open wound of ossicles, without mention of complication
C0273256|ICD9CM|AB|872.64|Open wound of cochlea
C0273256|ICD9CM|PT|872.64|Open wound of cochlea, without mention of complication
C0273259|ICD9CM|PT|873.0|Open wound of scalp, without mention of complication
C0273259|ICD9CM|AB|873.0|Open wound of scalp
C0273260|ICD9CM|HT|873.2|Open wound of nose, without mention of complication
C0273260|ICD9CM|PT|873.20|Open wound of nose, unspecified site, without mention of complication
C0273260|ICD9CM|AB|873.20|Open wound of nose NOS
C0273267|ICD9CM|AB|873.41|Open wound of cheek
C0273267|ICD9CM|PT|873.41|Open wound of cheek, without mention of complication
C0273268|ICD9CM|AB|873.42|Open wound of forehead
C0273268|ICD9CM|PT|873.42|Open wound of forehead, without mention of complication
C0273270|ICD9CM|AB|873.43|Open wound of lip
C0273270|ICD9CM|PT|873.43|Open wound of lip, without mention of complication
C0273271|ICD9CM|AB|873.44|Open wound of jaw
C0273271|ICD9CM|PT|873.44|Open wound of jaw, without mention of complication
C0273276|ICD9CM|AB|873.61|Open wound buccal mucosa
C0273276|ICD9CM|PT|873.61|Open wound of buccal mucosa, without mention of complication
C0273277|ICD9CM|AB|873.62|Open wound of gum
C0273277|ICD9CM|PT|873.62|Open wound of gum (alveolar process), without mention of complication
C0273282|ICD9CM|AB|873.65|Open wound of palate
C0273282|ICD9CM|PT|873.65|Open wound of palate, without mention of complication
C0273284|ICD9CM|PT|873.70|Open wound of mouth, unspecified site, complicated
C0273284|ICD9CM|AB|873.70|Open wnd mouth NOS-compl
C0273286|ICD9CM|PT|873.72|Open wound of gum (alveolar process), complicated
C0273286|ICD9CM|AB|873.72|Open wound gum-compl
C0273292|ICD9CM|PT|874.4|Open wound of pharynx, without mention of complication
C0273292|ICD9CM|AB|874.4|Open wound of pharynx
C0273300|ICD9CM|AB|874.01|Open wound of larynx
C0273300|ICD9CM|PT|874.01|Open wound of larynx, without mention of complication
C0273301|ICD9CM|AB|874.02|Open wound of trachea
C0273301|ICD9CM|PT|874.02|Open wound of trachea, without mention of complication
C0273302|ICD9CM|PT|874.2|Open wound of thyroid gland, without mention of complication
C0273302|ICD9CM|AB|874.2|Open wound thyroid gland
C0273313|ICD9CM|PT|875.0|Open wound of chest (wall), without mention of complication
C0273313|ICD9CM|AB|875.0|Open wound of chest
C0273314|ICD9CM|PT|875.1|Open wound of chest (wall), complicated
C0273314|ICD9CM|AB|875.1|Open wound chest-compl
C0273315|ICD9CM|AB|876.0|Open wound of back
C0273315|ICD9CM|PT|876.0|Open wound of back, without mention of complication
C0273318|ICD9CM|AB|877.0|Open wound of buttock
C0273318|ICD9CM|PT|877.0|Open wound of buttock, without mention of complication
C0273329|ICD9CM|PT|878.4|Open wound of vulva, without mention of complication
C0273329|ICD9CM|AB|878.4|Open wound of vulva
C0273330|ICD9CM|PT|878.6|Open wound of vagina, without mention of complication
C0273330|ICD9CM|AB|878.6|Open wound of vagina
C0273354|ICD9CM|PT|880.00|Open wound of shoulder region, without mention of complication
C0273354|ICD9CM|AB|880.00|Open wound of shoulder
C0273365|ICD9CM|PT|883.0|Open wound of finger(s), without mention of complication
C0273365|ICD9CM|AB|883.0|Open wound of finger
C0273387|ICD9CM|PT|887.3|Traumatic amputation of arm and hand (complete) (partial), unilateral, at or above elbow, complicated
C0273387|ICD9CM|AB|887.3|Amput abv elb, unil-comp
C0273389|ICD9CM|PT|887.1|Traumatic amputation of arm and hand (complete) (partial), unilateral, below elbow, complicated
C0273389|ICD9CM|AB|887.1|Amp below elb, unil-comp
C0273412|ICD9CM|PT|893.1|Open wound of toe(s), complicated
C0273412|ICD9CM|AB|893.1|Open wound toe-compl
C0273413|ICD9CM|PT|893.2|Open wound of toe(s), with tendon involvement
C0273413|ICD9CM|AB|893.2|Open wound toe w tendon
C0273417|ICD9CM|PT|896.1|Traumatic amputation of foot (complete) (partial), unilateral, complicated
C0273417|ICD9CM|AB|896.1|Amput foot, unilat-compl
C0273419|ICD9CM|PT|896.3|Traumatic amputation of foot (complete) (partial), bilateral, complicated
C0273419|ICD9CM|AB|896.3|Amputat foot, bilat-comp
C0273433|ICD9CM|PT|925.2|Crushing injury of neck
C0273433|ICD9CM|AB|925.2|Crush inj neck
C0273444|ICD9CM|AB|927.20|Crushing injury of hand
C0273444|ICD9CM|PT|927.20|Crushing injury of hand(s)
C0273445|ICD9CM|PT|927.3|Crushing injury of finger(s)
C0273445|ICD9CM|AB|927.3|Crushing injury finger
C0273448|ICD9CM|PT|928.3|Crushing injury of toe(s)
C0273448|ICD9CM|AB|928.3|Crushing injury toe
C0273454|ICD9CM|HT|901.4|Injury to pulmonary blood vessels
C0273454|ICD9CM|PT|901.40|Injury to pulmonary vessel(s), unspecified
C0273454|ICD9CM|AB|901.40|Inj pulmonary vessel NOS
C0273463|ICD9CM|PT|902.25|Injury to superior mesenteric artery (trunk)
C0273463|ICD9CM|AB|902.25|Inj super mesenteric art
C0273471|ICD9CM|HT|903.0|Injury to axillary blood vessels
C0273471|ICD9CM|PT|903.00|Injury to axillary vessel(s), unspecified
C0273471|ICD9CM|AB|903.00|Inj axillary vessel NOS
C0273478|ICD9CM|PT|904.8|Injury to unspecified blood vessel of lower extremity
C0273478|ICD9CM|AB|904.8|Injury leg vessel NOS
C0273480|ICD9CM|HT|904.4|Injury to popliteal blood vessels
C0273480|ICD9CM|PT|904.40|Injury to popliteal vessel(s), unspecified
C0273480|ICD9CM|AB|904.40|Inj popliteal vessel NOS
C0273483|ICD9CM|AB|951.9|Injury cranial nerve NOS
C0273483|ICD9CM|PT|951.9|Injury to unspecified cranial nerve
C0273520|ICD9CM|PT|952.2|Lumbar spinal cord injury without evidence of spinal bone injury
C0273520|ICD9CM|AB|952.2|Lumbar spinal cord injur
C0273521|ICD9CM|PT|952.3|Sacral spinal cord injury without evidence of spinal bone injury
C0273521|ICD9CM|AB|952.3|Sacral spinal cord injur
C0273529|ICD9CM|PT|955.9|Injury to unspecified nerve of shoulder girdle and upper limb
C0273529|ICD9CM|HT|955|Injury to peripheral nerve(s) of shoulder girdle and upper limb
C0273529|ICD9CM|AB|955.9|Inj nerve shldr/arm NOS
C0273531|ICD9CM|PT|956.9|Injury to unspecified nerve of pelvic girdle and lower limb
C0273531|ICD9CM|AB|956.9|Inj nerve pelv/leg NOS
C0273532|ICD9CM|PT|956.2|Injury to posterior tibial nerve
C0273532|ICD9CM|AB|956.2|Inj posterior tib nerve
C0273533|ICD9CM|PT|956.5|Injury to other specified nerve(s) of pelvic girdle and lower limb
C0273533|ICD9CM|AB|956.5|Inj nerve pelv/leg NEC
C0273631|ICD9CM|PT|911.4|Insect bite, nonvenomous of trunk, without mention of infection
C0273631|ICD9CM|AB|911.4|Insect bite trunk
C0273632|ICD9CM|PT|911.5|Insect bite, nonvenomous of trunk, infected
C0273632|ICD9CM|AB|911.5|Insect bite trunk-infec
C0273867|ICD9CM|PT|915.0|Abrasion or friction burn of finger(s), without mention of infection
C0273867|ICD9CM|AB|915.0|Abrasion finger
C0273869|ICD9CM|PT|915.4|Insect bite, nonvenomous, of finger(s), without mention of infection
C0273869|ICD9CM|AB|915.4|Insect bite finger
C0273934|ICD9CM|HT|940|Burn confined to eye and adnexa
C0273934|ICD9CM|PT|940.9|Unspecified burn of eye and adnexa
C0273934|ICD9CM|AB|940.9|Burn eye & adnexa NOS
C0273940|ICD9CM|PT|941.00|Burn of unspecified degree of face and head, unspecified site
C0273940|ICD9CM|AB|941.00|Burn NOS head-unspec
C0273941|ICD9CM|PT|941.10|Erythema [first degree] of face and head, unspecified site
C0273941|ICD9CM|AB|941.10|1st deg burn head NOS
C0273948|ICD9CM|PT|941.21|Blisters, epidermal loss [second degree] of ear [any part]
C0273948|ICD9CM|AB|941.21|2nd deg burn ear
C0273970|ICD9CM|AB|941.06|Burn NOS scalp
C0273970|ICD9CM|PT|941.06|Burn of unspecified degree of scalp [any part]
C0273982|ICD9CM|AB|941.08|Burn NOS neck
C0273982|ICD9CM|PT|941.08|Burn of unspecified degree of neck
C0273993|ICD9CM|AB|942.01|Burn NOS breast
C0273993|ICD9CM|PT|942.01|Burn of unspecified degree of breast
C0274005|ICD9CM|AB|942.03|Burn NOS abdominal wall
C0274005|ICD9CM|PT|942.03|Burn of unspecified degree of abdominal wall
C0274011|ICD9CM|AB|942.04|Burn NOS back
C0274011|ICD9CM|PT|942.04|Burn of unspecified degree of back [any part]
C0274035|ICD9CM|PT|943.00|Burn of unspecified degree of upper limb, except wrist and hand, unspecified site
C0274035|ICD9CM|AB|943.00|Burn NOS arm-unspec
C0274041|ICD9CM|AB|943.05|Burn NOS shoulder
C0274041|ICD9CM|PT|943.05|Burn of unspecified degree of shoulder
C0274047|ICD9CM|PT|943.06|Burn of unspecified degree of scapular region
C0274047|ICD9CM|AB|943.06|Burn NOS scapula
C0274053|ICD9CM|AB|943.04|Burn NOS axilla
C0274053|ICD9CM|PT|943.04|Burn of unspecified degree of axilla
C0274056|ICD9CM|PT|943.34|Full-thickness skin loss [third degree, not otherwise specified] of axilla
C0274056|ICD9CM|AB|943.34|3rd deg burn axilla
C0274065|ICD9CM|AB|943.02|Burn NOS elbow
C0274065|ICD9CM|PT|943.02|Burn of unspecified degree of elbow
C0274071|ICD9CM|AB|943.01|Burn NOS forearm
C0274071|ICD9CM|PT|943.01|Burn of unspecified degree of forearm
C0274083|ICD9CM|AB|944.07|Burn NOS wrist
C0274083|ICD9CM|PT|944.07|Burn of unspecified degree of wrist
C0274084|ICD9CM|PT|944.17|Erythema [first degree] of wrist
C0274084|ICD9CM|AB|944.17|1st deg burn wrist
C0274089|ICD9CM|PT|944.00|Burn of unspecified degree of hand, unspecified site
C0274089|ICD9CM|AB|944.00|Burn NOS hand-unspec
C0274090|ICD9CM|PT|944.10|Erythema [first degree] of hand, unspecified site
C0274090|ICD9CM|AB|944.10|1st deg burn hand NOS
C0274134|ICD9CM|HT|944.3|Full-thickness skin loss due to burn [third degree NOS] of wrist(s) and hand(s)
C0274137|ICD9CM|HT|945|Burn of lower limb(s)
C0274143|ICD9CM|AB|945.06|Burn NOS thigh
C0274143|ICD9CM|PT|945.06|Burn of unspecified degree of thigh [any part]
C0274149|ICD9CM|AB|945.05|Burn NOS knee
C0274149|ICD9CM|PT|945.05|Burn of unspecified degree of knee
C0274155|ICD9CM|AB|945.04|Burn NOS lower leg
C0274155|ICD9CM|PT|945.04|Burn of unspecified degree of lower leg
C0274161|ICD9CM|AB|945.03|Burn NOS ankle
C0274161|ICD9CM|PT|945.03|Burn of unspecified degree of ankle
C0274167|ICD9CM|AB|945.02|Burn NOS foot
C0274167|ICD9CM|PT|945.02|Burn of unspecified degree of foot
C0274220|ICD9CM|PT|922.32|Contusion of buttock
C0274220|ICD9CM|AB|922.32|Buttock contusion
C0274221|ICD9CM|PT|922.33|Contusion of interscapular region
C0274221|ICD9CM|AB|922.33|Interscplr reg contusion
C0274236|ICD9CM|PT|924.5|Contusion of unspecified part of lower limb
C0274236|ICD9CM|AB|924.5|Contusion leg NOS
C0274237|ICD9CM|HT|924.2|Contusion of ankle and foot, excluding toe(s)
C0274265|ICD9CM|AB|958.0|Air embolism
C0274265|ICD9CM|PT|958.0|Air embolism
C0274267|ICD9CM|PT|958.2|Secondary and recurrent hemorrhage
C0274267|ICD9CM|AB|958.2|Secondary/recur hemorr
C0274271|ICD9CM|PT|E929.9|Late effects of unspecified accident
C0274271|ICD9CM|AB|E929.9|Late eff accident NOS
C0274276|ICD9CM|AB|906.4|Late effect of crushing
C0274276|ICD9CM|PT|906.4|Late effect of crushing
C0274278|ICD9CM|PT|907.0|Late effect of intracranial injury without mention of skull fracture
C0274278|ICD9CM|AB|907.0|Lt eff intracranial inj
C0274287|ICD9CM|PT|992.9|Unspecified effects of heat and light
C0274287|ICD9CM|HT|992|Effects of heat and light
C0274287|ICD9CM|AB|992.9|Heat effect NOS
C0274288|ICD9CM|PT|992.3|Heat exhaustion, anhydrotic
C0274288|ICD9CM|AB|992.3|Heat exhaust-anhydrotic
C0274323|ICD9CM|HT|996.0|Mechanical complication of cardiac device, implant, and graft
C0274323|ICD9CM|PT|996.00|Mechanical complication of unspecified cardiac device, implant, and graft
C0274323|ICD9CM|AB|996.00|Malfunc card dev/grf NOS
C0274338|ICD9CM|PT|996.2|Mechanical complication of nervous system device, implant, and graft
C0274338|ICD9CM|AB|996.2|Malfun neuro device/graf
C0274344|ICD9CM|PT|996.30|Mechanical complication of unspecified genitourinary device, implant, and graft
C0274344|ICD9CM|HT|996.3|Mechanical complication of genitourinary device, implant, and graft
C0274344|ICD9CM|AB|996.30|Malfunc gu dev/graft NOS
C0274354|ICD9CM|PT|996.51|Mechanical complication due to corneal graft
C0274354|ICD9CM|AB|996.51|Corneal grft malfunction
C0274356|ICD9CM|PT|996.53|Mechanical complication due to ocular lens prosthesis
C0274356|ICD9CM|AB|996.53|Lens prosthesis malfunc
C0274357|ICD9CM|PT|996.54|Mechanical complication due to breast prosthesis
C0274357|ICD9CM|AB|996.54|Breast prosth malfunc
C0274370|ICD9CM|PT|996.87|Complications of transplanted intestine
C0274370|ICD9CM|AB|996.87|Comp intestine transplnt
C0274372|ICD9CM|PT|996.93|Complications of reattached finger(s)
C0274372|ICD9CM|AB|996.93|Compl reattached finger
C0274373|ICD9CM|PT|996.95|Complication of reattached foot and toe(s)
C0274373|ICD9CM|AB|996.95|Compl reattached foot
C0274397|ICD9CM|HT|998.1|Hemorrhage or hematoma complicating a procedure
C0274411|ICD9CM|PT|998.81|Emphysema (subcutaneous) (surgical) resulting from procedure
C0274411|ICD9CM|AB|998.81|Emphysema rsult frm proc
C0274435|ICD9CM|AB|999.80|Transfusion reaction NOS
C0274435|ICD9CM|PT|999.80|Transfusion reaction, unspecified
C0274484|ICD9CM|PT|960.6|Poisoning of antimycobacterial antibiotics
C0274484|ICD9CM|AB|960.6|Pois-antimycobac antibio
C0274507|ICD9CM|PT|960.4|Poisoning by tetracycline group
C0274507|ICD9CM|AB|960.4|Poisoning-tetracycline
C0274511|ICD9CM|PT|960.5|Poisoning of cephalosporin group
C0274511|ICD9CM|AB|960.5|Pois-cephalosporin group
C0274526|ICD9CM|HT|962|Poisoning by hormones and synthetic substitutes
C0274535|ICD9CM|PT|962.2|Poisoning by ovarian hormones and synthetic substitutes
C0274535|ICD9CM|AB|962.2|Poisoning-ovarian hormon
C0274594|ICD9CM|AB|964.3|Poisoning-vitamin k
C0274594|ICD9CM|PT|964.3|Poisoning by vitamin K (phytonadione)
C0274602|ICD9CM|PT|964.7|Poisoning by natural blood and blood products
C0274602|ICD9CM|AB|964.7|Poisoning-blood product
C0274609|ICD9CM|PT|965.9|Poisoning by unspecified analgesic and antipyretic
C0274609|ICD9CM|AB|965.9|Pois-analges/antipyr NOS
C0274638|ICD9CM|PT|967.9|Poisoning by unspecified sedative or hypnotic
C0274638|ICD9CM|HT|967|Poisoning by sedatives and hypnotics
C0274638|ICD9CM|AB|967.9|Pois-sedative/hypnot NOS
C0274659|ICD9CM|PT|970.81|Poisoning by cocaine
C0274659|ICD9CM|AB|970.81|Poisoning by cocaine
C0274669|ICD9CM|PT|969.01|Poisoning by monoamine oxidase inhibitors
C0274669|ICD9CM|AB|969.01|Pois monoamine oxidase
C0274692|ICD9CM|AB|969.72|Poisoning by amphetamine
C0274692|ICD9CM|PT|969.72|Poisoning by amphetamines
C0274693|ICD9CM|PT|969.71|Poisoning by caffeine
C0274693|ICD9CM|AB|969.71|Poisoning by caffeine
C0274702|ICD9CM|PT|971.0|Poisoning by parasympathomimetics (cholinergics)
C0274702|ICD9CM|AB|971.0|Pois-parasympathomimetic
C0274714|ICD9CM|PT|971.2|Poisoning by sympathomimetics [adrenergics]
C0274714|ICD9CM|AB|971.2|Poison-sympathomimetics
C0274717|ICD9CM|PT|971.3|Poisoning by sympatholytics [antiadrenergics]
C0274717|ICD9CM|AB|971.3|Poisoning-sympatholytics
C0274829|ICD9CM|HT|980-989.99|TOXIC EFFECTS OF SUBSTANCES CHIEFLY NONMEDICINAL AS TO SOURCE
C0274829|ICD9CM|PT|989.9|Toxic effect of unspecified substance, chiefly nonmedicinal as to source
C0274829|ICD9CM|AB|989.9|Tox eff nonmed subst NOS
C0274842|ICD9CM|HT|982|Toxic effect of solvents other than petroleum based
C0274869|ICD9CM|HT|985|Toxic effect of other metals
C0274870|ICD9CM|PT|987.9|Toxic effect of unspecified gas, fume, or vapor
C0274870|ICD9CM|AB|987.9|Toxic eff gas/vapor NOS
C0274908|ICD9CM|PT|989.6|Toxic effect of soaps and detergents
C0274908|ICD9CM|AB|989.6|Toxic eff soap/detergent
C0274967|ICD9CM|PT|969.1|Poisoning by phenothiazine-based tranquilizers
C0274967|ICD9CM|AB|969.1|Pois-phenothiazine tranq
C0275016|ICD9CM|PT|989.2|Toxic effect of chlorinated hydrocarbons
C0275016|ICD9CM|AB|989.2|Tox eff chlor hydrocarb
C0275551|ICD9CM|PT|567.23|Spontaneous bacterial peritonitis
C0275551|ICD9CM|AB|567.23|Spontan bact peritonitis
C0275566|ICD9CM|AB|039.1|Pulmonary actinomycosis
C0275566|ICD9CM|PT|039.1|Pulmonary actinomycotic infection
C0275567|ICD9CM|AB|039.0|Cutaneous actinomycosis
C0275567|ICD9CM|PT|039.0|Cutaneous actinomycotic infection
C0275590|ICD9CM|PT|005.2|Food poisoning due to Clostridium perfringens (C. welchii)
C0275590|ICD9CM|AB|005.2|Food pois d/t c. perfrin
C0275594|ICD9CM|AB|023.2|Brucella suis
C0275594|ICD9CM|PT|023.2|Brucella suis
C0275654|ICD9CM|PT|098.17|Gonococcal salpingitis, specified as acute
C0275654|ICD9CM|AB|098.17|Acute gc salpingitis
C0275667|ICD9CM|HT|647.1|Gonorrhea complicating pregnancy, childbirth, or the puerperium
C0275742|ICD9CM|AB|033.1|Bordetella parapertussis
C0275742|ICD9CM|PT|033.1|Whooping cough due to bordetella parapertussis [B. parapertussis]
C0275820|ICD9CM|HT|647.0|Syphilis complicating pregnancy, childbirth, or the puerperium
C0275834|ICD9CM|PT|091.4|Adenopathy due to secondary syphilis
C0275834|ICD9CM|AB|091.4|Syphilitic adenopathy
C0275836|ICD9CM|HT|091.5|Uveitis due to secondary syphilis
C0275836|ICD9CM|AB|091.50|Syphilitic uveitis NOS
C0275836|ICD9CM|PT|091.50|Syphilitic uveitis, unspecified
C0275842|ICD9CM|HT|092|Early syphilis, latent
C0275842|ICD9CM|PT|092.9|Early syphilis, latent, unspecified
C0275842|ICD9CM|AB|092.9|Early syphil latent NOS
C0275844|ICD9CM|PT|093.0|Aneurysm of aorta, specified as syphilitic
C0275844|ICD9CM|AB|093.0|Aortic aneurysm, syphil
C0275859|ICD9CM|PT|090.2|Early congenital syphilis, unspecified
C0275859|ICD9CM|AB|090.2|Early congen syph NOS
C0275874|ICD9CM|PT|090.6|Late congenital syphilis, latent
C0275874|ICD9CM|AB|090.6|Late congen syph latent
C0275891|ICD9CM|HT|011.6|Tuberculous pneumonia [any form]
C0275904|ICD9CM|HT|013.9|Unspecified tuberculosis of central nervous system
C0275904|ICD9CM|AB|013.90|Cns TB NOS-unspec
C0275904|ICD9CM|PT|013.90|Unspecified tuberculosis of central nervous system, unspecified
C0275956|ICD9CM|HT|015.6|Tuberculosis of mastoid
C0275976|ICD9CM|HT|002|Typhoid and paratyphoid fevers
C0275982|ICD9CM|PT|008.43|Intestinal infection due to campylobacter
C0275982|ICD9CM|AB|008.43|Int infec campylobacter
C0275990|ICD9CM|PT|102.0|Initial lesions of yaws
C0275990|ICD9CM|AB|102.0|Initial lesions yaws
C0276001|ICD9CM|AB|102.3|Hyperkeratosis of yaws
C0276001|ICD9CM|PT|102.3|Hyperkeratosis due to yaws
C0276007|ICD9CM|AB|102.4|Gummata and ulcers, yaws
C0276007|ICD9CM|PT|102.4|Gummata and ulcers due to yaws
C0276009|ICD9CM|AB|102.5|Gangosa
C0276009|ICD9CM|PT|102.5|Gangosa
C0276026|ICD9CM|PT|482.2|Pneumonia due to Hemophilus influenzae [H. influenzae]
C0276026|ICD9CM|AB|482.2|H.influenzae pneumonia
C0276029|ICD9CM|PT|038.41|Septicemia due to hemophilus influenzae [H. influenzae]
C0276029|ICD9CM|AB|038.41|H. influenae septicemia
C0276058|ICD9CM|PT|008.2|Intestinal infection due to aerobacter aerogenes
C0276058|ICD9CM|AB|008.2|Aerobacter enteritis
C0276063|ICD9CM|PT|038.49|Other septicemia due to gram-negative organisms
C0276063|ICD9CM|HT|038.4|Septicemia due to other gram-negative organisms
C0276063|ICD9CM|AB|038.49|Gram-neg septicemia NEC
C0276088|ICD9CM|PT|038.42|Septicemia due to escherichia coli [E. coli]
C0276088|ICD9CM|AB|038.42|E coli septicemia
C0276089|ICD9CM|PT|482.82|Pneumonia due to escherichia coli [E. coli]
C0276089|ICD9CM|AB|482.82|Pneumonia e coli
C0276148|ICD9CM|PT|049.9|Unspecified non-arthropod-borne viral diseases of central nervous system
C0276148|ICD9CM|AB|049.9|Viral encephalitis NOS
C0276156|ICD9CM|AB|480.0|Adenoviral pneumonia
C0276156|ICD9CM|PT|480.0|Pneumonia due to adenovirus
C0276162|ICD9CM|PT|008.62|Enteritis due to adenovirus
C0276162|ICD9CM|AB|008.62|Intes infec adenovirus
C0276180|ICD9CM|PT|059.01|Monkeypox
C0276180|ICD9CM|AB|059.01|Monkeypox
C0276191|ICD9CM|PT|059.12|Sealpox
C0276191|ICD9CM|AB|059.12|Sealpox
C0276214|ICD9CM|PT|059.21|Tanapox
C0276214|ICD9CM|AB|059.21|Tanapox
C0276249|ICD9CM|PT|053.8|Herpes zoster with unspecified complication
C0276249|ICD9CM|AB|053.8|H zoster complicated NOS
C0276253|ICD9CM|PT|484.1|Pneumonia in cytomegalic inclusion disease
C0276253|ICD9CM|AB|484.1|Pneum w cytomeg incl dis
C0276306|ICD9CM|PT|647.50|Rubella in the mother, unspecified as to episode of care or not applicable
C0276306|ICD9CM|AB|647.50|Rubella in preg-unspec
C0276308|ICD9CM|AB|056.71|Arthritis due to rubella
C0276308|ICD9CM|PT|056.71|Arthritis due to rubella
C0276333|ICD9CM|PT|480.2|Pneumonia due to parainfluenza virus
C0276333|ICD9CM|AB|480.2|Parinfluenza viral pneum
C0276430|ICD9CM|HT|047|Meningitis due to enterovirus
C0276431|ICD9CM|PT|047.0|Meningitis due to coxsackie virus
C0276431|ICD9CM|AB|047.0|Coxsackie virus mening
C0276682|ICD9CM|PT|771.7|Neonatal Candida infection
C0276682|ICD9CM|AB|771.7|Neonatal candida infect
C0276721|ICD9CM|PT|117.8|Infection by dematiacious fungi [Phaehyphomycosis]
C0276721|ICD9CM|AB|117.8|Dematiacious fungi inf
C0276774|ICD9CM|PT|007.9|Unspecified protozoal intestinal disease
C0276774|ICD9CM|AB|007.9|Protozoal intest dis NOS
C0276804|ICD9CM|AB|130.3|Toxoplasma myocarditis
C0276804|ICD9CM|PT|130.3|Myocarditis due to toxoplasmosis
C0276926|ICD9CM|AB|120.0|Schistosoma haematobium
C0276926|ICD9CM|PT|120.0|Schistosomiasis due to schistosoma haematobium
C0277056|ICD9CM|PT|122.6|Echinococcus multilocularis infection, other
C0277056|ICD9CM|AB|122.6|Echinococc multiloc NEC
C0277120|ICD9CM|PT|126.3|Ancylostomiasis due to ancylostoma ceylanicum
C0277120|ICD9CM|AB|126.3|Ancylostoma ceylanicum
C0277351|ICD9CM|PT|132.3|Mixed pediculosis infestation
C0277351|ICD9CM|AB|132.3|Mixed pedicul & phthirus
C0277538|ICD9CM|HT|799.8|Other ill-defined conditions
C0277538|ICD9CM|PT|799.89|Other ill-defined conditions
C0277538|ICD9CM|AB|799.89|Ill-define condition NEC
C0277590|ICD9CM|PT|798.2|Death occurring in less than 24 hours from onset of symptoms, not otherwise explained
C0277590|ICD9CM|AB|798.2|Death within 24 hr sympt
C0278061|ICD9CM|PT|780.97|Altered mental status
C0278061|ICD9CM|AB|780.97|Altered mental status
C0278314|ICD9CM|AB|55.02|Nephrostomy
C0278314|ICD9CM|PT|55.02|Nephrostomy
C0278321|ICD9CM|HT|65.5|Bilateral oophorectomy
C0278321|ICD9CM|PT|65.51|Other removal of both ovaries at same operative episode
C0278321|ICD9CM|AB|65.51|Oth remove both ovaries
C0278372|ICD9CM|PT|93.01|Functional evaluation
C0278372|ICD9CM|AB|93.01|Functional pt evaluation
C0278729|ICD9CM|AB|233.32|Carcinoma in situ vulva
C0278729|ICD9CM|PT|233.32|Carcinoma in situ, vulva
C0280803|ICD9CM|HT|200.5|Primary central nervous system lymphoma
C0281856|ICD9CM|PT|780.96|Generalized pain
C0281856|ICD9CM|AB|780.96|Generalized pain
C0281890|ICD9CM|AB|748.2|Laryngeal web
C0281890|ICD9CM|PT|748.2|Web of larynx
C0282312|ICD9CM|AB|020.0|Bubonic plague
C0282312|ICD9CM|PT|020.0|Bubonic plague
C0282528|ICD9CM|AB|277.86|Peroxisomal disorders
C0282528|ICD9CM|PT|277.86|Peroxisomal disorders
C0282615|ICD9CM|PT|03.1|Division of intraspinal nerve root
C0282615|ICD9CM|AB|03.1|Intraspin nerve root div
C0300922|ICD9CM|PT|12.52|Goniotomy without goniopuncture
C0300922|ICD9CM|AB|12.52|Goniotomy
C0302112|ICD9CM|PT|284.2|Myelophthisis
C0302112|ICD9CM|AB|284.2|Myelophthisis
C0302358|ICD9CM|AB|004.0|Shigella dysenteriae
C0302358|ICD9CM|PT|004.0|Shigella dysenteriae
C0302359|ICD9CM|AB|004.1|Shigella flexneri
C0302359|ICD9CM|PT|004.1|Shigella flexneri
C0302360|ICD9CM|AB|004.2|Shigella boydii
C0302360|ICD9CM|PT|004.2|Shigella boydii
C0302361|ICD9CM|AB|004.3|Shigella sonnei
C0302361|ICD9CM|PT|004.3|Shigella sonnei
C0302362|ICD9CM|AB|023.0|Brucella melitensis
C0302362|ICD9CM|PT|023.0|Brucella melitensis
C0302363|ICD9CM|AB|023.1|Brucella abortus
C0302363|ICD9CM|PT|023.1|Brucella abortus
C0302367|MTH|PN|NOCODE|Other specified megaloblastic anemias, NEC in ICD9CM
C0302367|ICD9CM|AB|281.3|Megaloblastic anemia NEC
C0302367|ICD9CM|PT|281.3|Other specified megaloblastic anemias not elsewhere classified
C0302369|ICD9CM|PT|291.3|Alcohol-induced psychotic disorder with hallucinations
C0302369|ICD9CM|AB|291.3|Alcoh psy dis w hallucin
C0302370|MTH|PN|NOCODE|Special symptoms or syndromes, NEC in ICD9CM_2014
C0302370|ICD9CM|HT|307|Special symptoms or syndromes, not elsewhere classified
C0302371|MTH|PN|NOCODE|Other and unspecified special symptoms or syndromes, NEC in ICD9CM_2014
C0302371|ICD9CM|PT|307.9|Other and unspecified special symptoms or syndromes, not elsewhere classified
C0302371|ICD9CM|AB|307.9|Special symptom NEC/NOS
C0302373|MTH|PN|NOCODE|Other specified disturbances of conduct, NEC in ICD9CM_2014
C0302373|ICD9CM|HT|312.8|Other specified disturbances of conduct, not elsewhere classified
C0302375|MTH|PN|NOCODE|Certain sequelae of myocardial infarction, NEC in ICD9CM_2014
C0302375|ICD9CM|HT|429.7|Certain sequelae of myocardial infarction, not elsewhere classified
C0302376|MTH|PN|NOCODE|Other sequelae of myocardial infarction, NEC in ICD9CM
C0302376|ICD9CM|PT|429.79|Certain sequelae of myocardial infarction, not elsewhere classified, other
C0302376|ICD9CM|AB|429.79|Other sequelae of MI NEC
C0302377|MTH|PN|NOCODE|Pneumonia due to other virus NEC in ICD9CM
C0302377|ICD9CM|AB|480.8|Viral pneumonia NEC
C0302377|ICD9CM|PT|480.8|Pneumonia due to other virus not elsewhere classified
C0302378|MTH|PN|NOCODE|Chronic airway obstruction, NEC in ICD9CM_2014
C0302378|ICD9CM|PT|496|Chronic airway obstruction, not elsewhere classified
C0302378|ICD9CM|AB|496|Chr airway obstruct NEC
C0302379|MTH|PN|NOCODE|Other pulmonary insufficiency, NEC in ICD9CM
C0302379|ICD9CM|PT|518.82|Other pulmonary insufficiency, not elsewhere classified
C0302379|ICD9CM|AB|518.82|Other pulmonary insuff
C0302382|MTH|PN|NOCODE|Functional digestive disorders, NEC in ICD9CM_2014
C0302382|ICD9CM|HT|564|Functional digestive disorders, not elsewhere classified
C0302384|MTH|PN|NOCODE|Other specified disorders of uterus, NEC in ICD9CM
C0302384|ICD9CM|PT|621.8|Other specified disorders of uterus, not elsewhere classified
C0302384|ICD9CM|AB|621.8|Disorders of uterus NEC
C0302388|MTH|PN|NOCODE|Other indications for care or intervention related to labor and delivery, NEC in ICD9CM
C0302388|ICD9CM|HT|659|Other indications for care or intervention related to labor and delivery, not elsewhere classified
C0302396|MTH|PN|NOCODE|Nonallopathic lesions of abdomen and other sites, NEC in ICD9CM
C0302396|ICD9CM|PT|739.9|Nonallopathic lesions, abdomen and other sites
C0302396|ICD9CM|AB|739.9|Somatic dysfunction NEC
C0302397|ICD9CM|PT|759.6|Other hamartoses, not elsewhere classified
C0302397|ICD9CM|AB|759.6|Hamartoses NEC
C0302401|ICD9CM|HT|959|Injury, other and unspecified
C0302406|MTH|PN|NOCODE|Poisoning by other mineral salts, NEC in ICD9CM_2014
C0302406|ICD9CM|PT|974.6|Poisoning by other mineral salts, not elsewhere classified
C0302406|ICD9CM|AB|974.6|Poison-mineral salts NEC
C0302408|MTH|PN|NOCODE|Toxic effect of other pesticides, NEC in ICD9CM_2014
C0302408|ICD9CM|PT|989.4|Toxic effect of other pesticides, not elsewhere classified
C0302408|ICD9CM|AB|989.4|Toxic eff pesticides NEC
C0302409|MTH|PN|NOCODE|Certain adverse effects NEC in ICD9CM_2014
C0302409|ICD9CM|HT|995|Certain adverse effects not elsewhere classified
C0302411|ICD9CM|PT|996.52|Mechanical complication due to graft of other tissue, not elsewhere classified
C0302411|ICD9CM|AB|996.52|Oth tissue graft malfunc
C0302412|ICD9CM|PT|996.59|Mechanical complication due to other implant and internal device, not elsewhere classified
C0302412|ICD9CM|AB|996.59|Malfunc oth device/graft
C0302414|MTH|PN|NOCODE|Central nervous system complications, NEC in ICD9CM_2014
C0302414|ICD9CM|HT|997.0|Central nervous system complications, not elsewhere classified
C0302415|MTH|PN|NOCODE|Complications affecting other specified body systems, NEC in ICD9CM
C0302415|ICD9CM|HT|997.9|Complications affecting other specified body systems, not elsewhere classified
C0302422|MTH|PN|NOCODE|Other specified complications of procedures, NEC in ICD9CM
C0302422|ICD9CM|HT|998.8|Other specified complications of procedures, not elsewhere classified
C0302424|MTH|PN|NOCODE|Generalized vaccinia as a complication of medical care, NEC in ICD9CM_2014
C0302424|ICD9CM|AB|999.0|Generalized vaccinia
C0302424|ICD9CM|PT|999.0|Generalized vaccinia as a complication of medical care, not elsewhere classified
C0302425|MTH|PN|NOCODE|Air embolism as a complication of medical care, NEC in ICD9CM_2014
C0302425|ICD9CM|PT|999.1|Air embolism as a complication of medical care, not elsewhere classified
C0302425|ICD9CM|AB|999.1|Air embol comp med care
C0302426|MTH|PN|NOCODE|Other vascular complications of medical care, NEC in ICD9CM
C0302426|ICD9CM|PT|999.2|Other vascular complications of medical care, not elsewhere classified
C0302426|ICD9CM|AB|999.2|Vasc comp med care NEC
C0302427|MTH|PN|NOCODE|Other infection due to medical care, NEC in ICD9CM
C0302427|ICD9CM|HT|999.3|Other infection due to medical care, not elsewhere classified
C0302428|MTH|PN|NOCODE|Other serum reaction, NEC in ICD9CM
C0302428|ICD9CM|HT|999.5|Other serum reaction, not elsewhere classified
C0302430|MTH|PN|NOCODE|Other and unspecified complications of medical care, NEC in ICD9CM_2014
C0302430|ICD9CM|PT|999.9|Other and unspecified complications of medical care, not elsewhere classified
C0302430|ICD9CM|AB|999.9|Complic med care NEC/NOS
C0302431|ICD9CM|HT|V62.8|Other psychological or physical stress, not elsewhere classified
C0302431|ICD9CM|PT|V62.89|Other psychological or physical stress, not elsewhere classified
C0302431|ICD9CM|AB|V62.89|Psychological stress NEC
C0302433|ICD9CM|PT|V67.51|Follow-up examination, following completed treatment with high-risk medication, not elsewhere classified
C0302433|ICD9CM|AB|V67.51|High-risk rx NEC exam
C0302434|ICD9CM|PT|V70.2|General psychiatric examination, other and unspecified
C0302434|ICD9CM|AB|V70.2|Gen psychiatric exam NEC
C0302440|ICD9CM|HT|E862|Accidental poisoning by petroleum products, other solvents and their vapors, not elsewhere classified
C0302441|ICD9CM|PT|E862.4|Accidental poisoning by other specified solvents, not elsewhere classified
C0302441|ICD9CM|AB|E862.4|Acc poisn-solvents NEC
C0302442|ICD9CM|PT|E862.9|Accidental poisoning by unspecified solvent, not elsewhere classified
C0302442|ICD9CM|AB|E862.9|Acc poisn-solvent NOS
C0302444|ICD9CM|PT|E864.0|Accidental poisoning by corrosive aromatics not elsewhere classified
C0302444|ICD9CM|AB|E864.0|Acc pois-corrosiv aromat
C0302445|ICD9CM|PT|E864.1|Accidental poisoning by acids not elsewhere classified
C0302445|ICD9CM|AB|E864.1|Acc poison-acids
C0302446|ICD9CM|PT|E864.2|Accidental poisoning by caustic alkalis not elsewhere classified
C0302446|ICD9CM|AB|E864.2|Acc poisn-caustic alkali
C0302447|ICD9CM|PT|E864.3|Accidental poisoning by other specified corrosives and caustics not elsewhere classified
C0302447|ICD9CM|AB|E864.3|Acc poison-caustic NEC
C0302448|ICD9CM|PT|E864.4|Accidental poisoning by unspecified corrosives and caustics not elsewhere classified
C0302448|ICD9CM|AB|E864.4|Acc poison-caustic NOS
C0302450|ICD9CM|PT|64.5|Operations for sex transformation, not elsewhere classified
C0302450|ICD9CM|AB|64.5|Sex transformat op NEC
C0302452|ICD9CM|PT|78.81|Diagnostic procedures on bone, not elsewhere classified, scapula, clavicle, and thorax [ribs and sternum]
C0302452|ICD9CM|AB|78.81|Oth dx proced-chest cage
C0302453|ICD9CM|PT|78.89|Diagnostic procedures on bone, not elsewhere classified, other bones
C0302453|ICD9CM|AB|78.89|Other bone dx proc NEC
C0302454|ICD9CM|PT|88.39|X-ray, other and unspecified
C0302454|ICD9CM|AB|88.39|X-ray NEC and NOS
C0302455|ICD9CM|HT|90.1|Microscopic examination of specimen from endocrine gland, not elsewhere classified
C0302456|ICD9CM|PT|90.11|Microscopic examination of specimen from endocrine gland, not elsewhere classified, bacterial smear
C0302456|ICD9CM|AB|90.11|Bact smear-endocrine
C0302457|ICD9CM|PT|90.12|Microscopic examination of specimen from endocrine gland, not elsewhere classified, culture
C0302457|ICD9CM|AB|90.12|Culture-endocrine
C0302458|ICD9CM|PT|90.13|Microscopic examination of specimen from endocrine gland, not elsewhere classified, culture and sensitivity
C0302458|ICD9CM|AB|90.13|C & s-endocrine
C0302459|ICD9CM|PT|90.14|Microscopic examination of specimen from endocrine gland, not elsewhere classified, parasitology
C0302459|ICD9CM|AB|90.14|Parasitology-endocrine
C0302460|ICD9CM|PT|90.15|Microscopic examination of specimen from endocrine gland, not elsewhere classified, toxicology
C0302460|ICD9CM|AB|90.15|Toxicology-endocrine
C0302461|ICD9CM|PT|90.19|Microscopic examination of specimen from endocrine gland, not elsewhere classified, other microscopic examination
C0302461|ICD9CM|AB|90.19|Micro exam-endocrine NEC
C0302462|ICD9CM|PT|97.84|Removal of sutures from trunk, not elsewhere classified
C0302462|ICD9CM|AB|97.84|Remov trunk suture NEC
C0302465|ICD9CM|PT|441.02|Dissection of aorta, abdominal
C0302465|ICD9CM|AB|441.02|Dsct of abdominal aorta
C0302467|ICD9CM|PT|747.20|Anomaly of aorta, unspecified
C0302467|ICD9CM|AB|747.20|Cong anom of aorta NOS
C0302468|ICD9CM|AB|747.62|Renal vessel anomaly
C0302468|ICD9CM|PT|747.62|Renal vessel anomaly
C0302472|ICD9CM|PT|575.12|Acute and chronic cholecystitis
C0302472|ICD9CM|AB|575.12|Acte & chr cholecystitis
C0302473|ICD9CM|HT|997.6|Amputation stump complication
C0302491|ICD9CM|PT|733.13|Pathologic fracture of vertebrae
C0302491|ICD9CM|AB|733.13|Path fx vertebrae
C0302501|ICD9CM|AB|524.02|Mandibular hyperplasia
C0302501|ICD9CM|PT|524.02|Major anomalies of jaw size, mandibular hyperplasia
C0302505|ICD9CM|PT|788.32|Stress incontinence, male
C0302505|ICD9CM|AB|788.32|Stress incontinence male
C0302540|ICD9CM|PT|789.67|Abdominal tenderness, generalized
C0302540|ICD9CM|AB|789.67|Abdmnal tndr generalized
C0302564|ICD9CM|HT|45.2|Diagnostic procedures on large intestine
C0302565|ICD9CM|PT|85.96|Removal of breast tissue expander
C0302565|ICD9CM|AB|85.96|Remov breast tissu expan
C0311223|ICD9CM|PT|726.0|Adhesive capsulitis of shoulder
C0311223|ICD9CM|AB|726.0|Adhesive capsulit shlder
C0311245|ICD9CM|HT|753.1|Cystic kidney disease
C0311245|ICD9CM|PT|753.10|Cystic kidney disease, unspecified
C0311245|ICD9CM|AB|753.10|Cystic kidney diseas NOS
C0311249|ICD9CM|AB|743.06|Cryptophthalmos
C0311249|ICD9CM|PT|743.06|Cryptophthalmos
C0311251|ICD9CM|AB|743.21|Simple buphthalmos
C0311251|ICD9CM|PT|743.21|Simple buphthalmos
C0311262|ICD9CM|PT|557.1|Chronic vascular insufficiency of intestine
C0311262|ICD9CM|AB|557.1|Chr vasc insuff intest
C0311274|ICD9CM|AB|994.2|Effects of hunger
C0311274|ICD9CM|PT|994.2|Effects of hunger
C0311334|ICD9CM|HT|345.1|Generalized convulsive epilepsy
C0311335|ICD9CM|AB|345.3|Grand mal status
C0311335|ICD9CM|PT|345.3|Grand mal status
C0311341|ICD9CM|PT|366.11|Pseudoexfoliation of lens capsule
C0311341|ICD9CM|AB|366.11|Pseudoexfol lens capsule
C0311355|ICD9CM|HT|258.0|Polyglandular activity in multiple endocrine adenomatosis
C0311375|ICD9CM|PT|985.1|Toxic effect of arsenic and its compounds
C0311375|ICD9CM|AB|985.1|Toxic effect arsenic
C0311376|ICD9CM|PT|027.9|Unspecified zoonotic bacterial disease
C0311376|ICD9CM|HT|020-027.99|ZOONOTIC BACTERIAL DISEASES
C0311376|ICD9CM|AB|027.9|Zoonotic bact dis NOS
C0311389|ICD9CM|AB|597.80|Urethritis NOS
C0311389|ICD9CM|PT|597.80|Urethritis, unspecified
C0311394|ICD9CM|AB|719.7|Difficulty in walking
C0311394|ICD9CM|PT|719.7|Difficulty in walking
C0312413|ICD9CM|AB|788.38|Overflow incontinence
C0312413|ICD9CM|PT|788.38|Overflow incontinence
C0314603|ICD9CM|HT|V83-V84.99|GENETICS
C0332544|ICD9CM|AB|783.1|Abnormal weight gain
C0332544|ICD9CM|PT|783.1|Abnormal weight gain
C0332671|ICD9CM|HT|910-919.99|SUPERFICIAL INJURY
C0332679|ICD9CM|HT|925-929.99|CRUSHING INJURY
C0332679|ICD9CM|AB|929.9|Crushing injury NOS
C0332679|ICD9CM|PT|929.9|Crushing injury of unspecified site
C0332686|ICD9CM|PT|949.1|Erythema [first degree], unspecified site
C0332686|ICD9CM|AB|949.1|1st degree burn NOS
C0332687|ICD9CM|PT|949.2|Blisters, epidermal loss [second degree], unspecified site
C0332687|ICD9CM|AB|949.2|2nd degree burn NOS
C0332691|ICD9CM|PT|E988.2|Injury by scald, undetermined whether accidentally or purposely inflicted
C0332691|ICD9CM|AB|E988.2|Undeterm circ-scald
C0332798|ICD9CM|HT|870-897.99|OPEN WOUNDS
C0332815|ICD9CM|PT|E906.4|Bite of nonvenomous arthropod
C0332815|ICD9CM|AB|E906.4|Nonvenom arthropod bite
C0333297|ICD9CM|PT|707.9|Chronic ulcer of unspecified site
C0333297|ICD9CM|AB|707.9|Chronic skin ulcer NOS
C0336949|ICD9CM|AB|E006.3|Bowling
C0336949|ICD9CM|PT|E006.3|Activities involving bowling
C0336962|ICD9CM|AB|E006.1|Horseback riding
C0336962|ICD9CM|PT|E006.1|Activities involving horseback riding
C0336967|ICD9CM|AB|E004.4|Hang gliding
C0336967|ICD9CM|PT|E004.4|Activities involving hang gliding
C0337203|ICD9CM|HT|E830-E838.9|WATER TRANSPORT ACCIDENTS
C0337212|ICD9CM|PT|E881.0|Accidental fall from ladder
C0337212|ICD9CM|AB|E881.0|Fall from ladder
C0337228|ICD9CM|AB|E884.4|Fall from bed
C0337228|ICD9CM|PT|E884.4|Accidental fall from bed
C0337231|ICD9CM|AB|E884.3|Fall from wheelchair
C0337231|ICD9CM|PT|E884.3|Accidental fall from wheelchair
C0337308|ICD9CM|HT|84.1|Amputation of lower limb
C0337308|ICD9CM|PT|84.10|Lower limb amputation, not otherwise specified
C0337308|ICD9CM|AB|84.10|Lower limb amputat NOS
C0337354|ICD9CM|PT|85.22|Resection of quadrant of breast
C0337354|ICD9CM|AB|85.22|Quadrant resect breast
C0337358|ICD9CM|HT|27.6|Palatoplasty
C0337361|ICD9CM|AB|25.4|Radical glossectomy
C0337361|ICD9CM|PT|25.4|Radical glossectomy
C0337363|ICD9CM|AB|42.25|Open biopsy of esophagus
C0337363|ICD9CM|PT|42.25|Open biopsy of esophagus
C0337380|ICD9CM|PT|52.13|Endoscopic retrograde pancreatography [ERP]
C0337380|ICD9CM|AB|52.13|Endosc retro pancreatog
C0337383|ICD9CM|PT|40.3|Regional lymph node excision
C0337383|ICD9CM|AB|40.3|Regional lymph node exc
C0337385|ICD9CM|AB|41.5|Total splenectomy
C0337385|ICD9CM|PT|41.5|Total splenectomy
C0337419|ICD9CM|PT|19.6|Revision of tympanoplasty
C0337419|ICD9CM|AB|19.6|Tympanoplasty revision
C0338381|ICD9CM|HT|320-389.99|DISEASES OF THE NERVOUS SYSTEM AND SENSE ORGANS
C0338388|ICD9CM|PT|047.1|Meningitis due to echo virus
C0338388|ICD9CM|AB|047.1|Echo virus meningitis
C0338439|ICD9CM|HT|013.5|Tuberculous abscess of spinal cord
C0338439|ICD9CM|HT|013.4|Tuberculoma of spinal cord
C0338439|ICD9CM|AB|013.50|TB sp crd abscess-unspec
C0338439|ICD9CM|AB|013.40|Tubrclma sp cord-unspec
C0338439|ICD9CM|PT|013.40|Tuberculoma of spinal cord, unspecified
C0338439|ICD9CM|PT|013.50|Tuberculous abscess of spinal cord, unspecified
C0338451|ICD9CM|HT|331.1|Frontotemporal dementia
C0338480|ICD9CM|HT|346.1|Migraine without aura
C0338502|ICD9CM|PT|377.43|Optic nerve hypoplasia
C0338502|ICD9CM|AB|377.43|Optic nerve hypoplasia
C0338585|ICD9CM|PT|443.21|Dissection of carotid artery
C0338585|ICD9CM|AB|443.21|Dissect carotid artery
C0338586|ICD9CM|PT|443.24|Dissection of vertebral artery
C0338586|ICD9CM|AB|443.24|Dissect vertebral artery
C0338591|ICD9CM|AB|437.7|Transient global amnesia
C0338591|ICD9CM|PT|437.7|Transient global amnesia
C0338608|ICD9CM|HT|300-316.99|NEUROTIC DISORDERS, PERSONALITY DISORDERS, AND OTHER NONPSYCHOTIC MENTAL DISORDERS
C0338629|ICD9CM|PT|290.13|Presenile dementia with depressive features
C0338629|ICD9CM|AB|290.13|Presenile depression
C0338631|ICD9CM|PT|290.21|Senile dementia with depressive features
C0338631|ICD9CM|AB|290.21|Senile depressive
C0338632|ICD9CM|HT|294.1|Dementia in conditions classified elsewhere
C0338738|ICD9CM|PT|304.61|Other specified drug dependence, continuous
C0338738|ICD9CM|AB|304.61|Drug depend NEC-contin
C0338739|ICD9CM|PT|304.62|Other specified drug dependence, episodic
C0338739|ICD9CM|AB|304.62|Drug depend NEC-episodic
C0338749|ICD9CM|PT|304.51|Hallucinogen dependence, continuous
C0338749|ICD9CM|AB|304.51|Hallucinogen dep-contin
C0338750|ICD9CM|PT|304.52|Hallucinogen dependence, episodic
C0338750|ICD9CM|AB|304.52|Hallucinogen dep-episod
C0338757|ICD9CM|PT|304.31|Cannabis dependence, continuous
C0338757|ICD9CM|AB|304.31|Cannabis depend-contin
C0338758|ICD9CM|PT|304.32|Cannabis dependence, episodic
C0338758|ICD9CM|AB|304.32|Cannabis depend-episodic
C0338762|ICD9CM|PT|304.21|Cocaine dependence, continuous
C0338762|ICD9CM|AB|304.21|Cocaine depend-contin
C0338763|ICD9CM|PT|304.22|Cocaine dependence, episodic
C0338763|ICD9CM|AB|304.22|Cocaine depend-episodic
C0338787|ICD9CM|PT|303.01|Acute alcoholic intoxication in alcoholism, continuous
C0338787|ICD9CM|AB|303.01|Ac alcohol intox-contin
C0338788|ICD9CM|PT|303.02|Acute alcoholic intoxication in alcoholism, episodic
C0338788|ICD9CM|AB|303.02|Ac alcohol intox-episod
C0338810|ICD9CM|PT|295.51|Latent schizophrenia, subchronic
C0338810|ICD9CM|AB|295.51|Lat schizophren-subchr
C0338811|ICD9CM|PT|295.52|Latent schizophrenia, chronic
C0338811|ICD9CM|AB|295.52|Latent schizophren-chr
C0338812|ICD9CM|PT|295.53|Latent schizophrenia, subchronic with acute exacerbation
C0338812|ICD9CM|AB|295.53|Lat schizo-subchr/exacer
C0338813|ICD9CM|PT|295.54|Latent schizophrenia, chronic with acute exacerbation
C0338813|ICD9CM|AB|295.54|Latent schizo-chr/exacer
C0338828|ICD9CM|AB|295.75|Schizoaffectve dis-remis
C0338828|ICD9CM|PT|295.75|Schizoaffective disorder, in remission
C0338832|ICD9CM|HT|296.1|Manic disorder, recurrent episode
C0338838|ICD9CM|PT|296.15|Manic affective disorder, recurrent episode, in partial or unspecified remission
C0338838|ICD9CM|AB|296.15|Recur manic-part remiss
C0338839|ICD9CM|PT|296.16|Manic affective disorder, recurrent episode, in full remission
C0338839|ICD9CM|AB|296.16|Recur manic-full remiss
C0338843|ICD9CM|PT|296.05|Bipolar I disorder, single manic episode, in partial or unspecified remission
C0338843|ICD9CM|AB|296.05|Bipol I sing man rem NOS
C0338886|ICD9CM|PT|296.25|Major depressive affective disorder, single episode, in partial or unspecified remission
C0338886|ICD9CM|AB|296.25|Depr psychos-part remiss
C0338893|ICD9CM|PT|296.35|Major depressive affective disorder, recurrent episode, in partial or unspecified remission
C0338893|ICD9CM|AB|296.35|Recur depr psyc-part rem
C0338930|ICD9CM|PT|298.1|Excitative type psychosis
C0338930|ICD9CM|AB|298.1|Excitativ type psychosis
C0338945|ICD9CM|PT|306.1|Respiratory malfunction arising from mental factors
C0338945|ICD9CM|AB|306.1|Psychogenic respir dis
C0338969|ICD9CM|AB|301.21|Introverted personality
C0338969|ICD9CM|PT|301.21|Introverted personality
C0338982|ICD9CM|PT|315.2|Other specific developmental learning difficulties
C0338982|ICD9CM|AB|315.2|Oth learning difficulty
C0338984|ICD9CM|PT|299.01|Autistic disorder, residual state
C0338984|ICD9CM|AB|299.01|Autistic disord-residual
C0339002|ICD9CM|PT|314.00|Attention deficit disorder without mention of hyperactivity
C0339002|ICD9CM|AB|314.00|Attn defic nonhyperact
C0339005|ICD9CM|PT|312.81|Conduct disorder, childhood onset type
C0339005|ICD9CM|AB|312.81|Cndct dsrdr chldhd onst
C0339022|ICD9CM|AB|11.71|Keratomileusis
C0339022|ICD9CM|PT|11.71|Keratomileusis
C0339034|ICD9CM|PT|360.24|Other metallosis of globe
C0339034|ICD9CM|AB|360.24|Other metallosis, eye
C0339058|ICD9CM|HT|374.0|Entropion and trichiasis of eyelid
C0339097|ICD9CM|PT|374.86|Retained foreign body of eyelid
C0339097|ICD9CM|AB|374.86|Old foreign body, eyelid
C0339121|ICD9CM|PT|375.14|Secondary lacrimal atrophy
C0339121|ICD9CM|AB|375.14|Secondary lacrim atrophy
C0339129|ICD9CM|HT|375.3|Acute and unspecified inflammation of lacrimal passages
C0339130|ICD9CM|PT|375.31|Acute canaliculitis, lacrimal
C0339130|ICD9CM|AB|375.31|Acute canaliculitis
C0339150|ICD9CM|PT|802.6|Closed fracture of orbital floor (blow-out)
C0339150|ICD9CM|AB|802.6|Fx orbital floor-closed
C0339151|ICD9CM|PT|802.7|Open fracture of orbital floor (blow-out)
C0339151|ICD9CM|AB|802.7|Fx orbital floor-open
C0339166|ICD9CM|PT|098.40|Gonococcal conjunctivitis (neonatorum)
C0339166|ICD9CM|AB|098.40|Gonococcal conjunctivit
C0339212|ICD9CM|PT|371.70|Corneal deformity, unspecified
C0339212|ICD9CM|AB|371.70|Corneal deformity NOS
C0339249|ICD9CM|HT|371.1|Corneal pigmentations and deposits
C0339277|ICD9CM|PT|371.51|Juvenile epithelial corneal dystrophy
C0339277|ICD9CM|AB|371.51|Juv epith cornea dystrph
C0339286|ICD9CM|PT|371.62|Keratoconus, acute hydrops
C0339286|ICD9CM|AB|371.62|Keratoconus, ac hydrops
C0339295|ICD9CM|PT|370.34|Exposure keratoconjunctivitis
C0339295|ICD9CM|AB|370.34|Expsure keratoconjunctiv
C0339308|ICD9CM|HT|364.8|Other disorders of iris and ciliary body
C0339319|ICD9CM|PT|364.11|Chronic iridocyclitis in diseases classified elsewhere
C0339319|ICD9CM|AB|364.11|Chr iridocyl in oth dis
C0339320|ICD9CM|PT|364.23|Lens-induced iridocyclitis
C0339320|ICD9CM|AB|364.23|Lens-induced iridocyclit
C0339394|ICD9CM|PT|363.04|Focal choroiditis and chorioretinitis, peripheral
C0339394|ICD9CM|AB|363.04|Periph focal choroiditis
C0339418|ICD9CM|PT|363.32|Other macular scars
C0339418|ICD9CM|AB|363.32|Macular scars NEC
C0339419|ICD9CM|PT|363.33|Other scars of posterior pole
C0339419|ICD9CM|AB|363.33|Posterior pole scar NEC
C0339427|ICD9CM|PT|363.53|Central dystrophy of choroid, partial
C0339427|ICD9CM|AB|363.53|Part cent choroid dystr
C0339436|ICD9CM|HT|362.5|Degeneration of macula and posterior pole of retina
C0339438|ICD9CM|HT|362|Other retinal disorders
C0339438|ICD9CM|HT|362.8|Other retinal disorders
C0339438|ICD9CM|PT|362.89|Other retinal disorders
C0339438|ICD9CM|AB|362.89|Retinal disorders NEC
C0339440|ICD9CM|HT|361.8|Other forms of retinal detachment
C0339440|ICD9CM|PT|361.89|Other forms of retinal detachment
C0339440|ICD9CM|AB|361.89|Retinal detachment NEC
C0339543|ICD9CM|AB|362.56|Macular puckering
C0339543|ICD9CM|PT|362.56|Macular puckering
C0339572|ICD9CM|PT|365.03|Steroid responders borderline glaucoma
C0339572|ICD9CM|AB|365.03|Steroid responders
C0339573|ICD9CM|PT|365.11|Primary open angle glaucoma
C0339573|ICD9CM|AB|365.11|Prim open angle glaucoma
C0339578|ICD9CM|HT|365.3|Corticosteroid-induced glaucoma
C0339579|ICD9CM|PT|365.31|Corticosteroid-induced glaucoma, glaucomatous stage
C0339579|ICD9CM|AB|365.31|Glauc stage-ster induced
C0339580|ICD9CM|PT|365.32|Corticosteroid-induced glaucoma, residual stage
C0339580|ICD9CM|AB|365.32|Glauc resid-ster induced
C0339593|ICD9CM|PT|365.62|Glaucoma associated with ocular inflammations
C0339593|ICD9CM|AB|365.62|Glaucoma w ocular inflam
C0339594|ICD9CM|PT|365.65|Glaucoma associated with ocular trauma
C0339594|ICD9CM|AB|365.65|Glaucoma w ocular trauma
C0339596|ICD9CM|PT|365.82|Glaucoma with increased episcleral venous pressure
C0339596|ICD9CM|AB|365.82|Glauc w inc episcl press
C0339598|ICD9CM|PT|365.61|Glaucoma associated with pupillary block
C0339598|ICD9CM|AB|365.61|Glauc w pupillary block
C0339611|ICD9CM|AB|378.34|Monofixation syndrome
C0339611|ICD9CM|PT|378.34|Monofixation syndrome
C0339666|ICD9CM|HT|379.5|Nystagmus and other irregular eye movements
C0339670|ICD9CM|HT|367|Disorders of refraction and accommodation
C0339670|ICD9CM|PT|367.9|Unspecified disorder of refraction and accommodation
C0339670|ICD9CM|AB|367.9|Refraction disorder NOS
C0339701|ICD9CM|HT|369.1|Moderate or severe vision impairment, better eye; profound vision impairment of lesser eye
C0339711|ICD9CM|PT|369.4|Legal blindness, as defined in U.S.A.
C0339711|ICD9CM|AB|369.4|Legal blindness-usa def
C0339781|ICD9CM|AB|386.41|Round window fistula
C0339781|ICD9CM|PT|386.41|Round window fistula
C0339782|ICD9CM|AB|386.42|Oval window fistula
C0339782|ICD9CM|PT|386.42|Oval window fistula
C0339876|ICD9CM|PT|464.20|Acute laryngotracheitis without mention of obstruction
C0339876|ICD9CM|AB|464.20|Ac laryngotrach no obstr
C0339877|ICD9CM|PT|464.10|Acute tracheitis without mention of obstruction
C0339877|ICD9CM|AB|464.10|Ac tracheitis no obstruc
C0339891|ICD9CM|PT|35.92|Creation of conduit between right ventricle and pulmonary artery
C0339891|ICD9CM|AB|35.92|Conduit rt vent-pul art
C0339901|ICD9CM|HT|460-466.99|ACUTE RESPIRATORY INFECTIONS
C0339904|ICD9CM|PT|517.2|Lung involvement in systemic sclerosis
C0339904|ICD9CM|AB|517.2|Syst sclerosis lung dis
C0339946|ICD9CM|AB|021.2|Pulmonary tularemia
C0339946|ICD9CM|PT|021.2|Pulmonary tularemia
C0339950|ICD9CM|AB|130.4|Toxoplasma pneumonitis
C0339950|ICD9CM|PT|130.4|Pneumonitis due to toxoplasmosis
C0339951|ICD9CM|PT|486|Pneumonia, organism unspecified
C0339951|ICD9CM|AB|486|Pneumonia, organism NOS
C0339959|ICD9CM|PT|483.1|Pneumonia due to chlamydia
C0339959|ICD9CM|AB|483.1|Pneumonia d/t chlamydia
C0339963|ICD9CM|PT|114.4|Chronic pulmonary coccidioidomycosis
C0339963|ICD9CM|AB|114.4|Ch pl coccidioidomycosis
C0340008|ICD9CM|HT|860|Traumatic pneumothorax and hemothorax
C0340270|ICD9CM|HT|451-459.99|DISEASES OF VEINS AND LYMPHATICS, AND OTHER DISEASES OF CIRCULATORY SYSTEM
C0340283|ICD9CM|PT|411.89|Other acute and subacute forms of ischemic heart disease, other
C0340283|ICD9CM|HT|411.8|Other acute and subacute forms of ischemic heart disease
C0340283|ICD9CM|HT|411|Other acute and subacute forms of ischemic heart disease
C0340283|ICD9CM|AB|411.89|Ac ischemic hrt dis NEC
C0340304|ICD9CM|HT|410.3|Acute myocardial infarction, of inferoposterior wall
C0340308|ICD9CM|HT|410.2|Acute myocardial infarction, of inferolateral wall
C0340334|ICD9CM|PT|093.20|Syphilitic endocarditis of valve, unspecified
C0340334|ICD9CM|AB|093.20|Syphil endocarditis NOS
C0340345|ICD9CM|PT|424.91|Endocarditis in diseases classified elsewhere
C0340345|ICD9CM|AB|424.91|Endocarditis in oth dis
C0340348|ICD9CM|PT|421.1|Acute and subacute infective endocarditis in diseases classified elsewhere
C0340348|ICD9CM|AB|421.1|Ac endocardit in oth dis
C0340419|ICD9CM|PT|425.4|Other primary cardiomyopathies
C0340419|ICD9CM|AB|425.4|Prim cardiomyopathy NEC
C0340422|ICD9CM|PT|425.7|Nutritional and metabolic cardiomyopathy
C0340422|ICD9CM|AB|425.7|Metabolic cardiomyopathy
C0340442|ICD9CM|HT|423|Other diseases of pericardium
C0340443|ICD9CM|PT|420.0|Acute pericarditis in diseases classified elsewhere
C0340443|ICD9CM|AB|420.0|Ac pericardit in oth dis
C0340464|ICD9CM|HT|427.6|Premature beats
C0340464|ICD9CM|AB|427.60|Premature beats NOS
C0340464|ICD9CM|PT|427.60|Premature beats, unspecified
C0340529|ICD9CM|PT|996.83|Complications of transplanted heart
C0340529|ICD9CM|AB|996.83|Compl heart transplant
C0340579|ICD9CM|HT|444.2|Embolism and thrombosis of arteries of the extremities
C0340589|ICD9CM|PT|444.22|Arterial embolism and thrombosis of lower extremity
C0340589|ICD9CM|AB|444.22|Lower extremity embolism
C0340629|ICD9CM|AB|441.9|Aortic aneurysm NOS
C0340629|ICD9CM|PT|441.9|Aortic aneurysm of unspecified site without mention of rupture
C0340643|ICD9CM|PT|441.00|Dissection of aorta, unspecified site
C0340643|ICD9CM|AB|441.00|Dsct of aorta unsp site
C0340648|ICD9CM|PT|414.12|Dissection of coronary artery
C0340648|ICD9CM|AB|414.12|Dissection cor artery
C0340649|ICD9CM|PT|443.22|Dissection of iliac artery
C0340649|ICD9CM|AB|443.22|Dissection iliac artery
C0340692|ICD9CM|HT|451.8|Phlebitis and thrombophlebitis of other sites
C0340692|ICD9CM|PT|451.89|Phlebitis and thrombophlebitis of other sites
C0340692|ICD9CM|AB|451.89|Thrombophlebitis NEC
C0340711|ICD9CM|HT|451.1|Phlebitis and thrombophlebitis of deep vessels of lower extremities
C0340712|ICD9CM|PT|451.2|Phlebitis and thrombophlebitis of lower extremities, unspecified
C0340712|ICD9CM|AB|451.2|Thrombophlebitis leg NOS
C0340797|ICD9CM|PT|747.60|Anomaly of the peripheral vascular system, unspecified site
C0340797|ICD9CM|AB|747.60|Unsp prpherl vasc anomal
C0340970|ICD9CM|PT|288.01|Congenital neutropenia
C0340970|ICD9CM|AB|288.01|Congenital neutropenia
C0341004|ICD9CM|AB|521.05|Odontoclasia
C0341004|ICD9CM|PT|521.05|Odontoclasia
C0341029|ICD9CM|AB|524.05|Macrogenia
C0341029|ICD9CM|PT|524.05|Major anomalies of jaw size, macrogenia
C0341030|ICD9CM|AB|524.06|Microgenia
C0341030|ICD9CM|PT|524.06|Major anomalies of jaw size, microgenia
C0341039|ICD9CM|AB|526.1|Fissural cysts of jaw
C0341039|ICD9CM|PT|526.1|Fissural cysts of jaw
C0341072|ICD9CM|AB|52.51|Proximal pancreatectomy
C0341072|ICD9CM|PT|52.51|Proximal pancreatectomy
C0341089|ICD9CM|PT|564.89|Other functional disorders of intestine
C0341089|ICD9CM|AB|564.89|Funct dis intestine NEC
C0341106|ICD9CM|PT|530.13|Eosinophilic esophagitis
C0341106|ICD9CM|AB|530.13|Eosinophilic esophagitis
C0341245|ICD9CM|PT|535.61|Duodenitis, with hemorrhage
C0341245|ICD9CM|AB|535.61|Duodenitis w hmrhg
C0341558|ICD9CM|HT|008.0|Intestinal infection due to escherichia coli [E. coli]
C0341558|ICD9CM|PT|008.00|Intestinal infection due to E. coli, unspecified
C0341558|ICD9CM|AB|008.00|Intest infec e coli NOS
C0341677|ICD9CM|HT|588|Disorders resulting from impaired renal function
C0341677|ICD9CM|PT|588.9|Unspecified disorder resulting from impaired renal function
C0341677|ICD9CM|AB|588.9|Impaired renal funct NOS
C0341692|ICD9CM|PT|580.0|Acute glomerulonephritis with lesion of proliferative glomerulonephritis
C0341692|ICD9CM|AB|580.0|Ac proliferat nephritis
C0341694|ICD9CM|PT|582.4|Chronic glomerulonephritis with lesion of rapidly progressive glomerulonephritis
C0341694|ICD9CM|AB|582.4|Chr rapid progr nephrit
C0341747|ICD9CM|PT|596.55|Detrusor sphincter dyssynergia
C0341747|ICD9CM|AB|596.55|Detrusr sphinc dyssnrgia
C0341803|ICD9CM|AB|68.23|Endometrial ablation
C0341803|ICD9CM|PT|68.23|Endometrial ablation
C0341804|ICD9CM|PT|65.13|Laparoscopic biopsy of ovary
C0341804|ICD9CM|AB|65.13|Lap biopsy of ovary
C0341858|ICD9CM|PT|617.0|Endometriosis of uterus
C0341858|ICD9CM|AB|617.0|Uterine endometriosis
C0341863|ICD9CM|PT|626.2|Excessive or frequent menstruation
C0341863|ICD9CM|AB|626.2|Excessive menstruation
C0341893|ICD9CM|HT|648.0|Diabetes mellitus complicating pregnancy, childbirth, or the puerperium
C0341893|ICD9CM|PT|648.00|Diabetes mellitus of mother, complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C0341893|ICD9CM|AB|648.00|Diabetes in preg-unspec
C0341894|ICD9CM|PT|648.04|Diabetes mellitus of mother, complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication
C0341894|ICD9CM|AB|648.04|Diabetes-postpartum
C0341896|ICD9CM|PT|648.02|Diabetes mellitus of mother, complicating pregnancy, childbirth, or the puerperium, delivered, with mention of postpartum complication
C0341896|ICD9CM|AB|648.02|Diabetes-delivered w p/p
C0341897|ICD9CM|PT|648.01|Diabetes mellitus of mother, complicating pregnancy, childbirth, or the puerperium, delivered, with or without mention of antepartum condition
C0341897|ICD9CM|AB|648.01|Diabetes-delivered
C0341909|ICD9CM|HT|642|Hypertension complicating pregnancy, childbirth, and the puerperium
C0341930|ICD9CM|HT|642.0|Benign essential hypertension complicating pregnancy, childbirth, and the puerperium
C0341934|ICD9CM|HT|642.3|Transient hypertension of pregnancy
C0341950|ICD9CM|HT|642.5|Severe pre-eclampsia
C0341966|ICD9CM|HT|669.2|Maternal hypotension syndrome
C0341973|ICD9CM|HT|659.2|Maternal pyrexia during labor, unspecified
C0342038|ICD9CM|HT|671.5|Other phlebitis and thrombosis in pregnancy and the puerperium
C0342039|ICD9CM|HT|671.4|Deep phlebothrombosis, postpartum
C0342039|ICD9CM|PT|671.44|Deep phlebothrombosis, postpartum, postpartum condition or complication
C0342039|ICD9CM|AB|671.44|Deep vein thromb-postpar
C0342044|ICD9CM|HT|671.3|Deep phlebothrombosis, antepartum
C0342044|ICD9CM|PT|671.33|Deep phlebothrombosis, antepartum, antepartum condition or complication
C0342044|ICD9CM|PT|671.30|Deep phlebothrombosis, antepartum, unspecified as to episode of care or not applicable
C0342044|ICD9CM|AB|671.30|Deep thromb antepar-unsp
C0342044|ICD9CM|AB|671.33|Deep vein thromb-antepar
C0342054|ICD9CM|PT|671.23|Superficial thrombophlebitis complicating pregnancy and the puerperium, antepartum condition or complication
C0342054|ICD9CM|AB|671.23|Thrombophlebit-antepart
C0342068|ICD9CM|HT|671.0|Varicose veins of legs in pregnancy and the puerperium
C0342105|ICD9CM|HT|240-279.99|ENDOCRINE, NUTRITIONAL AND METABOLIC DISEASES, AND IMMUNITY DISORDERS
C0342115|ICD9CM|PT|241.0|Nontoxic uninodular goiter
C0342115|ICD9CM|AB|241.0|Nontox uninodular goiter
C0342122|ICD9CM|HT|242.0|Toxic diffuse goiter
C0342127|ICD9CM|HT|242.3|Toxic nodular goiter, unspecified type
C0342132|ICD9CM|PT|242.40|Thyrotoxicosis from ectopic thyroid nodule without mention of thyrotoxic crisis or storm
C0342132|ICD9CM|AB|242.40|Thyrotox-ect nod no cris
C0342133|ICD9CM|PT|242.41|Thyrotoxicosis from ectopic thyroid nodule with mention of thyrotoxic crisis or storm
C0342133|ICD9CM|AB|242.41|Thyrotox-ect nod w cris
C0342245|ICD9CM|HT|250.5|Diabetes with ophthalmic manifestations
C0342257|ICD9CM|HT|250.9|Diabetes with unspecified complication
C0342565|ICD9CM|PT|254.8|Other specified diseases of thymus gland
C0342565|ICD9CM|AB|254.8|Diseases of thymus NEC
C0342580|ICD9CM|PT|276.0|Hyperosmolality and/or hypernatremia
C0342580|ICD9CM|AB|276.0|Hyperosmolality
C0342635|ICD9CM|PT|275.5|Hungry bone syndrome
C0342635|ICD9CM|AB|275.5|Hungry bone syndrome
C0342712|ICD9CM|PT|270.3|Disturbances of branched-chain amino-acid metabolism
C0342712|ICD9CM|AB|270.3|Bran-chain amin-acid dis
C0342788|ICD9CM|PT|277.81|Primary carnitine deficiency
C0342788|ICD9CM|AB|277.81|Primary carnitine defncy
C0342957|ICD9CM|PT|998.02|Postoperative shock, septic
C0342957|ICD9CM|AB|998.02|Postop shock, septic
C0342971|ICD9CM|AB|53.51|Incisional hernia repair
C0342971|ICD9CM|PT|53.51|Incisional hernia repair
C0342981|ICD9CM|PT|709.3|Degenerative skin disorders
C0342981|ICD9CM|AB|709.3|Degenerative skin disord
C0343065|ICD9CM|AB|708.3|Dermatographic urticaria
C0343065|ICD9CM|PT|708.3|Dermatographic urticaria
C0343139|ICD9CM|HT|730|Osteomyelitis, periostitis, and other infections involving bone
C0343161|ICD9CM|AB|717.6|Loose body in knee
C0343161|ICD9CM|PT|717.6|Loose body in knee
C0343175|ICD9CM|PT|711.00|Pyogenic arthritis, site unspecified
C0343175|ICD9CM|AB|711.00|Pyogen arthritis-unspec
C0343251|ICD9CM|HT|728.1|Muscular calcification and ossification
C0343312|ICD9CM|AB|771.3|Tetanus neonatorum
C0343312|ICD9CM|PT|771.3|Tetanus neonatorum
C0343372|ICD9CM|PT|001.1|Cholera due to vibrio cholerae el tor
C0343372|ICD9CM|AB|001.1|Cholera d/t vib el tor
C0343375|ICD9CM|AB|002.1|Paratyphoid fever a
C0343375|ICD9CM|PT|002.1|Paratyphoid fever A
C0343376|ICD9CM|AB|002.2|Paratyphoid fever b
C0343376|ICD9CM|PT|002.2|Paratyphoid fever B
C0343377|ICD9CM|AB|002.3|Paratyphoid fever c
C0343377|ICD9CM|PT|002.3|Paratyphoid fever C
C0343379|ICD9CM|PT|008.02|Intestinal infection due to enterotoxigenic E. coli
C0343379|ICD9CM|AB|008.02|Int inf e coli entrtoxgn
C0343380|ICD9CM|PT|008.01|Intestinal infection due to enteropathogenic E. coli
C0343380|ICD9CM|AB|008.01|Int inf e coli entrpath
C0343381|ICD9CM|PT|008.04|Intestinal infection due to enterohemorrhagic E. coli
C0343381|ICD9CM|AB|008.04|Int inf e coli entrhmrg
C0343382|ICD9CM|PT|008.03|Intestinal infection due to enteroinvasive E. coli
C0343382|ICD9CM|AB|008.03|Int inf e coli entrnvsv
C0343398|ICD9CM|AB|007.5|Cyclosporiasis
C0343398|ICD9CM|PT|007.5|Cyclosporiasis
C0343413|ICD9CM|PT|137.0|Late effects of respiratory or unspecified tuberculosis
C0343413|ICD9CM|AB|137.0|Late effect tb, resp/NOS
C0343422|ICD9CM|PT|137.2|Late effects of genitourinary tuberculosis
C0343422|ICD9CM|AB|137.2|Late effect gu TB
C0343487|ICD9CM|HT|034|Streptococcal sore throat and scarlet fever
C0343642|ICD9CM|PT|078.10|Viral warts, unspecified
C0343642|ICD9CM|AB|078.10|Viral warts NOS
C0343653|ICD9CM|PT|074.8|Other specified diseases due to Coxsackie virus
C0343653|ICD9CM|AB|074.8|Coxsackie virus NEC
C0343666|ICD9CM|PT|090.0|Early congenital syphilis, symptomatic
C0343666|ICD9CM|AB|090.0|Early cong syph symptom
C0343676|ICD9CM|HT|091.6|Secondary syphilis of viscera and bone
C0343677|ICD9CM|PT|091.3|Secondary syphilis of skin or mucous membranes
C0343677|ICD9CM|AB|091.3|Secondary syph skin
C0343689|ICD9CM|PT|095.8|Other specified forms of late symptomatic syphilis
C0343689|ICD9CM|AB|095.8|Late sympt syphilis NEC
C0343714|ICD9CM|PT|098.51|Gonococcal synovitis and tenosynovitis
C0343714|ICD9CM|AB|098.51|Gonococcal synovitis
C0343816|ICD9CM|PT|130.8|Multisystemic disseminated toxoplasmosis
C0343816|ICD9CM|AB|130.8|Multisystem toxoplasmos
C0343834|ICD9CM|PT|102.6|Bone and joint lesions due to yaws
C0343834|ICD9CM|AB|102.6|Yaws of bone & joint
C0343846|ICD9CM|HT|117|Other mycoses
C0343891|ICD9CM|PT|114.3|Other forms of progressive coccidioidomycosis
C0343891|ICD9CM|AB|114.3|Progress coccidioid NEC
C0344128|ICD9CM|HT|965.6|Poisoning by antirheumatics [antiphlogistics]
C0344133|ICD9CM|PT|969.2|Poisoning by butyrophenone-based tranquilizers
C0344133|ICD9CM|AB|969.2|Pois-butyrophenone tranq
C0344156|ICD9CM|PT|967.1|Poisoning by chloral hydrate group
C0344156|ICD9CM|AB|967.1|Poisoning-chloral hydrat
C0344213|ICD9CM|PT|93.99|Other respiratory procedures
C0344213|ICD9CM|AB|93.99|Other resp procedures
C0344225|ICD9CM|PT|V45.51|Presence of intrauterine contraceptive device
C0344225|ICD9CM|AB|V45.51|Prsc ntrutr cntrcptv dvc
C0344289|ICD9CM|AB|361.12|Bullous retinoschisis
C0344289|ICD9CM|PT|361.12|Bullous retinoschisis
C0344297|ICD9CM|HT|363.4|Choroidal degenerations
C0344297|ICD9CM|PT|363.40|Choroidal degeneration, unspecified
C0344297|ICD9CM|AB|363.40|Choroidal degen NOS
C0344304|ICD9CM|PT|789.07|Abdominal pain, generalized
C0344304|ICD9CM|AB|789.07|Abdmnal pain generalized
C0344365|ICD9CM|PT|788.21|Incomplete bladder emptying
C0344365|ICD9CM|AB|788.21|Incmplet bldder emptying
C0344436|ICD9CM|AB|599.83|Urethral instability
C0344436|ICD9CM|PT|599.83|Urethral instability
C0344528|ICD9CM|PT|743.41|Congenital anomalies of corneal size and shape
C0344528|ICD9CM|AB|743.41|Anom corneal size/shape
C0344538|ICD9CM|PT|743.47|Specified congenital anomalies of sclera
C0344538|ICD9CM|AB|743.47|Anomalies of sclera
C0344553|ICD9CM|PT|743.57|Specified congenital anomalies of optic disc
C0344553|ICD9CM|AB|743.57|Optic disc anomalies
C0344572|ICD9CM|PT|744.41|Branchial cleft sinus or fistula
C0344572|ICD9CM|AB|744.41|Branch cleft sinus/fistu
C0344616|ICD9CM|PT|745.12|Corrected transposition of great vessels
C0344616|ICD9CM|AB|745.12|Correct transpos grt ves
C0344724|ICD9CM|PT|745.5|Ostium secundum type atrial septal defect
C0344724|ICD9CM|AB|745.5|Secundum atrial sept def
C0345010|ICD9CM|PT|747.22|Atresia and stenosis of aorta
C0345010|ICD9CM|AB|747.22|Aortic atresia/stenosis
C0345205|ICD9CM|PT|751.2|Atresia and stenosis of large intestine, rectum, and anal canal
C0345205|ICD9CM|AB|751.2|Atresia large intestine
C0345377|ICD9CM|PT|755.13|Syndactyly of toes without fusion of bone
C0345377|ICD9CM|AB|755.13|Syndactyl toe-no fusion
C0345380|ICD9CM|PT|754.1|Congenital musculoskeletal deformities of sternocleidomastoid muscle
C0345380|ICD9CM|AB|754.1|Congenital torticollis
C0345904|ICD9CM|PT|155.2|Malignant neoplasm of liver, not specified as primary or secondary
C0345904|ICD9CM|AB|155.2|Malignant neo liver NOS
C0345975|ICD9CM|PT|212.6|Benign neoplasm of thymus
C0345975|ICD9CM|AB|212.6|Benign neoplasm thymus
C0346156|ICD9CM|PT|217|Benign neoplasm of breast
C0346156|ICD9CM|AB|217|Benign neoplasm breast
C0346613|ICD9CM|HT|165|Malignant neoplasm of other and ill-defined sites within the respiratory system and intrathoracic organs
C0346627|ICD9CM|PT|159.0|Malignant neoplasm of intestinal tract, part unspecified
C0346627|ICD9CM|AB|159.0|Malig neo intestine NOS
C0346647|ICD9CM|HT|157|Malignant neoplasm of pancreas
C0346647|ICD9CM|PT|157.9|Malignant neoplasm of pancreas, part unspecified
C0346647|ICD9CM|AB|157.9|Malig neo pancreas NOS
C0346773|ICD9CM|PT|172.2|Malignant melanoma of skin of ear and external auditory canal
C0346773|ICD9CM|AB|172.2|Malig melanoma ear
C0346782|ICD9CM|PT|172.4|Malignant melanoma of skin of scalp and neck
C0346782|ICD9CM|AB|172.4|Mal melanoma scalp/neck
C0346866|ICD9CM|PT|183.3|Malignant neoplasm of broad ligament of uterus
C0346866|ICD9CM|AB|183.3|Mal neo broad ligament
C0346867|ICD9CM|PT|183.5|Malignant neoplasm of round ligament of uterus
C0346867|ICD9CM|AB|183.5|Mal neo round ligament
C0346906|ICD9CM|PT|191.5|Malignant neoplasm of ventricles
C0346906|ICD9CM|AB|191.5|Mal neo cereb ventricle
C0346957|ICD9CM|PT|199.0|Disseminated malignant neoplasm without specification of site
C0346957|ICD9CM|AB|199.0|Malig neo disseminated
C0347055|ICD9CM|PT|196.5|Secondary and unspecified malignant neoplasm of lymph nodes of inguinal region and lower limb
C0347055|ICD9CM|AB|196.5|Mal neo lymph-inguin/leg
C0347071|ICD9CM|HT|190-199.99|MALIGNANT NEOPLASM OF OTHER AND UNSPECIFIED SITES
C0347071|ICD9CM|AB|199.1|Malignant neoplasm NOS
C0347071|ICD9CM|PT|199.1|Other malignant neoplasm without specification of site
C0347129|ICD9CM|PT|569.44|Dysplasia of anus
C0347129|ICD9CM|AB|569.44|Dysplasia of anus
C0347138|ICD9CM|PT|232.1|Carcinoma in situ of eyelid, including canthus
C0347138|ICD9CM|AB|232.1|Ca in situ eyelid
C0347139|ICD9CM|PT|232.2|Carcinoma in situ of skin of ear and external auditory canal
C0347139|ICD9CM|AB|232.2|Ca in situ skin ear
C0347243|ICD9CM|HT|212|Benign neoplasm of respiratory and intrathoracic organs
C0347243|ICD9CM|PT|212.9|Benign neoplasm of respiratory and intrathoracic organs, site unspecified
C0347243|ICD9CM|AB|212.9|Benign neo resp sys NOS
C0347277|ICD9CM|PT|211.5|Benign neoplasm of liver and biliary passages
C0347277|ICD9CM|AB|211.5|Ben neo liver/bile ducts
C0347406|ICD9CM|PT|211.8|Benign neoplasm of retroperitoneum and peritoneum
C0347406|ICD9CM|AB|211.8|Ben neo peritoneum
C0347491|ICD9CM|PT|219.8|Benign neoplasm of other specified parts of uterus
C0347491|ICD9CM|AB|219.8|Benign neo uterus NEC
C0347524|ICD9CM|PT|227.9|Benign neoplasm of endocrine gland, site unspecified
C0347524|ICD9CM|AB|227.9|Benign neo endocrine NOS
C0347525|ICD9CM|PT|227.3|Benign neoplasm of pituitary gland and craniopharyngeal duct
C0347525|ICD9CM|AB|227.3|Benign neo pituitary
C0347564|ICD9CM|AB|879.0|Open wound of breast
C0347564|ICD9CM|PT|879.0|Open wound of breast, without mention of complication
C0347619|ICD9CM|PT|860.1|Traumatic pneumothorax with open wound into thorax
C0347619|ICD9CM|AB|860.1|Traum pneumothorax-open
C0347620|ICD9CM|PT|860.0|Traumatic pneumothorax without mention of open wound into thorax
C0347620|ICD9CM|AB|860.0|Traum pneumothorax-close
C0347621|ICD9CM|PT|860.3|Traumatic hemothorax with open wound into thorax
C0347621|ICD9CM|AB|860.3|Traum hemothorax-open
C0347623|ICD9CM|PT|860.5|Traumatic pneumohemothorax with open wound into thorax
C0347623|ICD9CM|AB|860.5|Traum pneumohemothor-opn
C0347624|ICD9CM|PT|860.4|Traumatic pneumohemothorax without mention of open wound into thorax
C0347624|ICD9CM|AB|860.4|Traum pneumohemothor-cl
C0347815|ICD9CM|PT|825.23|Closed fracture of cuboid
C0347815|ICD9CM|AB|825.23|Fx cuboid-closed
C0347816|ICD9CM|PT|825.33|Open fracture of cuboid
C0347816|ICD9CM|AB|825.33|Fx cuboid-open
C0347854|ICD9CM|PT|008.61|Enteritis due to rotavirus
C0347854|ICD9CM|AB|008.61|Intes infec rotavirus
C0347894|ICD9CM|PT|729.2|Neuralgia, neuritis, and radiculitis, unspecified
C0347894|ICD9CM|AB|729.2|Neuralgia/neuritis NOS
C0347900|ICD9CM|HT|015.5|Tuberculosis of limb bones
C0347900|ICD9CM|PT|015.50|Tuberculosis of limb bones, unspecified
C0347900|ICD9CM|AB|015.50|TB of limb bones-unspec
C0347924|ICD9CM|PT|211.6|Benign neoplasm of pancreas, except islets of Langerhans
C0347924|ICD9CM|AB|211.6|Benign neoplasm pancreas
C0347966|ICD9CM|PT|961.3|Poisoning by quinoline and hydroxyquinoline derivatives
C0347966|ICD9CM|AB|961.3|Pois-quinoline/hydroxyqu
C0348087|ICD9CM|HT|V69|Problems related to lifestyle
C0348089|ICD9CM|PT|V69.2|High-risk sexual behavior
C0348089|ICD9CM|AB|V69.2|High-risk sexual behavr
C0348090|ICD9CM|AB|V69.3|Gambling and betting
C0348090|ICD9CM|PT|V69.3|Gambling and betting
C0348098|ICD9CM|PT|008.69|Enteritis due to other viral enteritis
C0348098|ICD9CM|AB|008.69|Other viral intes infec
C0348133|ICD9CM|PT|038.8|Other specified septicemias
C0348133|ICD9CM|AB|038.8|Septicemia NEC
C0348147|ICD9CM|HT|091.8|Other forms of secondary syphilis
C0348147|ICD9CM|PT|091.89|Other forms of secondary syphilis
C0348147|ICD9CM|AB|091.89|Secondary syphilis NEC
C0348149|ICD9CM|HT|095|Other forms of late syphilis, with symptoms
C0348157|ICD9CM|PT|099.55|Other venereal diseases due to chlamydia trachomatis, unspecified genitourinary site
C0348157|ICD9CM|AB|099.55|Ot VD chlm trch unspf gu
C0348168|ICD9CM|PT|062.8|Other specified mosquito-borne viral encephalitis
C0348168|ICD9CM|AB|062.8|Mosquit-borne enceph NEC
C0348187|ICD9CM|PT|052.8|Chickenpox with unspecified complication
C0348187|ICD9CM|AB|052.8|Varicella complicat NOS
C0348188|ICD9CM|AB|052.9|Varicella uncomplicated
C0348188|ICD9CM|PT|052.9|Varicella without mention of complication
C0348194|ICD9CM|PT|056.9|Rubella without mention of complication
C0348194|ICD9CM|AB|056.9|Rubella uncomplicated
C0348196|ICD9CM|HT|059.0|Other orthopoxvirus infections
C0348196|ICD9CM|PT|059.09|Other orthopoxvirus infections
C0348196|ICD9CM|AB|059.09|Orthopoxvirus infect NEC
C0348276|ICD9CM|PT|122.9|Echinococcosis, other and unspecified
C0348276|ICD9CM|AB|122.9|Echinococcosis NEC/NOS
C0348287|ICD9CM|PT|127.9|Intestinal helminthiasis, unspecified
C0348287|ICD9CM|AB|127.9|Intest helminthiasis NOS
C0348296|ICD9CM|HT|137-139.99|LATE EFFECTS OF INFECTIOUS AND PARASITIC DISEASES
C0348343|ICD9CM|PT|162.9|Malignant neoplasm of bronchus and lung, unspecified
C0348343|ICD9CM|AB|162.9|Mal neo bronch/lung NOS
C0348371|ICD9CM|PT|189.9|Malignant neoplasm of urinary organ, site unspecified
C0348371|ICD9CM|AB|189.9|Mal neo urinary NOS
C0348382|ICD9CM|PT|196.8|Secondary and unspecified malignant neoplasm of lymph nodes of multiple sites
C0348382|ICD9CM|AB|196.8|Mal neo lymph node-mult
C0348393|ICD9CM|HT|200-208.99|MALIGNANT NEOPLASM OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0348402|ICD9CM|HT|231|Carcinoma in situ of respiratory system
C0348402|ICD9CM|PT|231.9|Carcinoma in situ of respiratory system, part unspecified
C0348402|ICD9CM|AB|231.9|Ca in situ resp sys NOS
C0348455|ICD9CM|PT|252.08|Other hyperparathyroidism
C0348455|ICD9CM|AB|252.08|Hyperparathyroidism NEC
C0348461|ICD9CM|PT|255.3|Other corticoadrenal overactivity
C0348461|ICD9CM|AB|255.3|Corticoadren overact NEC
C0348483|ICD9CM|PT|270.2|Other disturbances of aromatic amino-acid metabolism
C0348483|ICD9CM|AB|270.2|Arom amin-acid metab NEC
C0348494|ICD9CM|PT|272.4|Other and unspecified hyperlipidemia
C0348494|ICD9CM|AB|272.4|Hyperlipidemia NEC/NOS
C0348499|ICD9CM|PT|277.39|Other amyloidosis
C0348499|ICD9CM|AB|277.39|Amyloidosis NEC
C0348526|ICD9CM|AB|370.8|Keratitis NEC
C0348526|ICD9CM|PT|370.8|Other forms of keratitis
C0348538|ICD9CM|PT|364.89|Other disorders of iris and ciliary body
C0348538|ICD9CM|AB|364.89|Iris/ciliary disord NEC
C0348579|ICD9CM|PT|394.9|Other and unspecified mitral valve diseases
C0348579|ICD9CM|AB|394.9|Mitral valve dis NEC/NOS
C0348586|ICD9CM|PT|405.99|Other unspecified secondary hypertension
C0348586|ICD9CM|AB|405.99|Second hypertension NEC
C0348588|ICD9CM|PT|413.9|Other and unspecified angina pectoris
C0348588|ICD9CM|AB|413.9|Angina pectoris NEC/NOS
C0348597|ICD9CM|PT|420.99|Other acute pericarditis
C0348597|ICD9CM|AB|420.99|Acute pericarditis NEC
C0348615|ICD9CM|PT|425.18|Other hypertrophic cardiomyopathy
C0348615|ICD9CM|AB|425.18|Oth hyprtrophic cardiomy
C0348621|ICD9CM|HT|426.1|Atrioventricular block, other and unspecified
C0348626|ICD9CM|HT|427.8|Other specified cardiac dysrhythmias
C0348626|ICD9CM|PT|427.89|Other specified cardiac dysrhythmias
C0348626|ICD9CM|AB|427.89|Cardiac dysrhythmias NEC
C0348650|ICD9CM|PT|444.89|Embolism and thrombosis of other specified artery
C0348650|ICD9CM|AB|444.89|Arterial embolism NEC
C0348651|ICD9CM|PT|448.9|Other and unspecified capillary diseases
C0348651|ICD9CM|AB|448.9|Capillary dis NEC/NOS
C0348668|ICD9CM|HT|459|Other disorders of circulatory system
C0348708|ICD9CM|AB|512.89|Other pneumothorax
C0348708|ICD9CM|PT|512.89|Other pneumothorax
C0348712|ICD9CM|HT|518.8|Other diseases of lung
C0348712|ICD9CM|HT|518|Other diseases of lung
C0348717|ICD9CM|HT|520-529.99|DISEASES OF ORAL CAVITY, SALIVARY GLANDS, AND JAWS
C0348719|ICD9CM|PT|521.09|Other dental caries
C0348719|ICD9CM|AB|521.09|Dental caries NEC
C0348727|ICD9CM|HT|530.8|Other specified disorders of esophagus
C0348727|ICD9CM|PT|530.89|Other specified disorders of esophagus
C0348727|ICD9CM|AB|530.89|Other dsrders esophagus
C0348731|ICD9CM|HT|537.8|Other specified disorders of stomach and duodenum
C0348731|ICD9CM|PT|537.89|Other specified disorders of stomach and duodenum
C0348731|ICD9CM|AB|537.89|Gastroduodenal dis NEC
C0348737|ICD9CM|AB|556.8|Other ulcerative colitis
C0348737|ICD9CM|PT|556.8|Other ulcerative colitis
C0348742|ICD9CM|HT|569.4|Other specified disorders of rectum and anus
C0348742|ICD9CM|PT|569.49|Other specified disorders of rectum and anus
C0348742|ICD9CM|AB|569.49|Rectal & anal dis NEC
C0348743|ICD9CM|HT|569.8|Other specified disorders of intestine
C0348743|ICD9CM|PT|569.89|Other specified disorders of intestine
C0348743|ICD9CM|AB|569.89|Intestinal disorders NEC
C0348751|ICD9CM|PT|573.8|Other specified disorders of liver
C0348751|ICD9CM|AB|573.8|Liver disorders NEC
C0348758|ICD9CM|AB|575.8|Dis of gallbladder NEC
C0348758|ICD9CM|PT|575.8|Other specified disorders of gallbladder
C0348759|ICD9CM|PT|576.8|Other specified disorders of biliary tract
C0348759|ICD9CM|AB|576.8|Dis of biliary tract NEC
C0348768|ICD9CM|PT|690.18|Other seborrheic dermatitis
C0348768|ICD9CM|AB|690.18|Sebrrheic dermatitis NEC
C0348769|ICD9CM|PT|599.84|Other specified disorders of urethra
C0348769|ICD9CM|AB|599.84|Oth spcf dsdr urethra
C0348773|ICD9CM|PT|V65.49|Other specified counseling
C0348773|ICD9CM|AB|V65.49|Other specfd counseling
C0348774|ICD9CM|PT|V69.8|Other problems related to lifestyle
C0348774|ICD9CM|AB|V69.8|Oth prblms rltd lfstyle
C0348775|ICD9CM|PT|V69.9|Unspecified problem related to lifestyle
C0348775|ICD9CM|AB|V69.9|Prblm rltd lfstyle NOS
C0348799|ICD9CM|PT|466.11|Acute bronchiolitis due to respiratory syncytial virus (RSV)
C0348799|ICD9CM|AB|466.11|Acu broncholitis d/t RSV
C0348801|ICD9CM|PT|482.32|Pneumonia due to Streptococcus, group B
C0348801|ICD9CM|AB|482.32|Pneumonia strptococcus b
C0348815|ICD9CM|PT|277.02|Cystic fibrosis with pulmonary manifestations
C0348815|ICD9CM|AB|277.02|Cystic fibros w pul man
C0348860|ICD9CM|PT|403.91|Hypertensive chronic kidney disease, unspecified, with chronic kidney disease stage V or end stage renal disease
C0348860|ICD9CM|AB|403.91|Hyp kid NOS w cr kid V
C0348879|ICD9CM|PT|404.92|Hypertensive heart and chronic kidney disease, unspecified, without heart failure and with chronic kidney disease stage V or end stage renal disease
C0348879|ICD9CM|AB|404.92|Hy ht/kd NOS st V w/o hf
C0348903|ICD9CM|PT|099.52|Other venereal diseases due to chlamydia trachomatis, anus and rectum
C0348903|ICD9CM|AB|099.52|Oth VD chlm trch ans rct
C0348904|ICD9CM|PT|099.53|Other venereal diseases due to chlamydia trachomatis, lower genitourinary sites
C0348904|ICD9CM|AB|099.53|Oth VD chlm trch lowr gu
C0349231|ICD9CM|AB|300.20|Phobia NOS
C0349231|ICD9CM|HT|300.2|Phobic disorders
C0349231|ICD9CM|PT|300.20|Phobia, unspecified
C0349249|ICD9CM|PT|300.89|Other somatoform disorders
C0349249|ICD9CM|AB|300.89|Somatoform disorders NEC
C0349403|ICD9CM|HT|V10.7|Personal history of other lymphatic and hematopoietic neoplasms
C0349403|ICD9CM|PT|V10.79|Personal history of other lymphatic and hematopoietic neoplasms
C0349403|ICD9CM|AB|V10.79|Hx-lymphatic malign NEC
C0349458|ICD9CM|AB|622.11|Mild dysplasia of cervix
C0349458|ICD9CM|PT|622.11|Mild dysplasia of cervix
C0349459|ICD9CM|PT|622.12|Moderate dysplasia of cervix
C0349459|ICD9CM|AB|622.12|Mod dysplasia of cervix
C0349579|ICD9CM|PT|621.33|Endometrial hyperplasia with atypia
C0349579|ICD9CM|AB|621.33|Endomet hyperpla w atyp
C0349588|ICD9CM|AB|783.43|Short stature
C0349588|ICD9CM|PT|783.43|Short stature
C0349632|ICD9CM|PT|200.37|Marginal zone lymphoma, spleen
C0349632|ICD9CM|AB|200.37|Margin zone lymph spleen
C0349693|ICD9CM|HT|727.4|Ganglion and cyst of synovium, tendon, and bursa
C0362047|ICD9CM|HT|797-799.99|ILL-DEFINED AND UNKNOWN CAUSES OF MORBIDITY AND MORTALITY
C0362049|ICD9CM|HT|E800-E848.9|TRANSPORT ACCIDENTS
C0362050|ICD9CM|PT|138|Late effects of acute poliomyelitis
C0362050|ICD9CM|AB|138|Late effect acute polio
C0362065|ICD9CM|AB|V25.2|Sterilization
C0362065|ICD9CM|PT|V25.2|Sterilization
C0362068|ICD9CM|AB|V25.3|Menstrual extraction
C0362068|ICD9CM|PT|V25.3|Menstrual extraction
C0362085|ICD9CM|PT|V72.7|Diagnostic skin and sensitization tests
C0362085|ICD9CM|AB|V72.7|Skin/sensitization tests
C0370618|ICD9CM|PT|85.71|Latissimus dorsi myocutaneous flap
C0370618|ICD9CM|AB|85.71|Latiss dorsi myocut flap
C0371436|ICD9CM|PT|34.04|Insertion of intercostal catheter for drainage
C0371436|ICD9CM|AB|34.04|Insert intercostal cath
C0371802|ICD9CM|HT|99.0|Transfusion of blood and blood components
C0372251|ICD9CM|PT|54.92|Removal of foreign body from peritoneal cavity
C0372251|ICD9CM|AB|54.92|Remove FB from periton
C0372415|ICD9CM|PT|60.95|Transurethral balloon dilation of the prostatic urethra
C0372415|ICD9CM|AB|60.95|Trans bal dil pros ureth
C0372525|ICD9CM|PT|47.01|Laparoscopic appendectomy
C0372525|ICD9CM|AB|47.01|Lap appendectomy
C0372565|ICD9CM|PT|70.71|Suture of laceration of vagina
C0372565|ICD9CM|AB|70.71|Suture vagina laceration
C0374921|ICD9CM|PT|005.81|Food poisoning due to Vibrio vulnificus
C0374921|ICD9CM|AB|005.81|Food poisn d/t v. vulnif
C0374931|ICD9CM|PT|008.46|Intestinal infection due to other anaerobes
C0374931|ICD9CM|AB|008.46|Intes infec oth anerobes
C0374932|ICD9CM|PT|008.47|Intestinal infection due to other gram-negative bacteria
C0374932|ICD9CM|AB|008.47|Int inf oth grm neg bctr
C0374933|ICD9CM|PT|008.63|Enteritis due to norwalk virus
C0374933|ICD9CM|AB|008.63|Int inf norwalk virus
C0374934|ICD9CM|PT|008.64|Enteritis due to other small round viruses [SRV's]
C0374934|ICD9CM|AB|008.64|Int inf oth sml rnd vrus
C0374936|ICD9CM|PT|008.66|Enteritis due to astrovirus
C0374936|ICD9CM|AB|008.66|Intes infec astrovirus
C0374937|ICD9CM|PT|008.67|Enteritis due to enterovirus nec
C0374937|ICD9CM|AB|008.67|Int inf enterovirus NEC
C0374939|ICD9CM|PT|010.01|Primary tuberculous infection, bacteriological or histological examination not done
C0374939|ICD9CM|AB|010.01|Prim TB complex-no exam
C0374940|ICD9CM|PT|010.02|Primary tuberculous infection, bacteriological or histological examination unknown (at present)
C0374940|ICD9CM|AB|010.02|Prim TB complex-exm unkn
C0374941|ICD9CM|PT|010.03|Primary tuberculous infection, tubercle bacilli found (in sputum) by microscopy
C0374941|ICD9CM|AB|010.03|Prim TB complex-micro dx
C0374942|ICD9CM|PT|010.04|Primary tuberculous infection, tubercle bacilli not found (in sputum) by microscopy, but found by bacterial culture
C0374942|ICD9CM|AB|010.04|Prim TB complex-cult dx
C0374943|ICD9CM|PT|010.05|Primary tuberculous infection, tubercle bacilli not found by bacteriological examination, but tuberculosis confirmed histologically
C0374943|ICD9CM|AB|010.05|Prim TB complex-histo dx
C0374944|ICD9CM|PT|010.06|Primary tuberculous infection, tubercle bacilli not found by bacteriological or histological examination, but tuberculosis confirmed by other methods [inoculation of animals]
C0374944|ICD9CM|AB|010.06|Prim TB complex-oth test
C0374945|ICD9CM|PT|010.10|Tuberculous pleurisy in primary progressive tuberculosis, unspecified
C0374945|ICD9CM|AB|010.10|Prim TB pleurisy-unspec
C0374946|ICD9CM|PT|010.80|Other primary progressive tuberculosis, unspecified
C0374946|ICD9CM|AB|010.80|Prim prog TB NEC-unspec
C0374952|ICD9CM|PT|011.60|Tuberculous pneumonia [any form], unspecified
C0374952|ICD9CM|AB|011.60|TB pneumonia-unspec
C0374954|ICD9CM|PT|011.80|Other specified pulmonary tuberculosis, unspecified
C0374954|ICD9CM|AB|011.80|Pulmonary TB NEC-unspec
C0374955|ICD9CM|PT|012.30|Tuberculous laryngitis, unspecified
C0374955|ICD9CM|AB|012.30|TB laryngitis-unspec
C0374958|ICD9CM|PT|013.30|Tuberculous abscess of brain, unspecified
C0374958|ICD9CM|AB|013.30|TB brain abscess-unspec
C0374959|ICD9CM|PT|013.80|Other specified tuberculosis of central nervous system, unspecified
C0374959|ICD9CM|AB|013.80|Cns TB NEC-unspec
C0374961|ICD9CM|AB|014.00|TB peritonitis-unspec
C0374961|ICD9CM|PT|014.00|Tuberculous peritonitis, unspecified
C0374962|ICD9CM|PT|014.80|Other tuberculosis of intestines, peritoneum, and mesenteric glands, unspecified
C0374962|ICD9CM|AB|014.80|Intestinal TB NEC-unspec
C0374963|ICD9CM|AB|015.10|TB of hip-unspec
C0374963|ICD9CM|PT|015.10|Tuberculosis of hip, unspecified
C0374964|ICD9CM|AB|015.20|TB of knee-unspec
C0374964|ICD9CM|PT|015.20|Tuberculosis of knee, unspecified
C0374965|ICD9CM|AB|015.60|TB of mastoid-unspec
C0374965|ICD9CM|PT|015.60|Tuberculosis of mastoid, unspecified
C0374966|ICD9CM|PT|015.70|Tuberculosis of other specified bone, unspecified
C0374966|ICD9CM|AB|015.70|TB of bone NEC-unspec
C0374967|ICD9CM|PT|015.80|Tuberculosis of other specified joint, unspecified
C0374967|ICD9CM|AB|015.80|TB of joint NEC-unspec
C0374968|ICD9CM|PT|015.90|Tuberculosis of unspecified bones and joints, unspecified
C0374968|ICD9CM|AB|015.90|TB bone/joint NOS-unspec
C0374969|ICD9CM|AB|016.20|TB of ureter-unspec
C0374969|ICD9CM|PT|016.20|Tuberculosis of ureter, unspecified
C0374970|ICD9CM|PT|016.30|Tuberculosis of other urinary organs, unspecified
C0374970|ICD9CM|AB|016.30|TB urinary NEC-unspec
C0374971|ICD9CM|PT|016.40|Tuberculosis of epididymis, unspecified
C0374971|ICD9CM|AB|016.40|TB epididymis-unspec
C0374972|ICD9CM|PT|016.60|Tuberculous oophoritis and salpingitis, unspecified
C0374972|ICD9CM|AB|016.60|TB ovary & tube-unspec
C0374973|ICD9CM|PT|016.90|Genitourinary tuberculosis, unspecified, unspecified
C0374973|ICD9CM|AB|016.90|Gu TB NOS-unspec
C0374974|ICD9CM|HT|017.0|Tuberculosis of skin and subcutaneous cellular tissue
C0374974|ICD9CM|AB|017.00|TB skin/subcutan-unspec
C0374974|ICD9CM|PT|017.00|Tuberculosis of skin and subcutaneous cellular tissue, unspecified
C0374976|ICD9CM|AB|017.40|TB of ear-unspec
C0374976|ICD9CM|PT|017.40|Tuberculosis of ear, unspecified
C0374977|ICD9CM|AB|017.70|TB of spleen-unspec
C0374977|ICD9CM|PT|017.70|Tuberculosis of spleen, unspecified
C0374978|ICD9CM|AB|017.80|TB esophagus-unspec
C0374978|ICD9CM|PT|017.80|Tuberculosis of esophagus, unspecified
C0374982|ICD9CM|PT|041.00|Streptococcus infection in conditions classified elsewhere and of unspecified site, streptococcus, unspecified
C0374982|ICD9CM|HT|041.0|Streptococcus infection in conditions classified elsewhere and of unspecified site
C0374982|ICD9CM|AB|041.00|Streptococcus unspecf
C0374983|ICD9CM|AB|041.01|Streptococcus group a
C0374983|ICD9CM|PT|041.01|Streptococcus infection in conditions classified elsewhere and of unspecified site, streptococcus, group A
C0374984|ICD9CM|AB|041.02|Streptococcus group b
C0374984|ICD9CM|PT|041.02|Streptococcus infection in conditions classified elsewhere and of unspecified site, streptococcus, group B
C0374985|ICD9CM|AB|041.03|Streptococcus group c
C0374985|ICD9CM|PT|041.03|Streptococcus infection in conditions classified elsewhere and of unspecified site, streptococcus, group C
C0374987|ICD9CM|AB|041.05|Streptococcus group g
C0374987|ICD9CM|PT|041.05|Streptococcus infection in conditions classified elsewhere and of unspecified site, streptococcus, group G
C0374988|ICD9CM|PT|041.09|Streptococcus infection in conditions classified elsewhere and of unspecified site, other streptococcus
C0374988|ICD9CM|AB|041.09|Other streptococcus
C0374989|ICD9CM|HT|041.1|Staphylococcus infection in conditions classified elsewhere and of unspecified site
C0374989|ICD9CM|PT|041.10|Staphylococcus infection in conditions classified elsewhere and of unspecified site, staphylococcus, unspecified
C0374989|ICD9CM|AB|041.10|Staphylococcus unspcfied
C0374990|ICD9CM|PT|041.11|Methicillin susceptible Staphylococcus aureus in conditions classified elsewhere and of unspecified site
C0374990|ICD9CM|AB|041.11|Mth sus Stph aur els/NOS
C0374991|ICD9CM|PT|041.19|Staphylococcus infection in conditions classified elsewhere and of unspecified site, other staphylococcus
C0374991|ICD9CM|AB|041.19|Other staphylococcus
C0374992|ICD9CM|AB|041.81|Mycoplasma
C0374992|ICD9CM|PT|041.81|Other specified bacterial infections in conditions classified elsewhere and of unspecified site, mycoplasma
C0374994|ICD9CM|AB|041.83|Clostridium perfringens
C0374994|ICD9CM|PT|041.83|Other specified bacterial infections in conditions classified elsewhere and of unspecified site, Clostridium perfringens
C0374995|ICD9CM|PT|041.84|Other specified bacterial infections in conditions classified elsewhere and of unspecified site, other anaerobes
C0374995|ICD9CM|AB|041.84|Other anaerobes
C0374996|ICD9CM|PT|041.85|Other specified bacterial infections in conditions classified elsewhere and of unspecified site, other gram-negative organisms
C0374996|ICD9CM|AB|041.85|Oth gram negatv bacteria
C0374997|ICD9CM|AB|041.86|Helicobacter pylori
C0374997|ICD9CM|PT|041.86|Helicobacter pylori [H. pylori]
C0374998|ICD9CM|PT|045.90|Acute poliomyelitis, unspecified, poliovirus, unspecified type
C0374998|ICD9CM|AB|045.90|Ac polio NOS-type NOS
C0375000|ICD9CM|PT|070.20|Viral hepatitis B with hepatic coma, acute or unspecified, without mention of hepatitis delta
C0375000|ICD9CM|AB|070.20|Hpt B acte coma wo dlta
C0375001|ICD9CM|PT|070.21|Viral hepatitis B with hepatic coma, acute or unspecified, with hepatitis delta
C0375001|ICD9CM|AB|070.21|Hpt B acte coma w dlta
C0375002|ICD9CM|PT|070.22|Chronic viral hepatitis B with hepatic coma without hepatitis delta
C0375002|ICD9CM|AB|070.22|Hpt B chrn coma wo dlta
C0375003|ICD9CM|PT|070.23|Chronic viral hepatitis B with hepatic coma with hepatitis delta
C0375003|ICD9CM|AB|070.23|Hpt B chrn coma w dlta
C0375004|ICD9CM|PT|070.30|Viral hepatitis B without mention of hepatic coma, acute or unspecified, without mention of hepatitis delta
C0375004|ICD9CM|AB|070.30|Hpt B acte wo cm wo dlta
C0375005|ICD9CM|PT|070.31|Viral hepatitis B without mention of hepatic coma, acute or unspecified, with hepatitis delta
C0375005|ICD9CM|AB|070.31|Hpt B acte wo cm w dlta
C0375006|ICD9CM|PT|070.32|Chronic viral hepatitis B without mention of hepatic coma without mention of hepatitis delta
C0375006|ICD9CM|AB|070.32|Hpt B chrn wo cm wo dlta
C0375007|ICD9CM|PT|070.33|Chronic viral hepatitis B without mention of hepatic coma with hepatitis delta
C0375007|ICD9CM|AB|070.33|Hpt B chrn wo cm w dlta
C0375009|ICD9CM|PT|070.44|Chronic hepatitis C with hepatic coma
C0375009|ICD9CM|AB|070.44|Chrnc hpt C w hepat Coma
C0375011|ICD9CM|PT|070.52|Hepatitis delta without mention of active hepatitis B disease or hepatic coma
C0375011|ICD9CM|AB|070.52|Hpt dlt wo b wo hpt coma
C0375012|ICD9CM|PT|070.54|Chronic hepatitis C without mention of hepatic coma
C0375012|ICD9CM|AB|070.54|Chrnc hpt C wo hpat coma
C0375013|ICD9CM|PT|078.19|Other specified viral warts
C0375013|ICD9CM|AB|078.19|Oth specfd viral warts
C0375014|ICD9CM|PT|078.88|Other specified diseases due to chlamydiae
C0375014|ICD9CM|AB|078.88|Oth spec dis chlamydiae
C0375016|ICD9CM|AB|079.4|Human papillomavirus
C0375016|ICD9CM|PT|079.4|Human papillomavirus in conditions classified elsewhere and of unspecified site
C0375018|ICD9CM|AB|079.50|Retrovirus, unspecified
C0375018|ICD9CM|PT|079.50|Retrovirus, unspecified
C0375018|ICD9CM|HT|079.5|Retrovirus infection in conditions classified elsewhere and of unspecified site
C0375019|ICD9CM|PT|079.51|Human T-cell lymphotrophic virus, type I [HTLV-I]
C0375019|ICD9CM|AB|079.51|Htlv-1 infection oth dis
C0375020|ICD9CM|PT|079.52|Human T-cell lymphotrophic virus, type II [HTLV-II]
C0375020|ICD9CM|AB|079.52|Htlv-ii infectn oth dis
C0375021|ICD9CM|PT|079.53|Human immunodeficiency virus, type 2 [HIV-2]
C0375021|ICD9CM|AB|079.53|Hiv-2 infection oth dis
C0375022|ICD9CM|PT|079.59|Other specified retrovirus
C0375022|ICD9CM|AB|079.59|Oth specfied retrovirus
C0375023|ICD9CM|PT|079.6|Respiratory syncytial virus (RSV)
C0375023|ICD9CM|AB|079.6|Resprtry syncytial virus
C0375024|ICD9CM|AB|079.81|Hantavirus infection
C0375024|ICD9CM|PT|079.81|Hantavirus infection
C0375025|ICD9CM|PT|079.88|Other specified chlamydial infection
C0375025|ICD9CM|AB|079.88|Oth spcf chlamydial infc
C0375026|ICD9CM|HT|079|Viral and chlamydial infection in conditions classified elsewhere and of unspecified site
C0375026|ICD9CM|HT|079.9|Unspecified viral and chlamydial infection in conditions classified elsewhere and of unspecified site
C0375027|ICD9CM|AB|079.98|Chlamydial infection NOS
C0375027|ICD9CM|PT|079.98|Unspecified chlamydial infection
C0375028|ICD9CM|HT|098.1|Gonococcal infection (acute) of upper genitourinary tract
C0375028|ICD9CM|PT|098.10|Gonococcal infection (acute) of upper genitourinary tract, site unspecified
C0375028|ICD9CM|AB|098.10|Gc (acute) upper gu NOS
C0375029|ICD9CM|PT|098.30|Chronic gonococcal infection of upper genitourinary tract, site unspecified
C0375029|ICD9CM|HT|098.3|Gonococcal infection, chronic, of upper genitourinary tract
C0375029|ICD9CM|AB|098.30|Chr gc upper gu NOS
C0375031|ICD9CM|PT|099.40|Other nongonococcal urethritis, unspecified
C0375031|ICD9CM|AB|099.40|Unspcf nongnccl urethrts
C0375033|ICD9CM|PT|099.49|Other nongonococcal urethritis, other specified organism
C0375033|ICD9CM|AB|099.49|Nongc urth oth spf orgsm
C0375034|ICD9CM|HT|099.5|Other venereal diseases due to Chlamydia trachomatis
C0375035|ICD9CM|PT|099.50|Other venereal diseases due to chlamydia trachomatis, unspecified site
C0375035|ICD9CM|AB|099.50|Oth VD chlm trch unsp st
C0375036|ICD9CM|PT|099.51|Other venereal diseases due to chlamydia trachomatis, pharynx
C0375036|ICD9CM|AB|099.51|Oth VD chlm trch pharynx
C0375039|ICD9CM|PT|099.54|Other venereal diseases due to chlamydia trachomatis, other genitourinary sites
C0375039|ICD9CM|AB|099.54|Oth VD chlm trch oth gu
C0375041|ICD9CM|PT|099.56|Other venereal diseases due to chlamydia trachomatis, peritoneum
C0375041|ICD9CM|AB|099.56|Ot VD chlm trch prtoneum
C0375042|ICD9CM|PT|099.59|Other venereal diseases due to chlamydia trachomatis, other specified site
C0375042|ICD9CM|AB|099.59|Oth VD chlm trch spcf st
C0375046|ICD9CM|PT|114.5|Pulmonary coccidioidomycosis, unspecified
C0375046|ICD9CM|AB|114.5|Pl cocidioidomycosis NOS
C0375065|ICD9CM|PT|171.7|Malignant neoplasm of connective and other soft tissue of trunk, unspecified
C0375065|ICD9CM|AB|171.7|Mal neopl trunk NOS
C0375071|ICD9CM|PT|184.4|Malignant neoplasm of vulva, unspecified site
C0375071|ICD9CM|AB|184.4|Malign neopl vulva NOS
C0375075|ICD9CM|PT|200.00|Reticulosarcoma, unspecified site, extranodal and solid organ sites
C0375075|ICD9CM|AB|200.00|Retclsrc unsp xtrndl org
C0375076|ICD9CM|PT|200.10|Lymphosarcoma, unspecified site, extranodal and solid organ sites
C0375076|ICD9CM|AB|200.10|Lymphsrc unsp xtrndl org
C0375077|ICD9CM|PT|200.20|Burkitt's tumor or lymphoma, unspecified site, extranodal and solid organ sites
C0375077|ICD9CM|AB|200.20|Brkt tmr unsp xtrndl org
C0375078|ICD9CM|PT|200.80|Other named variants of lymphosarcoma and reticulosarcoma, unspecified site, extranodal and solid organ sites
C0375078|ICD9CM|AB|200.80|Oth varn unsp xtrndl org
C0375080|ICD9CM|PT|201.10|Hodgkin's granuloma, unspecified site, extranodal and solid organ sites
C0375080|ICD9CM|AB|201.10|Hdgk grn unsp xtrndl org
C0375081|ICD9CM|PT|201.20|Hodgkin's sarcoma, unspecified site, extranodal and solid organ sites
C0375081|ICD9CM|AB|201.20|Hdgk src unsp xtrndl org
C0375082|ICD9CM|PT|201.40|Hodgkin's disease, lymphocytic-histiocytic predominance, unspecified site, extranodal and solid organ sites
C0375082|ICD9CM|AB|201.40|Lym-hst unsp xtrndl orgn
C0375083|ICD9CM|PT|201.50|Hodgkin's disease, nodular sclerosis, unspecified site, extranodal and solid organ sites
C0375083|ICD9CM|AB|201.50|Ndr sclr unsp xtrndl org
C0375084|ICD9CM|PT|201.60|Hodgkin's disease, mixed cellularity, unspecified site, extranodal and solid organ sites
C0375084|ICD9CM|AB|201.60|Mxd celr unsp xtrndl org
C0375085|ICD9CM|PT|201.70|Hodgkin's disease, lymphocytic depletion, unspecified site, extranodal and solid organ sites
C0375085|ICD9CM|AB|201.70|Lym dplt unsp xtrndl org
C0375086|ICD9CM|PT|201.90|Hodgkin's disease, unspecified type, unspecified site, extranodal and solid organ sites
C0375086|ICD9CM|AB|201.90|Hdgk dis unsp xtrndl org
C0375087|ICD9CM|PT|202.00|Nodular lymphoma, unspecified site, extranodal and solid organ sites
C0375087|ICD9CM|AB|202.00|Ndlr lym unsp xtrndl org
C0375088|ICD9CM|PT|202.10|Mycosis fungoides, unspecified site, extranodal and solid organ sites
C0375088|ICD9CM|AB|202.10|Mycs fng unsp xtrndl org
C0375089|ICD9CM|PT|202.20|Sezary's disease, unspecified site, extranodal and solid organ sites
C0375089|ICD9CM|AB|202.20|Szry dis unsp xtrndl org
C0375090|ICD9CM|PT|202.30|Malignant histiocytosis, unspecified site, extranodal and solid organ sites
C0375090|ICD9CM|AB|202.30|Mlg hist unsp xtrndl org
C0375091|ICD9CM|PT|202.40|Leukemic reticuloendotheliosis, unspecified site, extranodal and solid organ sites
C0375091|ICD9CM|AB|202.40|Lk rtctl unsp xtrndl org
C0375092|ICD9CM|PT|202.50|Letterer-siwe disease, unspecified site, extranodal and solid organ sites
C0375092|ICD9CM|AB|202.50|Ltr-siwe unsp xtrndl org
C0375093|ICD9CM|PT|202.60|Malignant mast cell tumors, unspecified site, extranodal and solid organ sites
C0375093|ICD9CM|AB|202.60|Mlg mast unsp xtrndl org
C0375094|ICD9CM|PT|202.80|Other malignant lymphomas, unspecified site, extranodal and solid organ sites
C0375094|ICD9CM|AB|202.80|Oth lymp unsp xtrndl org
C0375095|ICD9CM|PT|202.90|Other and unspecified malignant neoplasms of lymphoid and histiocytic tissue, unspecified site, extranodal and solid organ sites
C0375095|ICD9CM|AB|202.90|Unsp lym unsp xtrndl org
C0375098|ICD9CM|PT|215.7|Other benign neoplasm of connective and other soft tissue of trunk, unspecified
C0375098|ICD9CM|AB|215.7|Benign neo trunk NOS
C0375110|ICD9CM|PT|238.9|Neoplasm of uncertain behavior, site unspecified
C0375110|ICD9CM|AB|238.9|Uncert behavior neo NOS
C0375111|ICD9CM|PT|239.9|Neoplasm of unspecified nature, site unspecified
C0375111|ICD9CM|AB|239.9|Neoplasm NOS
C0375113|ICD9CM|PT|250.00|Diabetes mellitus without mention of complication, type II or unspecified type, not stated as uncontrolled
C0375113|ICD9CM|AB|250.00|DMII wo cmp nt st uncntr
C0375114|ICD9CM|PT|250.01|Diabetes mellitus without mention of complication, type I [juvenile type], not stated as uncontrolled
C0375114|ICD9CM|AB|250.01|DMI wo cmp nt st uncntrl
C0375115|ICD9CM|PT|250.02|Diabetes mellitus without mention of complication, type II or unspecified type, uncontrolled
C0375115|ICD9CM|AB|250.02|DMII wo cmp uncntrld
C0375116|ICD9CM|PT|250.03|Diabetes mellitus without mention of complication, type I [juvenile type], uncontrolled
C0375116|ICD9CM|AB|250.03|DMI wo cmp uncntrld
C0375117|ICD9CM|PT|250.10|Diabetes with ketoacidosis, type II or unspecified type, not stated as uncontrolled
C0375117|ICD9CM|AB|250.10|DMII keto nt st uncntrld
C0375118|ICD9CM|PT|250.11|Diabetes with ketoacidosis, type I [juvenile type], not stated as uncontrolled
C0375118|ICD9CM|AB|250.11|DMI keto nt st uncntrld
C0375119|ICD9CM|PT|250.12|Diabetes with ketoacidosis, type II or unspecified type, uncontrolled
C0375119|ICD9CM|AB|250.12|DMII ketoacd uncontrold
C0375120|ICD9CM|PT|250.13|Diabetes with ketoacidosis, type I [juvenile type], uncontrolled
C0375120|ICD9CM|AB|250.13|DMI ketoacd uncontrold
C0375121|ICD9CM|HT|250.2|Diabetes mellitus with hyperosmolarity
C0375122|ICD9CM|PT|250.20|Diabetes with hyperosmolarity, type II or unspecified type, not stated as uncontrolled
C0375122|ICD9CM|AB|250.20|DMII hprsm nt st uncntrl
C0375123|ICD9CM|PT|250.21|Diabetes with hyperosmolarity, type I [juvenile type], not stated as uncontrolled
C0375123|ICD9CM|AB|250.21|DMI hprsm nt st uncntrld
C0375124|ICD9CM|PT|250.22|Diabetes with hyperosmolarity, type II or unspecified type, uncontrolled
C0375124|ICD9CM|AB|250.22|DMII hprosmlr uncontrold
C0375125|ICD9CM|PT|250.23|Diabetes with hyperosmolarity, type I [juvenile type], uncontrolled
C0375125|ICD9CM|AB|250.23|DMI hprosmlr uncontrold
C0375126|ICD9CM|PT|250.30|Diabetes with other coma, type II or unspecified type, not stated as uncontrolled
C0375126|ICD9CM|AB|250.30|DMII o cm nt st uncntrld
C0375127|ICD9CM|PT|250.31|Diabetes with other coma, type I [juvenile type], not stated as uncontrolled
C0375127|ICD9CM|AB|250.31|DMI o cm nt st uncntrld
C0375128|ICD9CM|PT|250.32|Diabetes with other coma, type II or unspecified type, uncontrolled
C0375128|ICD9CM|AB|250.32|DMII oth coma uncontrold
C0375129|ICD9CM|PT|250.33|Diabetes with other coma, type I [juvenile type], uncontrolled
C0375129|ICD9CM|AB|250.33|DMI oth coma uncontrold
C0375130|ICD9CM|PT|250.40|Diabetes with renal manifestations, type II or unspecified type, not stated as uncontrolled
C0375130|ICD9CM|AB|250.40|DMII renl nt st uncntrld
C0375131|ICD9CM|PT|250.41|Diabetes with renal manifestations, type I [juvenile type], not stated as uncontrolled
C0375131|ICD9CM|AB|250.41|DMI renl nt st uncntrld
C0375132|ICD9CM|PT|250.42|Diabetes with renal manifestations, type II or unspecified type, uncontrolled
C0375132|ICD9CM|AB|250.42|DMII renal uncntrld
C0375133|ICD9CM|PT|250.43|Diabetes with renal manifestations, type I [juvenile type], uncontrolled
C0375133|ICD9CM|AB|250.43|DMI renal uncntrld
C0375134|ICD9CM|PT|250.50|Diabetes with ophthalmic manifestations, type II or unspecified type, not stated as uncontrolled
C0375134|ICD9CM|AB|250.50|DMII ophth nt st uncntrl
C0375135|ICD9CM|PT|250.51|Diabetes with ophthalmic manifestations, type I [juvenile type], not stated as uncontrolled
C0375135|ICD9CM|AB|250.51|DMI ophth nt st uncntrld
C0375136|ICD9CM|PT|250.53|Diabetes with ophthalmic manifestations, type I [juvenile type], uncontrolled
C0375136|ICD9CM|AB|250.53|DMI ophth uncntrld
C0375137|ICD9CM|PT|250.60|Diabetes with neurological manifestations, type II or unspecified type, not stated as uncontrolled
C0375137|ICD9CM|AB|250.60|DMII neuro nt st uncntrl
C0375138|ICD9CM|PT|250.61|Diabetes with neurological manifestations, type I [juvenile type], not stated as uncontrolled
C0375138|ICD9CM|AB|250.61|DMI neuro nt st uncntrld
C0375139|ICD9CM|PT|250.62|Diabetes with neurological manifestations, type II or unspecified type, uncontrolled
C0375139|ICD9CM|AB|250.62|DMII neuro uncntrld
C0375140|ICD9CM|PT|250.63|Diabetes with neurological manifestations, type I [juvenile type], uncontrolled
C0375140|ICD9CM|AB|250.63|DMI neuro uncntrld
C0375141|ICD9CM|PT|250.70|Diabetes with peripheral circulatory disorders, type II or unspecified type, not stated as uncontrolled
C0375141|ICD9CM|AB|250.70|DMII circ nt st uncntrld
C0375142|ICD9CM|PT|250.71|Diabetes with peripheral circulatory disorders, type I [juvenile type], not stated as uncontrolled
C0375142|ICD9CM|AB|250.71|DMI circ nt st uncntrld
C0375143|ICD9CM|PT|250.72|Diabetes with peripheral circulatory disorders, type II or unspecified type, uncontrolled
C0375143|ICD9CM|AB|250.72|DMII circ uncntrld
C0375144|ICD9CM|PT|250.73|Diabetes with peripheral circulatory disorders, type I [juvenile type], uncontrolled
C0375144|ICD9CM|AB|250.73|DMI circ uncntrld
C0375145|ICD9CM|PT|250.80|Diabetes with other specified manifestations, type II or unspecified type, not stated as uncontrolled
C0375145|ICD9CM|AB|250.80|DMII oth nt st uncntrld
C0375146|ICD9CM|PT|250.81|Diabetes with other specified manifestations, type I [juvenile type], not stated as uncontrolled
C0375146|ICD9CM|AB|250.81|DMI oth nt st uncntrld
C0375147|ICD9CM|PT|250.82|Diabetes with other specified manifestations, type II or unspecified type, uncontrolled
C0375147|ICD9CM|AB|250.82|DMII oth uncntrld
C0375148|ICD9CM|PT|250.83|Diabetes with other specified manifestations, type I [juvenile type], uncontrolled
C0375148|ICD9CM|AB|250.83|DMI oth uncntrld
C0375149|ICD9CM|PT|250.90|Diabetes with unspecified complication, type II or unspecified type, not stated as uncontrolled
C0375149|ICD9CM|AB|250.90|DMII unspf nt st uncntrl
C0375150|ICD9CM|PT|250.91|Diabetes with unspecified complication, type I [juvenile type], not stated as uncontrolled
C0375150|ICD9CM|AB|250.91|DMI unspf nt st uncntrld
C0375151|ICD9CM|PT|250.92|Diabetes with unspecified complication, type II or unspecified type, uncontrolled
C0375151|ICD9CM|AB|250.92|DMII unspf uncntrld
C0375152|ICD9CM|PT|250.93|Diabetes with unspecified complication, type I [juvenile type], uncontrolled
C0375152|ICD9CM|AB|250.93|DMI unspf uncntrld
C0375153|ICD9CM|PT|251.1|Other specified hypoglycemia
C0375153|ICD9CM|AB|251.1|Oth spcf hypoglycemia
C0375155|ICD9CM|PT|283.19|Other non-autoimmune hemolytic anemias
C0375155|ICD9CM|AB|283.19|Oth nonauto hem anemia
C0375157|ICD9CM|PT|295.10|Disorganized type schizophrenia, unspecified
C0375157|ICD9CM|AB|295.10|Hebephrenia-unspec
C0375158|ICD9CM|PT|295.20|Catatonic type schizophrenia, unspecified
C0375158|ICD9CM|AB|295.20|Catatonia-unspec
C0375162|ICD9CM|PT|295.70|Schizoaffective disorder, unspecified
C0375162|ICD9CM|AB|295.70|Schizoaffective dis NOS
C0375164|ICD9CM|PT|296.10|Manic affective disorder, recurrent episode, unspecified
C0375164|ICD9CM|AB|296.10|Recur manic dis-unspec
C0375172|ICD9CM|PT|304.10|Sedative, hypnotic or anxiolytic dependence, unspecified
C0375172|ICD9CM|AB|304.10|Sed,hyp,anxiolyt dep-NOS
C0375174|ICD9CM|PT|304.30|Cannabis dependence, unspecified
C0375174|ICD9CM|AB|304.30|Cannabis depend-unspec
C0375175|ICD9CM|PT|304.40|Amphetamine and other psychostimulant dependence, unspecified
C0375175|ICD9CM|HT|304.4|Amphetamine and other psychostimulant dependence
C0375175|ICD9CM|AB|304.40|Amphetamin depend-unspec
C0375176|ICD9CM|PT|304.70|Combinations of opioid type drug with any other drug dependence, unspecified
C0375176|ICD9CM|AB|304.70|Opioid/other dep-unspec
C0375177|ICD9CM|PT|304.80|Combinations of drug dependence excluding opioid type drug, unspecified
C0375177|ICD9CM|AB|304.80|Comb drug dep NEC-unspec
C0375178|ICD9CM|PT|304.90|Unspecified drug dependence, unspecified
C0375178|ICD9CM|AB|304.90|Drug depend NOS-unspec
C0375179|ICD9CM|PT|305.20|Cannabis abuse, unspecified
C0375179|ICD9CM|AB|305.20|Cannabis abuse-unspec
C0375180|ICD9CM|AB|305.30|Hallucinog abuse-unspec
C0375180|ICD9CM|PT|305.30|Hallucinogen abuse, unspecified
C0375181|ICD9CM|PT|305.40|Sedative, hypnotic or anxiolytic abuse, unspecified
C0375181|ICD9CM|AB|305.40|Sed,hyp,anxiolytc ab-NOS
C0375182|ICD9CM|AB|305.50|Opioid abuse-unspec
C0375182|ICD9CM|PT|305.50|Opioid abuse, unspecified
C0375184|ICD9CM|PT|305.70|Amphetamine or related acting sympathomimetic abuse, unspecified
C0375184|ICD9CM|AB|305.70|Amphetamine abuse-unspec
C0375185|ICD9CM|PT|305.80|Antidepressant type abuse, unspecified
C0375185|ICD9CM|AB|305.80|Antidepress abuse-unspec
C0375189|ICD9CM|PT|312.00|Undersocialized conduct disorder, aggressive type, unspecified
C0375189|ICD9CM|AB|312.00|Unsocial aggress-unspec
C0375190|ICD9CM|PT|312.10|Undersocialized conduct disorder, unaggressive type, unspecified
C0375190|ICD9CM|AB|312.10|Unsocial unaggress-unsp
C0375192|ICD9CM|PT|312.82|Conduct disorder, adolescent onset type
C0375192|ICD9CM|AB|312.82|Cndct dsrdr adlscnt onst
C0375193|ICD9CM|AB|312.89|Other conduct disorder
C0375193|ICD9CM|PT|312.89|Other conduct disorder
C0375197|ICD9CM|AB|320.81|Anaerobic meningitis
C0375197|ICD9CM|PT|320.81|Anaerobic meningitis
C0375198|MTH|PN|NOCODE|Meningitis due to gram-negative bacteria, NEC in ICD9CM_2014
C0375198|ICD9CM|PT|320.82|Meningitis due to gram-negative bacteria, not elsewhere classified
C0375198|ICD9CM|AB|320.82|Mningts gram-neg bct NEC
C0375200|ICD9CM|PT|333.93|Benign shuddering attacks
C0375200|ICD9CM|AB|333.93|Bnign shuddering attacks
C0375204|ICD9CM|PT|337.29|Reflex sympathetic dystrophy of other specified site
C0375204|ICD9CM|AB|337.29|Rflx sym dystrph oth st
C0375206|ICD9CM|HT|342|Hemiplegia and hemiparesis
C0375208|ICD9CM|PT|342.01|Flaccid hemiplegia and hemiparesis affecting dominant side
C0375208|ICD9CM|AB|342.01|Flccd hmiplga domnt side
C0375209|ICD9CM|PT|342.02|Flaccid hemiplegia and hemiparesis affecting nondominant side
C0375209|ICD9CM|AB|342.02|Flccd hmiplg nondmnt sde
C0375211|ICD9CM|PT|342.11|Spastic hemiplegia and hemiparesis affecting dominant side
C0375211|ICD9CM|AB|342.11|Spstc hmiplga domnt side
C0375212|ICD9CM|PT|342.12|Spastic hemiplegia and hemiparesis affecting nondominant side
C0375212|ICD9CM|AB|342.12|Spstc hmiplg nondmnt sde
C0375213|ICD9CM|HT|342.8|Other specified hemiplegia
C0375214|ICD9CM|PT|342.80|Other specified hemiplegia and hemiparesis affecting unspecified side
C0375214|ICD9CM|AB|342.80|Ot sp hmiplga unspf side
C0375215|ICD9CM|PT|342.81|Other specified hemiplegia and hemiparesis affecting dominant side
C0375215|ICD9CM|AB|342.81|Ot sp hmiplga domnt side
C0375216|ICD9CM|PT|342.82|Other specified hemiplegia and hemiparesis affecting nondominant side
C0375216|ICD9CM|AB|342.82|Ot sp hmiplg nondmnt sde
C0375218|ICD9CM|PT|342.90|Hemiplegia, unspecified, affecting unspecified side
C0375218|ICD9CM|AB|342.90|Unsp hemiplga unspf side
C0375219|ICD9CM|PT|342.91|Hemiplegia, unspecified, affecting dominant side
C0375219|ICD9CM|AB|342.91|Unsp hemiplga domnt side
C0375220|ICD9CM|PT|342.92|Hemiplegia, unspecified, affecting nondominant side
C0375220|ICD9CM|AB|342.92|Unsp hmiplga nondmnt sde
C0375221|ICD9CM|HT|344.0|Quadriplegia and quadriparesis
C0375223|ICD9CM|AB|344.09|Other quadriplegia
C0375223|ICD9CM|PT|344.09|Other quadriplegia
C0375224|ICD9CM|PT|344.30|Monoplegia of lower limb affecting unspecified side
C0375224|ICD9CM|AB|344.30|Monplga lwr lmb unsp sde
C0375225|ICD9CM|PT|344.31|Monoplegia of lower limb affecting dominant side
C0375225|ICD9CM|AB|344.31|Monplga lwr lmb dmnt sde
C0375228|ICD9CM|PT|344.41|Monoplegia of upper limb affecting dominant side
C0375228|ICD9CM|AB|344.41|Monplga upr lmb dmnt sde
C0375229|ICD9CM|PT|344.42|Monoplegia of upper limb affecting nondominant sde
C0375229|ICD9CM|AB|344.42|Mnplg upr lmb nondmnt sd
C0375239|ICD9CM|PT|346.90|Migraine, unspecified, without mention of intractable migraine without mention of status migrainosus
C0375239|ICD9CM|AB|346.90|Migrne unsp wo ntrc mgrn
C0375240|ICD9CM|PT|346.91|Migraine, unspecified, with intractable migraine, so stated, without mention of status migrainosus
C0375240|ICD9CM|AB|346.91|Mgrn unsp w ntrc mgr std
C0375242|ICD9CM|PT|355.71|Causalgia of lower limb
C0375242|ICD9CM|AB|355.71|Causalgia lower limb
C0375253|ICD9CM|PT|371.82|Corneal disorder due to contact lens
C0375253|ICD9CM|AB|371.82|Corneal dsdr contct lens
C0375257|ICD9CM|PT|388.40|Abnormal auditory perception, unspecified
C0375257|ICD9CM|AB|388.40|Abn auditory percept NOS
C0375259|ICD9CM|HT|396|Diseases of mitral and aortic valves
C0375259|ICD9CM|PT|396.9|Mitral and aortic valve diseases, unspecified
C0375259|ICD9CM|AB|396.9|Mitral/aortic v dis NOS
C0375264|ICD9CM|PT|414.04|Coronary atherosclerosis of artery bypass graft
C0375264|ICD9CM|AB|414.04|Cor ath artry bypas grft
C0375265|ICD9CM|PT|414.05|Coronary atherosclerosis of unspecified bypass graft
C0375265|ICD9CM|AB|414.05|Cor ath bypass graft NOS
C0375267|ICD9CM|PT|415.19|Other pulmonary embolism and infarction
C0375267|ICD9CM|AB|415.19|Pulm embol/infarct NEC
C0375268|ICD9CM|PT|421.9|Acute endocarditis, unspecified
C0375268|ICD9CM|AB|421.9|Ac/subac endocardit NOS
C0375273|ICD9CM|PT|433.00|Occlusion and stenosis of basilar artery without mention of cerebral infarction
C0375273|ICD9CM|AB|433.00|Ocl bslr art wo infrct
C0375274|ICD9CM|PT|433.01|Occlusion and stenosis of basilar artery with cerebral infarction
C0375274|ICD9CM|AB|433.01|Ocl bslr art w infrct
C0375275|ICD9CM|PT|433.10|Occlusion and stenosis of carotid artery without mention of cerebral infarction
C0375275|ICD9CM|AB|433.10|Ocl crtd art wo infrct
C0375276|ICD9CM|PT|433.11|Occlusion and stenosis of carotid artery with cerebral infarction
C0375276|ICD9CM|AB|433.11|Ocl crtd art w infrct
C0375277|ICD9CM|PT|433.20|Occlusion and stenosis of vertebral artery without mention of cerebral infarction
C0375277|ICD9CM|AB|433.20|Ocl vrtb art wo infrct
C0375278|ICD9CM|PT|433.21|Occlusion and stenosis of vertebral artery with cerebral infarction
C0375278|ICD9CM|AB|433.21|Ocl vrtb art w infrct
C0375279|ICD9CM|PT|433.30|Occlusion and stenosis of multiple and bilateral precerebral arteries without mention of cerebral infarction
C0375279|ICD9CM|AB|433.30|Ocl mlt bi art wo infrct
C0375280|ICD9CM|PT|433.31|Occlusion and stenosis of multiple and bilateral precerebral arteries with cerebral infarction
C0375280|ICD9CM|AB|433.31|Ocl mlt bi art w infrct
C0375281|ICD9CM|PT|433.80|Occlusion and stenosis of other specified precerebral artery without mention of cerebral infarction
C0375281|ICD9CM|AB|433.80|Ocl spcf art wo infrct
C0375282|ICD9CM|PT|433.81|Occlusion and stenosis of other specified precerebral artery with cerebral infarction
C0375282|ICD9CM|AB|433.81|Ocl spcf art w infrct
C0375283|ICD9CM|PT|433.90|Occlusion and stenosis of unspecified precerebral artery without mention of cerebral infarction
C0375283|ICD9CM|AB|433.90|Ocl art NOS wo infrct
C0375284|ICD9CM|PT|433.91|Occlusion and stenosis of unspecified precerebral artery with cerebral infarction
C0375284|ICD9CM|AB|433.91|Ocl art NOS w infrct
C0375285|ICD9CM|PT|434.00|Cerebral thrombosis without mention of cerebral infarction
C0375285|ICD9CM|AB|434.00|Crbl thrmbs wo infrct
C0375286|ICD9CM|PT|434.01|Cerebral thrombosis with cerebral infarction
C0375286|ICD9CM|AB|434.01|Crbl thrmbs w infrct
C0375287|ICD9CM|PT|434.10|Cerebral embolism without mention of cerebral infarction
C0375287|ICD9CM|AB|434.10|Crbl emblsm wo infrct
C0375288|ICD9CM|PT|434.11|Cerebral embolism with cerebral infarction
C0375288|ICD9CM|AB|434.11|Crbl emblsm w infrct
C0375290|ICD9CM|PT|434.90|Cerebral artery occlusion, unspecified without mention of cerebral infarction
C0375290|ICD9CM|AB|434.90|Crbl art oc NOS wo infrc
C0375291|ICD9CM|PT|434.91|Cerebral artery occlusion, unspecified with cerebral infarction
C0375291|ICD9CM|AB|434.91|Crbl art ocl NOS w infrc
C0375294|ICD9CM|PT|440.20|Atherosclerosis of native arteries of the extremities, unspecified
C0375294|ICD9CM|AB|440.20|Athscl extrm ntv art NOS
C0375295|ICD9CM|PT|440.21|Atherosclerosis of native arteries of the extremities with intermittent claudication
C0375295|ICD9CM|AB|440.21|Ath ext ntv at w claudct
C0375297|ICD9CM|PT|440.23|Atherosclerosis of native arteries of the extremities with ulceration
C0375297|ICD9CM|AB|440.23|Ath ext ntv art ulcrtion
C0375298|ICD9CM|PT|440.24|Atherosclerosis of native arteries of the extremities with gangrene
C0375298|ICD9CM|AB|440.24|Ath ext ntv art gngrene
C0375299|ICD9CM|PT|440.29|Other atherosclerosis of native arteries of the extremities
C0375299|ICD9CM|AB|440.29|Athrsc extrm ntv art oth
C0375300|ICD9CM|HT|440.3|Of bypass graft of the extremities
C0375301|ICD9CM|PT|440.30|Atherosclerosis of unspecified bypass graft of the extremities
C0375301|ICD9CM|AB|440.30|Athscl extrm bps gft NOS
C0375302|ICD9CM|PT|440.31|Atherosclerosis of autologous vein bypass graft of the extremities
C0375302|ICD9CM|AB|440.31|Ath ext autologs bps gft
C0375305|ICD9CM|PT|441.03|Dissection of aorta, thoracoabdominal
C0375305|ICD9CM|AB|441.03|Dsct of thoracoabd aorta
C0375306|ICD9CM|PT|441.7|Thoracoabdominal aneurysm, without mention of rupture
C0375306|ICD9CM|AB|441.7|Thracabd anurysm wo rupt
C0375311|ICD9CM|PT|451.82|Phlebitis and thrombophlebitis of superficial veins of upper extremities
C0375311|ICD9CM|AB|451.82|Phlbts sprfc vn up extrm
C0375312|ICD9CM|PT|451.83|Phlebitis and thrombophlebitis of deep veins of upper extremities
C0375312|ICD9CM|AB|451.83|Phlbts deep vn up extrm
C0375313|ICD9CM|PT|451.84|Phlebitis and thrombophlebitis of upper extremities, unspecified
C0375313|ICD9CM|AB|451.84|Phlbts vn NOS up extrm
C0375314|ICD9CM|HT|458.2|Iatrogenic hypotension
C0375319|ICD9CM|PT|466.19|Acute bronchiolitis due to other infectious organisms
C0375319|ICD9CM|AB|466.19|Acu brnchlts d/t oth org
C0375321|ICD9CM|PT|478.8|Upper respiratory tract hypersensitivity reaction, site unspecified
C0375321|ICD9CM|AB|478.8|Urt hypersens react NOS
C0375324|ICD9CM|PT|482.31|Pneumonia due to Streptococcus, group A
C0375324|ICD9CM|AB|482.31|Pneumonia strptococcus a
C0375326|ICD9CM|PT|482.39|Pneumonia due to other Streptococcus
C0375326|ICD9CM|AB|482.39|Pneumonia oth strep
C0375327|ICD9CM|PT|482.81|Pneumonia due to anaerobes
C0375327|ICD9CM|AB|482.81|Pneumonia anaerobes
C0375333|ICD9CM|PT|493.20|Chronic obstructive asthma, unspecified
C0375333|ICD9CM|AB|493.20|Chronic obst asthma NOS
C0375334|ICD9CM|PT|493.21|Chronic obstructive asthma with status asthmaticus
C0375334|ICD9CM|AB|493.21|Ch ob asthma w stat asth
C0375336|ICD9CM|AB|512.1|Iatrogenic pneumothorax
C0375336|ICD9CM|PT|512.1|Iatrogenic pneumothorax
C0375340|ICD9CM|PT|524.09|Major anomalies of jaw size, other specified anomaly
C0375340|ICD9CM|AB|524.09|Oth spcf anmly jaw size
C0375343|ICD9CM|AB|524.12|Other jaw asymmetry
C0375343|ICD9CM|PT|524.12|Anomalies of relationship of jaw to cranial base, other jaw asymmetry
C0375344|ICD9CM|PT|524.19|Anomalies of relationship of jaw to cranial base, other specified anomaly
C0375344|ICD9CM|AB|524.19|Spcfd anom jaw cranl bse
C0375346|ICD9CM|HT|524.7|Dental alveolar anomalies
C0375346|ICD9CM|PT|524.70|Dental alveolar anomalies, unspecified alveolar anomaly
C0375346|ICD9CM|AB|524.70|Unspf dent alvelr anmaly
C0375347|ICD9CM|PT|524.71|Alveolar maxillary hyperplasia
C0375347|ICD9CM|AB|524.71|Alveolar maxil hyprplsia
C0375348|ICD9CM|PT|524.72|Alveolar mandibular hyperplasia
C0375348|ICD9CM|AB|524.72|Alveolar mandib hyprplas
C0375349|ICD9CM|PT|524.73|Alveolar maxillary hypoplasia
C0375349|ICD9CM|AB|524.73|Alveolar maxil hypoplsia
C0375350|ICD9CM|PT|524.74|Alveolar mandibular hypoplasia
C0375350|ICD9CM|AB|524.74|Alveolar mandb hypoplsia
C0375352|ICD9CM|AB|530.19|Other esophagitis
C0375352|ICD9CM|PT|530.19|Other esophagitis
C0375354|ICD9CM|PT|550.02|Inguinal hernia, with gangrene, bilateral (not specified as recurrent)
C0375354|ICD9CM|AB|550.02|Bilat ing hernia w gang
C0375359|ICD9CM|PT|556.5|Left-sided ulcerative (chronic) colitis
C0375359|ICD9CM|AB|556.5|Lftsded ulcertve colitis
C0375360|ICD9CM|PT|556.6|Universal ulcerative (chronic) colitis
C0375360|ICD9CM|AB|556.6|Univrsl ulcertve colitis
C0375362|ICD9CM|PT|568.0|Peritoneal adhesions (postoperative) (postinfection)
C0375362|ICD9CM|AB|568.0|Peritoneal adhesions
C0375363|ICD9CM|PT|569.61|Infection of colostomy or enterostomy
C0375363|ICD9CM|AB|569.61|Colosty/enterost infectn
C0375364|ICD9CM|PT|569.69|Other colostomy and enterostomy complication
C0375364|ICD9CM|AB|569.69|Colstmy/enteros comp NEC
C0375365|ICD9CM|HT|574.6|Calculus of gallbladder and bile duct with acute cholecystitis
C0375366|ICD9CM|PT|574.60|Calculus of gallbladder and bile duct with acute cholecystitis, without mention of obstruction
C0375366|ICD9CM|AB|574.60|Gall&bil cal w/ac w/o ob
C0375367|ICD9CM|PT|574.61|Calculus of gallbladder and bile duct with acute cholecystitis, with obstruction
C0375367|ICD9CM|AB|574.61|Gall&bil cal w/ac w obs
C0375368|ICD9CM|HT|574.7|Calculus of gallbladder and bile duct with other cholecystitis
C0375369|ICD9CM|PT|574.70|Calculus of gallbladder and bile duct with other cholecystitis, without mention of obstruction
C0375369|ICD9CM|AB|574.70|Gal&bil cal w/oth w/o ob
C0375370|ICD9CM|PT|574.71|Calculus of gallbladder and bile duct with other cholecystitis, with obstruction
C0375370|ICD9CM|AB|574.71|Gall&bil cal w/oth w obs
C0375371|ICD9CM|HT|574.8|Calculus of gallbladder and bile duct with acute and chronic cholecystitis
C0375372|ICD9CM|PT|574.80|Calculus of gallbladder and bile duct with acute and chronic cholecystitis, without mention of obstruction
C0375372|ICD9CM|AB|574.80|Gal&bil cal w/ac&chr w/o
C0375373|ICD9CM|PT|574.81|Calculus of gallbladder and bile duct with acute and chronic cholecystitis, with obstruction
C0375373|ICD9CM|AB|574.81|Gal&bil cal w/ac&ch w ob
C0375374|ICD9CM|HT|574.9|Calculus of gallbladder and bile duct without cholecystitis
C0375375|ICD9CM|PT|574.90|Calculus of gallbladder and bile duct without cholecystitis, without mention of obstruction
C0375375|ICD9CM|AB|574.90|Gall&bil cal w/o cho w/o
C0375376|ICD9CM|PT|574.91|Calculus of gallbladder and bile duct without cholecystitis, with obstruction
C0375376|ICD9CM|AB|574.91|Gall&bil cal w/o ch w ob
C0375377|ICD9CM|PT|593.71|Vesicoureteral reflux with reflux nephropathy, unilateral
C0375377|ICD9CM|AB|593.71|Vscurt rflx npht uniltrl
C0375378|ICD9CM|PT|593.72|Vesicoureteral reflux with reflux nephropathy, bilateral
C0375378|ICD9CM|AB|593.72|Vscourtl rflx npht bltrl
C0375379|ICD9CM|PT|593.73|Other vesicoureteral reflux with reflux nephropathy NOS
C0375379|ICD9CM|AB|593.73|Vscourtl rflx w npht NOS
C0375380|ICD9CM|AB|599.81|Urethral hypermobility
C0375380|ICD9CM|PT|599.81|Urethral hypermobility
C0375381|ICD9CM|PT|599.82|Intrinsic (urethral) sphincter deficiency [ISD]
C0375381|ICD9CM|AB|599.82|Intrinsc sphnctr dficncy
C0375384|ICD9CM|PT|614.6|Pelvic peritoneal adhesions, female (postoperative) (postinfection)
C0375384|ICD9CM|AB|614.6|Fem pelvic periton adhes
C0375389|ICD9CM|PT|647.23|Other venereal diseases of mother, complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C0375389|ICD9CM|AB|647.23|Other vd-antepartum
C0375390|ICD9CM|PT|647.24|Other venereal diseases of mother, complicating pregnancy, childbirth, or the puerperium,postpartum condition or complication
C0375390|ICD9CM|AB|647.24|Other vd-postpartum
C0375391|ICD9CM|PT|652.30|Transverse or oblique presentation, unspecified as to episode of care or not applicable
C0375391|ICD9CM|AB|652.30|Transv/obliq lie-unspec
C0375392|ICD9CM|PT|652.31|Transverse or oblique presentation, delivered, with or without mention of antepartum condition
C0375392|ICD9CM|AB|652.31|Transver/obliq lie-deliv
C0375393|ICD9CM|PT|652.33|Transverse or oblique presentation, antepartum condition or complication
C0375393|ICD9CM|AB|652.33|Transv/obliq lie-antepar
C0375394|ICD9CM|HT|654.2|Previous cesarean section complicating pregnancy or childbirth
C0375395|ICD9CM|PT|654.21|Previous cesarean delivery, delivered, with or without mention of antepartum condition
C0375395|ICD9CM|AB|654.21|Prev c-delivery-delivrd
C0375434|ICD9CM|PT|657.01|Polyhydramnios, delivered, with or without mention of antepartum condition
C0375434|ICD9CM|AB|657.01|Polyhydramnios-delivered
C0375436|ICD9CM|PT|657.03|Polyhydramnios, antepartum condition or complication
C0375436|ICD9CM|AB|657.03|Polyhydramnios-antepart
C0375465|ICD9CM|PT|659.60|Elderly multigravida, unspecified as to episode of care or not applicable
C0375465|ICD9CM|AB|659.60|Elderly multigravida-uns
C0375466|ICD9CM|PT|659.61|Elderly multigravida, delivered with or without mention of antepartum condition
C0375466|ICD9CM|AB|659.61|Elderly multigravida-del
C0375468|ICD9CM|PT|659.63|Elderly multigravida, antepartum condition or complication
C0375468|ICD9CM|AB|659.63|Elderly multigravd-antep
C0375475|ICD9CM|PT|669.43|Other complications of obstetrical surgery and procedures, antepartum condition or complication
C0375475|ICD9CM|AB|669.43|Complc ob surg anteprtm
C0375476|ICD9CM|PT|670.00|Major puerperal infection, unspecified as to episode of care or not applicable
C0375476|ICD9CM|AB|670.00|Maj puerp inf NOS-unsp
C0375477|ICD9CM|PT|670.04|Major puerperal infection, postpartum condition or complication
C0375477|ICD9CM|AB|670.04|Major puerp inf NOS-p/p
C0375478|ICD9CM|PT|672.02|Pyrexia of unknown origin during the puerperium, delivered, with mention of postpartum complication
C0375478|ICD9CM|AB|672.02|Puerp pyrexia-del w p/p
C0375479|ICD9CM|PT|672.04|Pyrexia of unknown origin during the puerperium, postpartum condition or complication
C0375479|ICD9CM|AB|672.04|Puerp pyrexia-postpartum
C0375480|ICD9CM|PT|677|Late effect of complication of pregnancy, childbirth, and the puerperium
C0375480|ICD9CM|AB|677|Late effct cmplcatn preg
C0375481|ICD9CM|PT|690.8|Other erythematosquamous dermatosis
C0375481|ICD9CM|AB|690.8|Erythmtsquamous derm NEC
C0375482|ICD9CM|PT|692.72|Acute dermatitis due to solar radiation
C0375482|ICD9CM|AB|692.72|Act drmtitis solar rdiat
C0375483|ICD9CM|PT|692.73|Actinic reticuloid and actinic granuloma
C0375483|ICD9CM|AB|692.73|Actnc retic actnc grnlma
C0375484|ICD9CM|PT|692.74|Other chronic dermatitis due to solar radiation
C0375484|ICD9CM|AB|692.74|Oth chr drmtit solar rad
C0375485|ICD9CM|PT|692.79|Other dermatitis due to solar radiation
C0375485|ICD9CM|AB|692.79|Oth dermatitis solar rad
C0375486|ICD9CM|PT|692.82|Dermatitis due to other radiation
C0375486|ICD9CM|AB|692.82|Dermatitis oth radiation
C0375487|ICD9CM|PT|692.9|Contact dermatitis and other eczema, unspecified cause
C0375487|ICD9CM|AB|692.9|Dermatitis NOS
C0375488|ICD9CM|PT|702.19|Other seborrheic keratosis
C0375488|ICD9CM|AB|702.19|Other sborheic keratosis
C0375489|ICD9CM|AB|709.09|Other dyschromia
C0375489|ICD9CM|PT|709.09|Other dyschromia
C0375492|ICD9CM|PT|719.60|Other symptoms referable to joint, site unspecified
C0375492|ICD9CM|AB|719.60|Joint sympt NEC-unsp jt
C0375497|ICD9CM|PT|722.70|Intervertebral disc disorder with myelopathy, unspecified region
C0375497|ICD9CM|AB|722.70|Disc dis w myelopath NOS
C0375504|ICD9CM|PT|733.11|Pathologic fracture of humerus
C0375504|ICD9CM|AB|733.11|Path fx humerus
C0375505|ICD9CM|PT|733.12|Pathologic fracture of distal radius and ulna
C0375505|ICD9CM|AB|733.12|Path fx dstl radius ulna
C0375507|ICD9CM|PT|733.15|Pathologic fracture of other specified part of femur
C0375507|ICD9CM|AB|733.15|Path fx oth spcf prt fmr
C0375508|ICD9CM|PT|733.16|Pathologic fracture of tibia or fibula
C0375508|ICD9CM|AB|733.16|Path fx tibia fibula
C0375509|ICD9CM|PT|733.19|Pathologic fracture of other specified site
C0375509|ICD9CM|AB|733.19|Path fx oth specif site
C0375512|ICD9CM|AB|738.12|Zygomatic hypoplasia
C0375512|ICD9CM|PT|738.12|Zygomatic hypoplasia
C0375513|ICD9CM|PT|738.19|Other specified acquired deformity of head
C0375513|ICD9CM|AB|738.19|Oth spcf deformity head
C0375518|ICD9CM|AB|747.61|Gstrontest vesl anomaly
C0375518|ICD9CM|PT|747.61|Gastrointestinal vessel anomaly
C0375519|ICD9CM|AB|747.63|Upr limb vessel anomaly
C0375519|ICD9CM|PT|747.63|Upper limb vessel anomaly
C0375520|ICD9CM|AB|747.64|Lwr limb vessel anomaly
C0375520|ICD9CM|PT|747.64|Lower limb vessel anomaly
C0375521|ICD9CM|PT|747.69|Anomalies of other specified sites of peripheral vascular system
C0375521|ICD9CM|AB|747.69|Oth spcf prph vscl anoml
C0375522|ICD9CM|AB|747.82|Spinal vessel anomaly
C0375522|ICD9CM|PT|747.82|Spinal vessel anomaly
C0375526|ICD9CM|HT|752.6|Hypospadias and epispadias and other penile anomalies
C0375528|ICD9CM|PT|752.69|Other penile anomalies
C0375528|ICD9CM|AB|752.69|Penile anomalies NEC
C0375533|ICD9CM|PT|755.22|Longitudinal deficiency of upper limb, not elsewhere classified
C0375533|ICD9CM|AB|755.22|Longitud defic arm NEC
C0375534|ICD9CM|PT|755.32|Longitudinal deficiency of lower limb, not elsewhere classified
C0375534|ICD9CM|AB|755.32|Longitudin defic leg NEC
C0375536|ICD9CM|HT|756.5|Congenital osteodystrophies
C0375536|ICD9CM|AB|756.50|Osteodystrophy NOS
C0375536|ICD9CM|PT|756.50|Congenital osteodystrophy, unspecified
C0375539|ICD9CM|PT|760.76|Diethylstilbestrol [DES] affecting fetus or newborn via placenta or breast milk
C0375539|ICD9CM|AB|760.76|Maternal DES af NB/fetus
C0375543|ICD9CM|PT|774.30|Neonatal jaundice due to delayed conjugation, cause unspecified
C0375543|ICD9CM|AB|774.30|Delay conjugat jaund NOS
C0375546|ICD9CM|PT|785.2|Undiagnosed cardiac murmurs
C0375546|ICD9CM|AB|785.2|Cardiac murmurs NEC
C0375548|ICD9CM|AB|787.02|Nausea alone
C0375548|ICD9CM|PT|787.02|Nausea alone
C0375549|ICD9CM|PT|788.29|Other specified retention of urine
C0375549|ICD9CM|AB|788.29|Oth spcf retention urine
C0375551|ICD9CM|PT|788.34|Incontinence without sensory awareness
C0375551|ICD9CM|AB|788.34|Incontnce wo sensr aware
C0375552|ICD9CM|AB|788.35|Post-void dribbling
C0375552|ICD9CM|PT|788.35|Post-void dribbling
C0375553|ICD9CM|AB|788.37|Continuous leakage
C0375553|ICD9CM|PT|788.37|Continuous leakage
C0375554|ICD9CM|PT|788.39|Other urinary incontinence
C0375554|ICD9CM|AB|788.39|Oth urinry incontinence
C0375555|ICD9CM|PT|789.09|Abdominal pain, other specified site
C0375555|ICD9CM|AB|789.09|Abdmnal pain oth spcf st
C0375556|ICD9CM|PT|789.30|Abdominal or pelvic swelling, mass, or lump, unspecified site
C0375556|ICD9CM|AB|789.30|Abdmnal mass unspcf site
C0375557|ICD9CM|PT|789.31|Abdominal or pelvic swelling, mass, or lump, right upper quadrant
C0375557|ICD9CM|AB|789.31|Abdmnal mass rt upr quad
C0375558|ICD9CM|PT|789.32|Abdominal or pelvic swelling, mass, or lump, left upper quadrant
C0375558|ICD9CM|AB|789.32|Abdmnal mass lft up quad
C0375559|ICD9CM|PT|789.33|Abdominal or pelvic swelling, mass, or lump, right lower quadrant
C0375559|ICD9CM|AB|789.33|Abdmnal mass rt lwr quad
C0375560|ICD9CM|PT|789.34|Abdominal or pelvic swelling, mass, or lump, left lower quadrant
C0375560|ICD9CM|AB|789.34|Abdmnal mass lt lwr quad
C0375561|ICD9CM|PT|789.35|Abdominal or pelvic swelling, mass, or lump, periumbilic
C0375561|ICD9CM|AB|789.35|Abdmnal mass periumbilic
C0375562|ICD9CM|PT|789.36|Abdominal or pelvic swelling, mass, or lump, epigastric
C0375562|ICD9CM|AB|789.36|Abdmnal mass epigastric
C0375563|ICD9CM|PT|789.37|Abdominal or pelvic swelling, mass, or lump, generalized
C0375563|ICD9CM|AB|789.37|Abdmnal mass generalized
C0375564|ICD9CM|PT|789.39|Abdominal or pelvic swelling, mass, or lump, other specified site
C0375564|ICD9CM|AB|789.39|Abdmnal mass oth spcf st
C0375565|ICD9CM|PT|789.41|Abdominal rigidity, right upper quadrant
C0375565|ICD9CM|AB|789.41|Abdmnal rgdt rt upr quad
C0375570|ICD9CM|PT|789.46|Abdominal rigidity, epigastric
C0375570|ICD9CM|AB|789.46|Abdmnal rgdt epigastric
C0375571|ICD9CM|PT|789.47|Abdominal rigidity, generalized
C0375571|ICD9CM|AB|789.47|Abdmnal rgdt generalized
C0375572|ICD9CM|PT|789.49|Abdominal rigidity, other specified site
C0375572|ICD9CM|AB|789.49|Abdmnal rgdt oth spcf st
C0375573|ICD9CM|PT|789.65|Abdominal tenderness, periumbilic
C0375573|ICD9CM|AB|789.65|Abdmnal tndr periumbilic
C0375574|ICD9CM|PT|789.69|Abdominal tenderness, other specified site
C0375574|ICD9CM|AB|789.69|Abdmnal tndr oth spcf st
C0375575|ICD9CM|PT|790.91|Abnormal arterial blood gases
C0375575|ICD9CM|AB|790.91|Abnrml art blood gases
C0375576|ICD9CM|PT|790.92|Abnormal coagulation profile
C0375576|ICD9CM|AB|790.92|Abnrml coagultion prfile
C0375579|ICD9CM|PT|795.71|Nonspecific serologic evidence of human immunodeficiency virus [HIV]
C0375579|ICD9CM|AB|795.71|Nonspcf serlgc evdnc hiv
C0375580|ICD9CM|PT|795.79|Other and unspecified nonspecific immunological findings
C0375580|ICD9CM|HT|795.7|Other nonspecific immunological findings
C0375580|ICD9CM|AB|795.79|Oth unspcf nspf imun fnd
C0375581|ICD9CM|PT|800.19|Closed fracture of vault of skull with cerebral laceration and contusion, with concussion, unspecified
C0375581|ICD9CM|AB|800.19|Cl skl vlt fx-concus NOS
C0375582|ICD9CM|PT|800.29|Closed fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with concussion, unspecified
C0375582|ICD9CM|AB|800.29|Cl skl vlt fx-concus NOS
C0375583|ICD9CM|PT|800.39|Closed fracture of vault of skull with other and unspecified intracranial hemorrhage, with concussion, unspecified
C0375583|ICD9CM|AB|800.39|Cl skl vlt fx-concus NOS
C0375585|ICD9CM|PT|800.69|Open fracture of vault of skull with cerebral laceration and contusion, with concussion, unspecified
C0375585|ICD9CM|AB|800.69|Op skl vlt fx-concus NOS
C0375586|ICD9CM|PT|800.79|Open fracture of vault of skull with subarachnoid, subdural, and extradural hemorrhage, with concussion, unspecified
C0375586|ICD9CM|AB|800.79|Op skl vlt fx-concus NOS
C0375587|ICD9CM|PT|800.89|Open fracture of vault of skull with other and unspecified intracranial hemorrhage, with concussion, unspecified
C0375587|ICD9CM|AB|800.89|Op skl vlt fx-concus NOS
C0375589|ICD9CM|PT|801.19|Closed fracture of base of skull with cerebral laceration and contusion, with concussion, unspecified
C0375589|ICD9CM|AB|801.19|Cl skull base fx-concuss
C0375590|ICD9CM|PT|801.29|Closed fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with concussion, unspecified
C0375590|ICD9CM|AB|801.29|Cl skull base fx-concuss
C0375591|ICD9CM|PT|801.39|Closed fracture of base of skull with other and unspecified intracranial hemorrhage, with concussion, unspecified
C0375591|ICD9CM|AB|801.39|Cl skull base fx-concuss
C0375593|ICD9CM|PT|801.69|Open fracture of base of skull with cerebral laceration and contusion, with concussion, unspecified
C0375593|ICD9CM|AB|801.69|Opn skul base fx-concuss
C0375594|ICD9CM|PT|801.79|Open fracture of base of skull with subarachnoid, subdural, and extradural hemorrhage, with concussion, unspecified
C0375594|ICD9CM|AB|801.79|Opn skul base fx-concuss
C0375595|ICD9CM|PT|801.89|Open fracture of base of skull with other and unspecified intracranial hemorrhage, with concussion, unspecified
C0375595|ICD9CM|AB|801.89|Opn skul base fx-concuss
C0375598|ICD9CM|PT|803.19|Other closed skull fracture with cerebral laceration and contusion, with concussion, unspecified
C0375598|ICD9CM|AB|803.19|Cl skull fx NEC-concuss
C0375599|ICD9CM|PT|803.29|Other closed skull fracture with subarachnoid, subdural, and extradural hemorrhage, with concussion, unspecified
C0375599|ICD9CM|AB|803.29|Cl skull fx NEC-concuss
C0375600|ICD9CM|PT|803.39|Other closed skull fracture with other and unspecified intracranial hemorrhage, with concussion, unspecified
C0375600|ICD9CM|AB|803.39|Cl skull fx NEC-concuss
C0375603|ICD9CM|PT|803.69|Other open skull fracture with cerebral laceration and contusion, with concussion, unspecified
C0375603|ICD9CM|AB|803.69|Opn skull fx NEC-concuss
C0375604|ICD9CM|PT|803.79|Other open skull fracture with subarachnoid, subdural, and extradural hemorrhage, with concussion, unspecified
C0375604|ICD9CM|AB|803.79|Opn skull fx NEC-concuss
C0375605|ICD9CM|PT|803.89|Other open skull fracture with other and unspecified intracranial hemorrhage, with concussion, unspecified
C0375605|ICD9CM|AB|803.89|Opn skull fx NEC-concuss
C0375608|ICD9CM|PT|804.19|Closed fractures involving skull or face with other bones, with cerebral laceration and contusion, with concussion, unspecified
C0375608|ICD9CM|AB|804.19|Cl skul w oth fx-concuss
C0375609|ICD9CM|PT|804.29|Closed fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with concussion, unspecified
C0375609|ICD9CM|AB|804.29|Cl skul w oth fx-concuss
C0375610|ICD9CM|PT|804.39|Closed fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with concussion, unspecified
C0375610|ICD9CM|AB|804.39|Cl skul w oth fx-concuss
C0375613|ICD9CM|PT|804.69|Open fractures involving skull or face with other bones, with cerebral laceration and contusion, with concussion, unspecified
C0375613|ICD9CM|AB|804.69|Opn skull/oth fx-concuss
C0375614|ICD9CM|PT|804.79|Open fractures involving skull or face with other bones with subarachnoid, subdural, and extradural hemorrhage, with concussion, unspecified
C0375614|ICD9CM|AB|804.79|Opn skull/oth fx-concuss
C0375615|ICD9CM|PT|804.89|Open fractures involving skull or face with other bones, with other and unspecified intracranial hemorrhage, with concussion, unspecified
C0375615|ICD9CM|AB|804.89|Opn skull/oth fx-concuss
C0375617|ICD9CM|PT|805.00|Closed fracture of cervical vertebra, unspecified level
C0375617|ICD9CM|AB|805.00|Fx cervical vert NOS-cl
C0375618|ICD9CM|PT|805.10|Open fracture of cervical vertebra, unspecified level
C0375618|ICD9CM|AB|805.10|Fx cervical vert NOS-opn
C0375623|ICD9CM|PT|813.00|Closed fracture of upper end of forearm, unspecified
C0375623|ICD9CM|AB|813.00|Fx upper forearm NOS-cl
C0375624|ICD9CM|PT|813.10|Open fracture of upper end of forearm, unspecified
C0375624|ICD9CM|AB|813.10|Fx upper forearm NOS-opn
C0375625|ICD9CM|PT|831.00|Closed dislocation of shoulder, unspecified
C0375625|ICD9CM|AB|831.00|Disloc shoulder NOS-clos
C0375626|ICD9CM|PT|831.10|Open dislocation of shoulder, unspecified
C0375626|ICD9CM|AB|831.10|Disloc shoulder NOS-open
C0375627|ICD9CM|PT|832.00|Closed dislocation of elbow, unspecified
C0375627|ICD9CM|AB|832.00|Dislocat elbow NOS-close
C0375629|ICD9CM|PT|833.10|Open dislocation of wrist, unspecified part
C0375629|ICD9CM|AB|833.10|Dislocat wrist NOS-open
C0375630|ICD9CM|PT|834.00|Closed dislocation of finger, unspecified part
C0375630|ICD9CM|AB|834.00|Disl finger NOS-closed
C0375631|ICD9CM|PT|834.10|Open dislocation of finger, unspecified part
C0375631|ICD9CM|AB|834.10|Disloc finger NOS-open
C0375632|ICD9CM|PT|835.00|Closed dislocation of hip, unspecified site
C0375632|ICD9CM|AB|835.00|Dislocat hip NOS-closed
C0375633|ICD9CM|PT|835.10|Open dislocation of hip, unspecified site
C0375633|ICD9CM|AB|835.10|Dislocation hip NOS-open
C0375634|ICD9CM|PT|836.50|Dislocation of knee, unspecified, closed
C0375634|ICD9CM|AB|836.50|Dislocat knee NOS-closed
C0375635|ICD9CM|PT|838.00|Closed dislocation of foot, unspecified
C0375635|ICD9CM|AB|838.00|Dislocat foot NOS-closed
C0375636|ICD9CM|PT|838.10|Open dislocation of foot, unspecified
C0375636|ICD9CM|AB|838.10|Dislocat foot NOS-open
C0375639|ICD9CM|PT|864.05|Injury to liver without mention of open wound into cavity laceration, unspecified
C0375639|ICD9CM|AB|864.05|Liver lacerat unspcf cls
C0375641|ICD9CM|PT|872.00|Open wound of external ear, unspecified site, without mention of complication
C0375641|ICD9CM|AB|872.00|Opn wound extern ear NOS
C0375643|ICD9CM|PT|872.02|Open wound of auditory canal, without mention of complication
C0375643|ICD9CM|AB|872.02|Opn wound auditory canal
C0375646|ICD9CM|PT|872.63|Open wound of eustachian tube, without mention of complication
C0375646|ICD9CM|AB|872.63|Open wnd eustachian tube
C0375650|ICD9CM|PT|873.21|Open wound of nasal septum, without mention of complication
C0375650|ICD9CM|AB|873.21|Open wound nasal septum
C0375653|ICD9CM|PT|873.29|Open wound of multiple sites of nose, without mention of complication
C0375653|ICD9CM|AB|873.29|Mult open wound nose
C0375654|ICD9CM|PT|873.40|Open wound of face, unspecified site, without mention of complication
C0375654|ICD9CM|AB|873.40|Open wound of face NOS
C0375659|ICD9CM|PT|873.60|Open wound of mouth, unspecified site, without mention of complication
C0375659|ICD9CM|AB|873.60|Open wound of mouth NOS
C0375662|ICD9CM|PT|873.63|Open wound of tooth (broken) (fractured) (due to trauma), without mention of complication
C0375662|ICD9CM|AB|873.63|Broken tooth-uncomplic
C0375663|ICD9CM|PT|873.64|Open wound of tongue and floor of mouth, without mention of complication
C0375663|ICD9CM|AB|873.64|Opn wnd tongue/mouth flr
C0375668|ICD9CM|PT|909.5|Late effect of adverse effect of drug, medicinal or biological substance
C0375668|ICD9CM|AB|909.5|Lte efct advrs efct drug
C0375669|ICD9CM|PT|925.1|Crushing injury of face and scalp
C0375669|ICD9CM|AB|925.1|Crush inj face scalp
C0375673|ICD9CM|PT|941.16|Erythema [first degree] of scalp [any part]
C0375673|ICD9CM|AB|941.16|1st deg burn scalp
C0375674|ICD9CM|PT|941.20|Blisters, epidermal loss [second degree] of face and head, unspecified site
C0375674|ICD9CM|AB|941.20|2nd deg burn head NOS
C0375675|ICD9CM|PT|942.43|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of abdominal wall
C0375675|ICD9CM|AB|942.43|Deep 3rd burn abdom wall
C0375676|ICD9CM|PT|942.44|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of back [any part]
C0375676|ICD9CM|AB|942.44|Deep 3rd deg burn back
C0375677|ICD9CM|PT|942.45|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of genitalia
C0375677|ICD9CM|AB|942.45|Deep 3rd burn genitalia
C0375678|ICD9CM|PT|942.53|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of abdominal wall
C0375678|ICD9CM|AB|942.53|3rd brn w loss-abdom wll
C0375679|ICD9CM|PT|942.54|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of back [any part]
C0375679|ICD9CM|AB|942.54|3rd deg burn w loss-back
C0375680|ICD9CM|PT|942.55|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of genitalia
C0375680|ICD9CM|AB|942.55|3rd brn w loss-genitalia
C0375681|ICD9CM|HT|943.0|Burn of upper limb, except wrist and hand, unspecified degree
C0375683|ICD9CM|PT|945.41|Deep necrosis of underlying tissues [deep third degree] without mention of loss of a body part, of toe(s)(nail)
C0375683|ICD9CM|AB|945.41|Deep 3rd deg burn toe
C0375684|ICD9CM|PT|945.51|Deep necrosis of underlying tissues [deep third degree] with loss of a body part, of toe(s) (nail)
C0375684|ICD9CM|AB|945.51|3 deg burn w loss-toe
C0375688|ICD9CM|PT|949.3|Full-thickness skin loss [third degree nos]
C0375688|ICD9CM|AB|949.3|3rd degree burn NOS
C0375691|ICD9CM|PT|983.9|Toxic effect of caustic, unspecified
C0375691|ICD9CM|AB|983.9|Toxic effect caustic NOS
C0375692|ICD9CM|AB|989.81|Toxic effect of asbestos
C0375692|ICD9CM|PT|989.81|Toxic effect of asbestos
C0375693|ICD9CM|AB|989.82|Toxic effect of latex
C0375693|ICD9CM|PT|989.82|Toxic effect of latex
C0375694|ICD9CM|AB|989.83|Toxic effect of silicone
C0375694|ICD9CM|PT|989.83|Toxic effect of silicone
C0375695|ICD9CM|AB|989.84|Toxic effect of tobacco
C0375695|ICD9CM|PT|989.84|Toxic effect of tobacco
C0375699|ICD9CM|PT|995.51|Child emotional/psychological abuse
C0375699|ICD9CM|AB|995.51|Child emotnl/psych abuse
C0375700|ICD9CM|PT|995.52|Child neglect (nutritional)
C0375700|ICD9CM|AB|995.52|Child neglect-nutrition
C0375702|ICD9CM|PT|995.59|Other child abuse and neglect
C0375702|ICD9CM|AB|995.59|Child abuse/neglect NEC
C0375703|ICD9CM|PT|995.60|Anaphylactic reaction due to unspecified food
C0375703|ICD9CM|AB|995.60|Anphylct react food NOS
C0375707|ICD9CM|PT|995.64|Anaphylactic reaction due to tree nuts and seeds
C0375707|ICD9CM|AB|995.64|Anphyl react tr nts seed
C0375714|ICD9CM|PT|995.80|Adult maltreatment, unspecified
C0375714|ICD9CM|AB|995.80|Adult maltreatment NOS
C0375715|ICD9CM|PT|995.82|Adult emotional/psychological abuse
C0375715|ICD9CM|AB|995.82|Adult emotnl/psych abuse
C0375716|ICD9CM|PT|995.84|Adult neglect (nutritional)
C0375716|ICD9CM|AB|995.84|Adult neglect-nutrition
C0375717|ICD9CM|PT|995.85|Other adult abuse and neglect
C0375717|ICD9CM|AB|995.85|Oth adult abuse/neglect
C0375718|ICD9CM|PT|996.04|Mechanical complication of automatic implantable cardiac defibrillator
C0375718|ICD9CM|AB|996.04|Mch cmp autm mplnt dfbrl
C0375720|ICD9CM|PT|996.80|Complications of transplanted organ, unspecified
C0375720|ICD9CM|AB|996.80|Comp organ transplnt NOS
C0375722|ICD9CM|PT|997.02|Iatrogenic cerebrovascular infarction or hemorrhage
C0375722|ICD9CM|AB|997.02|Iatrogen CV infarc/hmrhg
C0375723|ICD9CM|PT|997.09|Other nervous system complications
C0375723|ICD9CM|AB|997.09|Surg comp nerv systm NEC
C0375724|MTH|PN|NOCODE|Other complications affecting other specified body systems, NEC in ICD9CM
C0375724|ICD9CM|PT|997.99|Complications affecting other specified body systems, not elsewhere classified
C0375724|ICD9CM|AB|997.99|Surg compl-body syst NEC
C0375725|ICD9CM|PT|998.11|Hemorrhage complicating a procedure
C0375725|ICD9CM|AB|998.11|Hemorrhage complic proc
C0375726|ICD9CM|PT|998.12|Hematoma complicating a procedure
C0375726|ICD9CM|AB|998.12|Hematoma complic proc
C0375727|ICD9CM|PT|998.13|Seroma complicating a procedure
C0375727|ICD9CM|AB|998.13|Seroma complicting proc
C0375728|ICD9CM|PT|998.51|Infected postoperative seroma
C0375728|ICD9CM|AB|998.51|Infected postop seroma
C0375729|ICD9CM|PT|998.59|Other postoperative infection
C0375729|ICD9CM|AB|998.59|Other postop infection
C0375731|ICD9CM|PT|998.82|Cataract fragments in eye following cataract surgery
C0375731|ICD9CM|AB|998.82|Ctrct frgmt frm ctr surg
C0375732|ICD9CM|PT|998.83|Non-healing surgical wound
C0375732|ICD9CM|AB|998.83|Non-healing surgcl wound
C0375733|ICD9CM|HT|E865|Accidental poisoning from poisonous foodstuffs and poisonous plants
C0375734|ICD9CM|PT|E869.4|Second hand tobacco smoke
C0375734|ICD9CM|AB|E869.4|Scndhnd tbcco smoke
C0375735|ICD9CM|PT|E880.1|Accidental fall on or from sidewalk curb
C0375735|ICD9CM|AB|E880.1|Fall on sidewalk curb
C0375736|ICD9CM|PT|E884.5|Accidental fall from other furniture
C0375736|ICD9CM|AB|E884.5|Fall from furniture NEC
C0375737|ICD9CM|PT|E884.6|Accidental fall from commode
C0375737|ICD9CM|AB|E884.6|Fall from commode
C0375739|ICD9CM|PT|E908.0|Hurricane
C0375739|ICD9CM|AB|E908.0|Accident d/t hurricane
C0375740|ICD9CM|PT|E908.1|Tornado
C0375740|ICD9CM|AB|E908.1|Accident d/t tornado
C0375741|ICD9CM|PT|E908.2|Floods
C0375741|ICD9CM|AB|E908.2|Accident d/t floods
C0375742|ICD9CM|PT|E908.3|Blizzard (snow) (ice)
C0375742|ICD9CM|AB|E908.3|Acc d/t snow blizzard
C0375743|ICD9CM|AB|E908.4|Accident d/t dust storm
C0375743|ICD9CM|PT|E908.4|Dust storm
C0375744|ICD9CM|AB|E908.8|Accident d/t storm NEC
C0375744|ICD9CM|PT|E908.8|Other cataclysmic storms
C0375746|ICD9CM|PT|E909.1|Volcanic eruptions
C0375746|ICD9CM|AB|E909.1|Acc d/t volcanic erupt
C0375747|ICD9CM|AB|E909.2|Acc d/t avalanche
C0375747|ICD9CM|PT|E909.2|Avalanche, landslide, or mudslide
C0375748|ICD9CM|PT|E909.3|Collapse of dam or man-made structure
C0375748|ICD9CM|AB|E909.3|Acc d/t dam collapse
C0375750|ICD9CM|PT|E909.8|Other cataclysmic earth surface movements and eruptions
C0375750|ICD9CM|AB|E909.8|Acc d/t eruptions NEC
C0375751|ICD9CM|PT|E909.9|Unspecified cataclysmic earth surface movements and eruptions
C0375751|ICD9CM|AB|E909.9|Acc d/t eruptions NOS
C0375752|ICD9CM|PT|E920.5|Accidents caused by hypodermic needle
C0375752|ICD9CM|AB|E920.5|Acc-hypodermic needle
C0375753|ICD9CM|PT|E924.2|Accident caused by hot (boiling) tap water
C0375753|ICD9CM|AB|E924.2|Acc-hot tap water
C0375754|ICD9CM|PT|E955.9|Suicide and self-inflicted injury by firearms and explosives, unspecified
C0375754|ICD9CM|AB|E955.9|Injury-firearm/expl NOS
C0375757|ICD9CM|PT|E967.3|Perpetrator of child and adult abuse, by spouse or partner
C0375757|ICD9CM|AB|E967.3|Batter by spouse/partner
C0375758|ICD9CM|PT|E967.4|Perpetrator of child and adult abuse, by child
C0375758|ICD9CM|AB|E967.4|Battering by child
C0375759|ICD9CM|PT|E967.5|Perpetrator of child and adult abuse, by sibling
C0375759|ICD9CM|AB|E967.5|Battering by sibling
C0375760|ICD9CM|PT|E967.6|Perpetrator of child and adult abuse, by grandparent
C0375760|ICD9CM|AB|E967.6|Battering by grandparent
C0375761|ICD9CM|PT|E967.7|Perpetrator of child and adult abuse, by other relative
C0375761|ICD9CM|AB|E967.7|Batter by other relative
C0375762|ICD9CM|PT|E967.8|Perpetrator of child and adult abuse, by non-related caregiver
C0375762|ICD9CM|AB|E967.8|Batter by non-relative
C0375763|ICD9CM|AB|E967.9|Child abuse NOS
C0375763|ICD9CM|PT|E967.9|Perpetrator of child and adult abuse, by unspecified person
C0375764|ICD9CM|PT|E968.5|Assault by transport vehicle
C0375764|ICD9CM|AB|E968.5|Asslt-transport vehicle
C0375765|ICD9CM|PT|V03.81|Other specified vaccinations against hemophilus influenza, type B [Hib]
C0375765|ICD9CM|AB|V03.81|Nd vac hmophlus inflnz b
C0375766|ICD9CM|PT|V03.82|Other specified vaccinations against streptococcus pneumoniae [pneumococcus]
C0375766|ICD9CM|AB|V03.82|Nd vac strptcs pneumni b
C0375767|ICD9CM|HT|V04|Need for prophylactic vaccination and inoculation against certain diseases
C0375768|ICD9CM|HT|V05|Need for prophylactic vaccination and inoculation against single diseases
C0375770|ICD9CM|PT|V05.4|Need for prophylactic vaccination and inoculation against varicella
C0375770|ICD9CM|AB|V05.4|Need prphyl vc varicella
C0375771|ICD9CM|PT|V06.5|Need for prophylactic vaccination and inoculation against tetanus-diphtheria [Td] (DT)
C0375771|ICD9CM|AB|V06.5|Vaccination for Td-DT
C0375772|ICD9CM|PT|V06.6|Need for prophylactic vaccination and inoculation against streptococcus pneumoniae [pneumococcus] and influenza
C0375772|ICD9CM|AB|V06.6|Nd vac strp pnumn/inflnz
C0375773|ICD9CM|PT|V07.31|Need for prophylactic fluoride administration
C0375773|ICD9CM|AB|V07.31|Prophylac fluoride admin
C0375777|ICD9CM|PT|V09.0|Infection with microorganisms resistant to penicillins
C0375777|ICD9CM|AB|V09.0|Inf mcrg rstn pncllins
C0375778|ICD9CM|PT|V09.1|Infection with microorganisms resistant to cephalosporins and other B-lactam antibiotics
C0375778|ICD9CM|AB|V09.1|Inf mcrg rstn b-lactam
C0375779|ICD9CM|PT|V09.2|Infection with microorganisms resistant to macrolides
C0375779|ICD9CM|AB|V09.2|Inf mcrg rstn macrolides
C0375780|ICD9CM|PT|V09.3|Infection with microorganisms resistant to tetracyclines
C0375780|ICD9CM|AB|V09.3|Inf mcrg rstn ttrcycln
C0375781|ICD9CM|PT|V09.4|Infection with microorganisms resistant to aminoglycosides
C0375781|ICD9CM|AB|V09.4|Inf mcrg rstn amnglcsds
C0375782|ICD9CM|HT|V09.5|Infection with microorganisms resistant to quinolones and fluoroquinolones
C0375783|ICD9CM|PT|V09.50|Infection with microorganisms without mention of resistance to multiple quinolones and fluroquinolones
C0375783|ICD9CM|AB|V09.50|Inf mcr rst qn flr nt ml
C0375784|ICD9CM|PT|V09.51|Infection with microorganisms with resistance to multiple quinolones and fluroquinolones
C0375784|ICD9CM|AB|V09.51|Inf mcrg rstn qn flrq ml
C0375785|ICD9CM|PT|V09.6|Infection with microorganisms resistant to sulfonamides
C0375785|ICD9CM|AB|V09.6|Inf mcrg rstn sulfnmides
C0375786|ICD9CM|HT|V09.7|Infection with microorganisms resistant to other specified antimycobacterial agents
C0375787|ICD9CM|PT|V09.70|Infection with microorganisms without mention of resistance to multiple antimycobacterial agents
C0375787|ICD9CM|AB|V09.70|Inf mcr rst oth ag nt ml
C0375788|ICD9CM|PT|V09.71|Infection with microorganisms with resistance to multiple antimycobacterial agents
C0375788|ICD9CM|AB|V09.71|Inf mcrg rstn oth ag mlt
C0375789|ICD9CM|HT|V09.8|Infection with microorganisms resistant to other specified drugs
C0375790|ICD9CM|PT|V09.80|Infection with microorganisms without mention of resistance to multiple drugs
C0375790|ICD9CM|AB|V09.80|Inf mcr rst ot drg nt ml
C0375791|ICD9CM|PT|V09.81|Infection with microorganisms with resistance to multiple drugs
C0375791|ICD9CM|AB|V09.81|Inf mcrg rstn oth drg ml
C0375792|ICD9CM|HT|V09|Infection with drug-resistant microorganisms
C0375792|ICD9CM|HT|V09.9|Infection with drug-resistant microorganisms, unspecified
C0375793|ICD9CM|PT|V09.90|Infection with drug-resistant microorganisms, unspecified, without mention of multiple drug resistance
C0375793|ICD9CM|AB|V09.90|Infc mcrg drgrst nt mult
C0375794|ICD9CM|PT|V09.91|Infection with drug-resistant microorganisms, unspecified, with multiple drug resistance
C0375794|ICD9CM|AB|V09.91|Infc mcrg drgrst mult
C0375795|ICD9CM|PT|V12.00|Personal history of unspecified infectious and parasitic disease
C0375795|ICD9CM|AB|V12.00|Prsnl hst unsp nfct prst
C0375796|ICD9CM|PT|V12.01|Personal history of tuberculosis
C0375796|ICD9CM|AB|V12.01|Prsnl hst tuberculosis
C0375797|ICD9CM|PT|V12.02|Personal history of poliomyelitis
C0375797|ICD9CM|AB|V12.02|Prsnl hst poliomyelitis
C0375798|ICD9CM|PT|V12.03|Personal history of malaria
C0375798|ICD9CM|AB|V12.03|Personal histry malaria
C0375799|ICD9CM|PT|V12.09|Personal history of other infectious and parasitic diseases
C0375799|ICD9CM|AB|V12.09|Prsnl hst oth nfct parst
C0375800|ICD9CM|PT|V12.51|Personal history of venous thrombosis and embolism
C0375800|ICD9CM|AB|V12.51|Hx-ven thrombosis/embols
C0375801|ICD9CM|PT|V12.52|Personal history of thrombophlebitis
C0375801|ICD9CM|AB|V12.52|Hx-thrombophlebitis
C0375802|ICD9CM|PT|V12.59|Personal history of other diseases of circulatory system
C0375802|ICD9CM|AB|V12.59|Hx-circulatory dis NEC
C0375803|ICD9CM|PT|V12.71|Personal history of peptic ulcer disease
C0375803|ICD9CM|AB|V12.71|Prsnl hst peptic ulcr ds
C0375804|ICD9CM|PT|V12.72|Personal history of colonic polyps
C0375804|ICD9CM|AB|V12.72|Prsnl hst colonic polyps
C0375805|ICD9CM|PT|V12.79|Personal history of other diseases of digestive system
C0375805|ICD9CM|AB|V12.79|Prsnl hst ot spf dgst ds
C0375806|ICD9CM|PT|V13.01|Personal history of urinary calculi
C0375806|ICD9CM|AB|V13.01|Prsnl hst urnr dsrd calc
C0375807|ICD9CM|PT|V13.09|Personal history of other specified urinary system disorders
C0375807|ICD9CM|AB|V13.09|Prsn hst ot spf urn dsrd
C0375810|ICD9CM|PT|V15.49|Other psychological trauma
C0375810|ICD9CM|AB|V15.49|Psychological trauma NEC
C0375815|ICD9CM|PT|V25.9|Unspecified contraceptive management
C0375815|ICD9CM|HT|V25|Encounter for contraceptive management
C0375815|ICD9CM|AB|V25.9|Contraceptive mangmt NOS
C0375816|ICD9CM|HT|V25.0|Encounter for general counseling and advice on contraceptive management
C0375817|ICD9CM|PT|V25.01|General counseling on prescription of oral contraceptives
C0375817|ICD9CM|AB|V25.01|Prescrip-oral contracept
C0375818|ICD9CM|PT|V25.02|General counseling on initiation of other contraceptive measures
C0375818|ICD9CM|AB|V25.02|Initiate contracept NEC
C0375820|ICD9CM|PT|V25.11|Encounter for insertion of intrauterine contraceptive device
C0375820|ICD9CM|AB|V25.11|Insertion of iud
C0375823|ICD9CM|HT|V25.4|Encounter for surveillance of previously prescribed contraceptive methods
C0375824|ICD9CM|PT|V25.40|Contraceptive surveillance, unspecified
C0375824|ICD9CM|AB|V25.40|Contracept surveill NOS
C0375825|ICD9CM|PT|V25.41|Surveillance of contraceptive pill
C0375825|ICD9CM|AB|V25.41|Contracept pill surveill
C0375827|ICD9CM|PT|V25.43|Surveillance of implantable subdermal contraceptive
C0375827|ICD9CM|AB|V25.43|Srvl mplnt sbdrm cntrcep
C0375828|ICD9CM|PT|V25.49|Surveillance of other contraceptive method
C0375828|ICD9CM|AB|V25.49|Contracept surveill NEC
C0375829|ICD9CM|PT|V25.5|Insertion of implantable subdermal contraceptive
C0375829|ICD9CM|AB|V25.5|Nsrt mplnt sbdrm cntrcep
C0375832|ICD9CM|HT|V29|Observation and evaluation of newborns for suspected condition not found
C0375833|ICD9CM|PT|V29.0|Observation for suspected infectious condition
C0375833|ICD9CM|AB|V29.0|NB obsrv suspct infect
C0375834|ICD9CM|PT|V29.1|Observation for suspected neurological conditions
C0375834|ICD9CM|AB|V29.1|NB obsrv suspct neurlgcl
C0375835|ICD9CM|PT|V29.2|Observation and evaluation of newborn for suspected respiratory condition
C0375835|ICD9CM|AB|V29.2|Obsrv NB suspc resp cond
C0375836|ICD9CM|PT|V43.60|Unspecified joint replacement
C0375836|ICD9CM|AB|V43.60|Joint replaced unspcf
C0375838|ICD9CM|PT|V43.62|Elbow joint replacement
C0375838|ICD9CM|AB|V43.62|Joint replaced elbow
C0375839|ICD9CM|AB|V43.63|Joint replaced wrist
C0375839|ICD9CM|PT|V43.63|Wrist joint replacement
C0375841|ICD9CM|PT|V43.65|Knee joint replacement
C0375841|ICD9CM|AB|V43.65|Joint replaced knee
C0375842|ICD9CM|PT|V43.66|Ankle joint replacement
C0375842|ICD9CM|AB|V43.66|Joint replaced ankle
C0375843|ICD9CM|PT|V43.69|Other joint replacement
C0375843|ICD9CM|AB|V43.69|Oth spcf joint replaced
C0375844|ICD9CM|AB|V43.81|Larynx replacement
C0375844|ICD9CM|PT|V43.81|Larynx replacement
C0375845|ICD9CM|AB|V43.82|Breast replacement
C0375845|ICD9CM|PT|V43.82|Breast replacement
C0375846|ICD9CM|PT|V45.00|Unspecified cardiac device in situ
C0375846|ICD9CM|AB|V45.00|Status cardc dvce unspcf
C0375848|ICD9CM|PT|V45.09|Other specified cardiac device in situ
C0375848|ICD9CM|AB|V45.09|Status oth spcf crdc dvc
C0375849|ICD9CM|HT|V45.5|Presence of contraceptive device
C0375850|ICD9CM|PT|V45.52|Presence of subdermal contraceptive implant
C0375850|ICD9CM|AB|V45.52|Prsc sbdrml cntrcp mplnt
C0375851|ICD9CM|PT|V45.59|Presence of other contraceptive device
C0375851|ICD9CM|AB|V45.59|Prsc other cntrcptv dvc
C0375852|ICD9CM|PT|V45.82|Percutaneous transluminal coronary angioplasty status
C0375852|ICD9CM|AB|V45.82|Status-post ptca
C0375853|ICD9CM|PT|V45.83|Breast implant removal status
C0375853|ICD9CM|AB|V45.83|Breast impl remov status
C0375854|ICD9CM|PT|V49.62|Other finger(s) amputation status
C0375854|ICD9CM|AB|V49.62|Status amput oth fingers
C0375855|ICD9CM|HT|V50.4|Prophylactic organ removal
C0375859|ICD9CM|HT|V52|Fitting and adjustment of prosthetic device and implant
C0375860|ICD9CM|PT|V52.4|Fitting and adjustment of breast prosthesis and implant
C0375860|ICD9CM|AB|V52.4|Fit/adj breast pros/impl
C0375861|ICD9CM|PT|V53.32|Fitting and adjustment of automatic implantable cardiac defibrillator
C0375861|ICD9CM|AB|V53.32|Ftng autmtc dfibrillator
C0375862|ICD9CM|PT|V53.39|Fitting and adjustment of other cardiac device
C0375862|ICD9CM|AB|V53.39|Ftng oth cardiac device
C0375864|ICD9CM|HT|V56|Encounter for dialysis and dialysis catheter care
C0375866|ICD9CM|PT|V57.22|Encounter for vocational therapy
C0375866|ICD9CM|AB|V57.22|Encntr vocational thrpy
C0375867|ICD9CM|PT|V58.41|Encounter for planned post-operative wound closure
C0375867|ICD9CM|AB|V58.41|Encntr plnd po wnd clsr
C0375868|ICD9CM|PT|V58.49|Other specified aftercare following surgery
C0375868|ICD9CM|AB|V58.49|Postop oth specfd aftrcr
C0375869|ICD9CM|HT|V58.6|Encounter for long-term (current) drug use
C0375871|ICD9CM|PT|V58.69|Long-term (current) use of other medications
C0375871|ICD9CM|AB|V58.69|Long-term use meds NEC
C0375872|ICD9CM|HT|V58.8|Encounter for other specified procedures and aftercare
C0375873|ICD9CM|PT|V58.81|Fitting and adjustment of vascular catheter
C0375873|ICD9CM|AB|V58.81|Fit/adj vascular cathetr
C0375874|ICD9CM|PT|V58.82|Fitting and adjustment of nonvascular catheter, NEC
C0375874|ICD9CM|AB|V58.82|Fit/adj non-vsc cath NEC
C0375878|ICD9CM|PT|V59.09|Other blood donors
C0375878|ICD9CM|AB|V59.09|Blood donor NEC
C0375879|ICD9CM|HT|V61.1|Counseling for marital and partner problems
C0375880|ICD9CM|PT|V61.10|Counseling for marital and partner problems, unspecified
C0375880|ICD9CM|AB|V61.10|Consl partner prob
C0375882|ICD9CM|PT|V61.20|Counseling for parent-child problem, unspecified
C0375882|ICD9CM|AB|V61.20|Cnsl prnt-chld prob NOS
C0375883|ICD9CM|PT|V61.21|Counseling for victim of child abuse
C0375883|ICD9CM|AB|V61.21|Cnsl victim child abuse
C0375885|ICD9CM|PT|V62.83|Counseling for perpetrator of physical/sexual abuse
C0375885|ICD9CM|AB|V62.83|Cnsl perp phys/sex abuse
C0375886|ICD9CM|AB|V65.41|Exercise counseling
C0375886|ICD9CM|PT|V65.41|Exercise counseling
C0375888|ICD9CM|PT|V65.43|Counseling on injury prevention
C0375888|ICD9CM|AB|V65.43|Counseling injry prevent
C0375890|ICD9CM|PT|V65.45|Counseling on other sexually transmitted diseases
C0375890|ICD9CM|AB|V65.45|Consln ot sex trnsmt dis
C0375891|ICD9CM|HT|V66|Convalescence and palliative care
C0375892|ICD9CM|PT|V66.7|Encounter for palliative care
C0375892|ICD9CM|AB|V66.7|Encountr palliative care
C0375893|ICD9CM|HT|V71|Observation and evaluation for suspected conditions not found
C0375894|ICD9CM|PT|V72.81|Pre-operative cardiovascular examination
C0375894|ICD9CM|AB|V72.81|Preop cardiovsclr exam
C0375895|ICD9CM|PT|V72.82|Pre-operative respiratory examination
C0375895|ICD9CM|AB|V72.82|Preop respiratory exam
C0375896|ICD9CM|PT|V72.83|Other specified pre-operative examination
C0375896|ICD9CM|AB|V72.83|Oth spcf preop exam
C0375897|ICD9CM|PT|V72.84|Pre-operative examination, unspecified
C0375897|ICD9CM|AB|V72.84|Preop exam unspcf
C0375898|ICD9CM|HT|V73|Special screening examination for viral and chlamydial diseases
C0375899|ICD9CM|PT|V73.88|Special screening examination for other specified chlamydial diseases
C0375899|ICD9CM|AB|V73.88|Scrn oth spcf chlmyd dis
C0375900|ICD9CM|PT|V73.98|Special screening examination for unspecified chlamydial disease
C0375900|ICD9CM|AB|V73.98|Scrn unspcf chlmyd dis
C0375901|ICD9CM|PT|02.96|Insertion of sphenoidal electrodes
C0375901|ICD9CM|AB|02.96|Insert sphenoid electrod
C0375906|ICD9CM|PT|07.15|Biopsy of pituitary gland, unspecified approach
C0375906|ICD9CM|AB|07.15|Pituitary biopsy NOS
C0375917|ICD9CM|PT|13.65|Excision of secondary membrane [after cataract]
C0375917|ICD9CM|AB|13.65|After-cataract excision
C0375921|ICD9CM|PT|16.93|Excision of lesion of eye, unspecified structure
C0375921|ICD9CM|AB|16.93|Excision eye lesion NOS
C0375926|ICD9CM|PT|22.50|Sinusotomy, not otherwise specified
C0375926|ICD9CM|AB|22.50|Sinusotomy NOS
C0375934|ICD9CM|PT|34.05|Creation of pleuroperitoneal shunt
C0375934|ICD9CM|AB|34.05|PlEuroperitoneal shunt
C0375941|ICD9CM|PT|36.17|Abdominal-coronary artery bypass
C0375941|ICD9CM|AB|36.17|Abd-coron artery bypass
C0375945|ICD9CM|PT|37.70|Initial insertion of lead [electrode], not otherwise specified
C0375945|ICD9CM|AB|37.70|Int insert pacemak lead
C0375946|ICD9CM|PT|37.76|Replacement of transvenous atrial and/or ventricular lead(s) [electrode]
C0375946|ICD9CM|AB|37.76|Repl tv atri-vent lead
C0375949|ICD9CM|PT|38.10|Endarterectomy, unspecified site
C0375949|ICD9CM|AB|38.10|Endarterectomy NOS
C0375951|ICD9CM|PT|38.40|Resection of vessel with replacement, unspecified site
C0375951|ICD9CM|AB|38.40|Vessel resect/replac NOS
C0375952|ICD9CM|PT|38.50|Ligation and stripping of varicose veins, unspecified site
C0375952|ICD9CM|AB|38.50|Varicose v lig-strip NOS
C0375953|ICD9CM|PT|38.60|Other excision of vessels, unspecified site
C0375953|ICD9CM|AB|38.60|Excision of vessel NOS
C0375954|ICD9CM|PT|38.80|Other surgical occlusion of vessels, unspecified site
C0375954|ICD9CM|AB|38.80|Surg vessel occlus NEC
C0375956|ICD9CM|HT|39.6|Extracorporeal circulation and procedures auxiliary to heart surgery
C0375961|ICD9CM|HT|41.0|Bone marrow or hematopoietic stem cell transplant
C0375969|ICD9CM|PT|45.27|Intestinal biopsy, site unspecified
C0375969|ICD9CM|AB|45.27|Intestinal biopsy NOS
C0375970|ICD9CM|PT|45.29|Other diagnostic procedures on intestine, site unspecified
C0375970|ICD9CM|AB|45.29|Bowel diagnost proc NEC
C0375971|ICD9CM|PT|45.43|Endoscopic destruction of other lesion or tissue of large intestine
C0375971|ICD9CM|AB|45.43|Endosc destru lg int les
C0375972|ICD9CM|HT|45.5|Isolation of intestinal segment
C0375972|ICD9CM|PT|45.50|Isolation of intestinal segment, not otherwise specified
C0375972|ICD9CM|AB|45.50|Intest seg isolat NOS
C0375979|ICD9CM|PT|47.11|Laparoscopic incidental appendectomy
C0375979|ICD9CM|AB|47.11|Lap incid appendectomy
C0375980|ICD9CM|PT|47.19|Other incidental appendectomy
C0375980|ICD9CM|AB|47.19|Other incid appendectomy
C0375981|ICD9CM|PT|48.36|[Endoscopic] polypectomy of rectum
C0375981|ICD9CM|AB|48.36|Polypectomy of rectum
C0375982|ICD9CM|PT|51.21|Other partial cholecystectomy
C0375982|ICD9CM|AB|51.21|Oth part cholecystectomy
C0375983|ICD9CM|PT|51.24|Laparoscopic partial cholecystectomy
C0375983|ICD9CM|AB|51.24|Lap part cholecystectomy
C0375984|ICD9CM|PT|51.51|Exploration of common duct
C0375984|ICD9CM|AB|51.51|Common duct exploration
C0375985|ICD9CM|PT|51.59|Other incision of other bile duct
C0375985|ICD9CM|AB|51.59|Bile duct incision NEC
C0375987|ICD9CM|PT|52.84|Autotransplantation of cells of Islets of Langerhans
C0375987|ICD9CM|AB|52.84|Autotrnsplnt islets lang
C0375988|ICD9CM|PT|52.85|Allotransplantation of cells of Islets of Langerhans
C0375988|ICD9CM|AB|52.85|Allotrnsplnt islets lang
C0375989|ICD9CM|PT|52.86|Transplantation of cells of Islets of Langerhans, not otherwise specified
C0375989|ICD9CM|AB|52.86|Trnsplnt islets lang NOS
C0375996|ICD9CM|PT|54.59|Other lysis of peritoneal adhesions
C0375996|ICD9CM|AB|54.59|Oth periton adhesiolysis
C0376001|ICD9CM|PT|59.03|Laparoscopic lysis of perirenal or periureteral adhesions
C0376001|ICD9CM|AB|59.03|Lap lys periren/uret adh
C0376002|ICD9CM|PT|59.11|Other lysis of perivesical adhesions
C0376002|ICD9CM|AB|59.11|Oth lys perives adhesio
C0376003|ICD9CM|PT|59.72|Injection of implant into urethra and/or bladder neck
C0376003|ICD9CM|AB|59.72|Inject implant urethra
C0376004|ICD9CM|PT|60.21|Transurethral (ultrasound) guided laser induced prostatectomy (TULIP)
C0376004|ICD9CM|AB|60.21|Transureth prostatectomy
C0376005|ICD9CM|PT|60.29|Other transurethral prostatectomy
C0376005|ICD9CM|AB|60.29|Oth transureth prostatec
C0376007|ICD9CM|AB|65.01|Laparoscopic oophorotomy
C0376007|ICD9CM|PT|65.01|Laparoscopic oophorotomy
C0376008|ICD9CM|AB|65.09|Other oophorotomy
C0376008|ICD9CM|PT|65.09|Other oophorotomy
C0376009|ICD9CM|PT|65.14|Other laparoscopic diagnostic procedures on ovaries
C0376009|ICD9CM|AB|65.14|Oth lap dx proc ovaries
C0376011|ICD9CM|PT|65.24|Laparoscopic wedge resection of ovary
C0376011|ICD9CM|AB|65.24|Lap wedge resect ovary
C0376012|ICD9CM|PT|65.25|Other laparoscopic local excision or destruction of ovary
C0376012|ICD9CM|AB|65.25|Oth lap loc exc dest ova
C0376013|ICD9CM|PT|65.31|Laparoscopic unilateral oophorectomy
C0376013|ICD9CM|AB|65.31|Lap unilat oophorectomy
C0376014|ICD9CM|PT|65.39|Other unilateral oophorectomy
C0376014|ICD9CM|AB|65.39|Oth unilat oophorectomy
C0376015|ICD9CM|PT|65.41|Laparoscopic unilateral salpingo-oophorectomy
C0376015|ICD9CM|AB|65.41|Lap uni salpingo-oophor
C0376016|ICD9CM|PT|65.49|Other unilateral salpingo-oophorectomy
C0376016|ICD9CM|AB|65.49|Oth uni salpingo-oophor
C0376018|ICD9CM|PT|65.52|Other removal of remaining ovary
C0376018|ICD9CM|AB|65.52|Oth remove remain ovary
C0376019|ICD9CM|PT|65.53|Laparoscopic removal of both ovaries at same operative episode
C0376019|ICD9CM|AB|65.53|Lap remove both ovaries
C0376020|ICD9CM|PT|65.54|Laparoscopic removal of remaining ovary
C0376020|ICD9CM|AB|65.54|Lap remove remain ovary
C0376021|ICD9CM|PT|65.61|Other removal of both ovaries and tubes at same operative episode
C0376021|ICD9CM|AB|65.61|Oth remove ovaries/tubes
C0376022|ICD9CM|PT|65.62|Other removal of remaining ovary and tube
C0376022|ICD9CM|AB|65.62|Oth remove rem ova/tube
C0376023|ICD9CM|PT|65.63|Laparoscopic removal of both ovaries and tubes at same operative episode
C0376023|ICD9CM|AB|65.63|Lap remove ovaries/tubes
C0376024|ICD9CM|PT|65.64|Laparoscopic removal of remaining ovary and tube
C0376024|ICD9CM|AB|65.64|Lap remove rem ova/tube
C0376025|ICD9CM|PT|65.71|Other simple suture of ovary
C0376025|ICD9CM|AB|65.71|Oth simple suture ovary
C0376026|ICD9CM|PT|65.72|Other reimplantation of ovary
C0376026|ICD9CM|AB|65.72|Oth reimplant of ovary
C0376027|ICD9CM|PT|65.73|Other salpingo-oophoroplasty
C0376027|ICD9CM|AB|65.73|Oth salpingo-oophoroplas
C0376028|ICD9CM|PT|65.74|Laparoscopic simple suture of ovary
C0376028|ICD9CM|AB|65.74|Lap simple suture ovary
C0376029|ICD9CM|PT|65.75|Laparoscopic reimplantation of ovary
C0376029|ICD9CM|AB|65.75|Lap reimplant of ovary
C0376030|ICD9CM|PT|65.76|Laparoscopic salpingo-oophoroplasty
C0376030|ICD9CM|AB|65.76|Lap salpingo-oophoroplas
C0376031|ICD9CM|PT|65.81|Laparoscopic lysis of adhesions of ovary and fallopian tube
C0376031|ICD9CM|AB|65.81|Lap adhesiolys ova/tube
C0376032|ICD9CM|PT|65.89|Other lysis of adhesions of ovary and fallopian tube
C0376032|ICD9CM|AB|65.89|Adhesiolysis ovary/tube
C0376037|ICD9CM|PT|68.9|Other and unspecified hysterectomy
C0376037|ICD9CM|AB|68.9|Hysterectomy NEC/NOS
C0376038|ICD9CM|PT|69.09|Other dilation and curettage
C0376038|ICD9CM|AB|69.09|D & C NEC
C0376039|ICD9CM|PT|69.21|Interposition operation
C0376039|ICD9CM|AB|69.21|Interposit op uterin lig
C0376040|ICD9CM|PT|74.3|Removal of extratubal ectopic pregnancy
C0376040|ICD9CM|AB|74.3|Rem extratub ectop preg
C0376044|ICD9CM|PT|77.10|Other incision of bone without division, unspecified site
C0376044|ICD9CM|AB|77.10|Other bone incision NOS
C0376047|ICD9CM|PT|77.60|Local excision of lesion or tissue of bone, unspecified site
C0376047|ICD9CM|AB|77.60|Loc exc bone lesion NOS
C0376048|ICD9CM|PT|77.70|Excision of bone for graft, unspecified site
C0376048|ICD9CM|AB|77.70|Excise bone for grft NOS
C0376049|ICD9CM|PT|77.80|Other partial ostectomy, unspecified site
C0376049|ICD9CM|HT|77.8|Other partial ostectomy
C0376049|ICD9CM|AB|77.80|Oth part ostectomy NOS
C0376050|ICD9CM|PT|77.90|Total ostectomy, unspecified site
C0376050|ICD9CM|AB|77.90|Total ostectomy NOS
C0376052|ICD9CM|PT|78.10|Application of external fixator device, unspecified site
C0376052|ICD9CM|AB|78.10|Applic ext fix dev NOS
C0376053|ICD9CM|PT|78.20|Limb shortening procedures, unspecified site
C0376053|ICD9CM|AB|78.20|Limb shorten proc NOS
C0376055|ICD9CM|PT|78.40|Other repair or plastic operations on bone, unspecified site
C0376055|ICD9CM|HT|78.4|Other repair or plastic operations on bone
C0376055|ICD9CM|AB|78.40|Oth bone repair/plast op
C0376056|ICD9CM|PT|78.50|Internal fixation of bone without fracture reduction, unspecified site
C0376056|ICD9CM|AB|78.50|Int fix w/o fx reduc NOS
C0376057|ICD9CM|PT|78.60|Removal of implanted devices from bone, unspecified site
C0376057|ICD9CM|AB|78.60|Remove imp device NOS
C0376059|ICD9CM|PT|78.80|Diagnostic procedures on bone, not elsewhere classified, unspecified site
C0376059|ICD9CM|HT|78.8|Diagnostic procedures on bone, not elsewhere classified
C0376059|ICD9CM|AB|78.80|Other bone dx proc NOS
C0376063|ICD9CM|PT|79.20|Open reduction of fracture without internal fixation, unspecified site
C0376063|ICD9CM|AB|79.20|Open fx reduction NOS
C0376064|ICD9CM|PT|79.30|Open reduction of fracture with internal fixation, unspecified site
C0376064|ICD9CM|AB|79.30|Opn fx red w int fix NOS
C0376065|ICD9CM|PT|79.40|Closed reduction of separated epiphysis, unspecified site
C0376065|ICD9CM|AB|79.40|Cls reduc-sep epiphy NOS
C0376066|ICD9CM|PT|79.50|Open reduction of separated epiphysis, unspecified site
C0376066|ICD9CM|AB|79.50|Open red-sep epiphy NOS
C0376067|ICD9CM|PT|79.90|Unspecified operation on bone injury, unspecified site
C0376067|ICD9CM|AB|79.90|Unspec op bone inj NOS
C0376069|ICD9CM|PT|80.10|Other arthrotomy, unspecified site
C0376069|ICD9CM|AB|80.10|Other arthrotomy NOS
C0376070|ICD9CM|PT|80.20|Arthroscopy, unspecified site
C0376070|ICD9CM|AB|80.20|Arthroscopy NOS
C0376071|ICD9CM|AB|80.30|Joint biopsy NOS
C0376071|ICD9CM|PT|80.30|Biopsy of joint structure, unspecified site
C0376072|ICD9CM|PT|80.40|Division of joint capsule, ligament, or cartilage, unspecified site
C0376072|ICD9CM|AB|80.40|Jt structur division NOS
C0376073|ICD9CM|PT|80.50|Excision or destruction of intervertebral disc, unspecified
C0376073|ICD9CM|AB|80.50|Exc/dest intvrt disc NOS
C0376075|ICD9CM|PT|80.80|Other local excision or destruction of lesion of joint, unspecified site
C0376075|ICD9CM|AB|80.80|Destruct joint les NOS
C0376076|ICD9CM|PT|80.90|Other excision of joint, unspecified site
C0376076|ICD9CM|AB|80.90|Excision of joint NOS
C0376078|ICD9CM|PT|81.59|Revision of joint replacement of lower extremity, not elsewhere classified
C0376078|ICD9CM|AB|81.59|Rev jt repl low ext NEC
C0376079|ICD9CM|PT|81.97|Revision of joint replacement of upper extremity
C0376079|ICD9CM|AB|81.97|Rev jt repl upper extrem
C0376083|ICD9CM|PT|85.20|Excision or destruction of breast tissue, not otherwise specified
C0376083|ICD9CM|HT|85.2|Excision or destruction of breast tissue
C0376083|ICD9CM|AB|85.20|Breast tissu destruc NOS
C0376086|ICD9CM|PT|86.70|Pedicle or flap graft, not otherwise specified
C0376086|ICD9CM|HT|86.7|Pedicle grafts or flaps
C0376086|ICD9CM|AB|86.70|Pedicle graft/flap NOS
C0376089|ICD9CM|PT|88.40|Arteriography using contrast material, unspecified site
C0376089|ICD9CM|AB|88.40|Contrast arteriogram NOS
C0376091|ICD9CM|PT|88.60|Phlebography using contrast material, unspecified site
C0376091|ICD9CM|AB|88.60|Contrast phlebogram NOS
C0376094|ICD9CM|PT|89.10|Intracarotid amobarbital test
C0376094|ICD9CM|AB|89.10|Intracarot amobarb test
C0376100|ICD9CM|PT|98.59|Extracorporeal shockwave lithotripsy of other sites
C0376100|ICD9CM|AB|98.59|Eswl other sites
C0376101|ICD9CM|PT|99.00|Perioperative autologous transfusion of whole blood or blood components
C0376101|ICD9CM|AB|99.00|Periop aut trans hol bld
C0376102|ICD9CM|PT|99.02|Transfusion of previously collected autologous blood
C0376102|ICD9CM|AB|99.02|Transfus prev auto blood
C0376103|ICD9CM|PT|99.28|Injection or infusion of biological response modifier [BRM] as an antineoplastic agent
C0376103|ICD9CM|AB|99.28|Immunotherapy as antineo
C0376105|ICD9CM|PT|99.79|Other therapeutic apheresis
C0376105|ICD9CM|AB|99.79|Other therapeu apheresis
C0376106|ICD9CM|HT|860-869.99|INTERNAL INJURY OF THORAX, ABDOMEN, AND PELVIS
C0376108|ICD9CM|HT|V07-V09.99|PERSONS WITH NEED FOR ISOLATION, OTHER POTENTIAL HEALTH HAZARDS AND PROPHYLACTIC MEASURES
C0376109|ICD9CM|HT|E000-E999.9|SUPPLEMENTARY CLASSIFICATION OF EXTERNAL CAUSES OF INJURY AND POISONING
C0376110|ICD9CM|PT|077.98|Unspecified diseases of conjunctiva due to chlamydiae
C0376110|ICD9CM|AB|077.98|Unsp ds conjuc chlamydia
C0376111|ICD9CM|PT|077.99|Unspecified diseases of conjunctiva due to viruses
C0376111|ICD9CM|AB|077.99|Unsp ds conjuc viruses
C0376115|ICD9CM|PT|429.71|Acquired cardiac septal defect
C0376115|ICD9CM|AB|429.71|Acq cardiac septl defect
C0376117|ICD9CM|PT|702.11|Inflamed seborrheic keratosis
C0376117|ICD9CM|AB|702.11|Inflamed sbrheic keratos
C0376124|ICD9CM|PT|V49.75|Below knee amputation status
C0376124|ICD9CM|AB|V49.75|Status amput below knee
C0376125|ICD9CM|PT|V49.76|Above knee amputation status
C0376125|ICD9CM|AB|V49.76|Status amput above knee
C0376128|ICD9CM|PT|250.52|Diabetes with ophthalmic manifestations, type II or unspecified type, uncontrolled
C0376128|ICD9CM|AB|250.52|DMII ophth uncntrld
C0376129|ICD9CM|PT|344.01|Quadriplegia, C1-C4, complete
C0376129|ICD9CM|AB|344.01|Quadrplg c1-c4, complete
C0376130|ICD9CM|PT|344.02|Quadriplegia, C1-C4, incomplete
C0376130|ICD9CM|AB|344.02|Quadrplg c1-c4, incomplt
C0376131|ICD9CM|PT|344.03|Quadriplegia, C5-C7, complete
C0376131|ICD9CM|AB|344.03|Quadrplg c5-c7, complete
C0376132|ICD9CM|PT|344.04|Quadriplegia, C5-C7, incomplete
C0376132|ICD9CM|AB|344.04|Quadrplg c5-c7, incomplt
C0376137|ICD9CM|HT|V49.6|Status post amputation of upper limb
C0376138|ICD9CM|PT|V49.60|Unspecified level upper limb amputation status
C0376138|ICD9CM|AB|V49.60|Status amput up lmb NOS
C0376139|ICD9CM|PT|V49.61|Thumb amputation status
C0376139|ICD9CM|AB|V49.61|Status amput thumb
C0376140|ICD9CM|PT|V49.63|Hand amputation status
C0376140|ICD9CM|AB|V49.63|Status amput hand
C0376141|ICD9CM|PT|V49.64|Wrist amputation status
C0376141|ICD9CM|AB|V49.64|Status amput wrist
C0376142|ICD9CM|PT|V49.65|Below elbow amputation status
C0376142|ICD9CM|AB|V49.65|Status amput below elbow
C0376143|ICD9CM|PT|V49.66|Above elbow amputation status
C0376143|ICD9CM|AB|V49.66|Status amput above elbow
C0376144|ICD9CM|PT|V49.67|Shoulder amputation status
C0376144|ICD9CM|AB|V49.67|Status amput shoulder
C0376175|ICD9CM|AB|351.0|Bell's palsy
C0376175|ICD9CM|PT|351.0|Bell's palsy
C0376329|ICD9CM|PT|046.11|Variant Creutzfeldt-Jakob disease
C0376329|ICD9CM|AB|046.11|Varnt Creutzfeldt-Jakob
C0376356|ICD9CM|AB|625.4|Premenstrual tension
C0376356|ICD9CM|PT|625.4|Premenstrual tension syndromes
C0376358|ICD9CM|PT|185|Malignant neoplasm of prostate
C0376358|ICD9CM|AB|185|Malign neopl prostate
C0376379|ICD9CM|PT|054.2|Herpetic gingivostomatitis
C0376379|ICD9CM|AB|054.2|Herpetic gingivostomat
C0376620|ICD9CM|AB|569.71|Pouchitis
C0376620|ICD9CM|PT|569.71|Pouchitis
C0391820|ICD9CM|HT|274.1|Gouty nephropathy
C0391820|ICD9CM|AB|274.10|Gouty nephropathy NOS
C0391820|ICD9CM|PT|274.10|Gouty nephropathy, unspecified
C0391870|ICD9CM|HT|790.0|Abnormality of red blood cells
C0391983|ICD9CM|HT|532.5|Chronic or unspecified duodenal ulcer with perforation
C0391984|ICD9CM|HT|532.9|Duodenal ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation
C0391994|ICD9CM|AB|V45.4|Arthrodesis status
C0391994|ICD9CM|PT|V45.4|Arthrodesis status
C0392044|ICD9CM|PT|901.81|Injury to intercostal artery or vein
C0392044|ICD9CM|AB|901.81|Inj intercostal art/vein
C0392054|ICD9CM|PT|031.0|Pulmonary diseases due to other mycobacteria
C0392054|ICD9CM|AB|031.0|Pulmonary mycobacteria
C0392098|ICD9CM|PT|V42.6|Lung replaced by transplant
C0392098|ICD9CM|AB|V42.6|Lung transplant status
C0392099|ICD9CM|PT|V42.3|Skin replaced by transplant
C0392099|ICD9CM|AB|V42.3|Skin transplant status
C0392440|ICD9CM|PT|701.2|Acquired acanthosis nigricans
C0392440|ICD9CM|AB|701.2|Acq acanthosis nigricans
C0392470|ICD9CM|PT|426.7|Anomalous atrioventricular excitation
C0392470|ICD9CM|AB|426.7|Anomalous av excitation
C0392477|ICD9CM|AB|754.61|Congenital pes planus
C0392477|ICD9CM|PT|754.61|Congenital pes planus
C0392485|ICD9CM|AB|750.27|Diverticulum of pharynx
C0392485|ICD9CM|PT|750.27|Diverticulum of pharynx
C0392492|ICD9CM|PT|522.6|Chronic apical periodontitis
C0392492|ICD9CM|AB|522.6|Chr apical periodontitis
C0392494|ICD9CM|PT|529.3|Hypertrophy of tongue papillae
C0392494|ICD9CM|AB|529.3|Hypertroph tongue papill
C0392499|ICD9CM|HT|533.3|Acute peptic ulcer of unspecified site without mention of hemorrhage and perforation
C0392501|ICD9CM|HT|534.3|Acute gastrojejunal ulcer without mention of hemorrhage or perforation
C0392502|ICD9CM|HT|534.7|Chronic gastrojejunal ulcer without mention of hemorrhage or perforation
C0392503|ICD9CM|HT|560.3|Impaction of intestine
C0392503|ICD9CM|AB|560.30|Impaction intestine NOS
C0392503|ICD9CM|PT|560.30|Impaction of intestine, unspecified
C0392514|ICD9CM|PT|275.01|Hereditary hemochromatosis
C0392514|ICD9CM|AB|275.01|Heredit hemochromatosis
C0392530|ICD9CM|PT|618.3|Uterovaginal prolapse, complete
C0392530|ICD9CM|AB|618.3|Uterovag prolaps-complet
C0392531|ICD9CM|AB|608.23|Torsion appendix testis
C0392531|ICD9CM|PT|608.23|Torsion of appendix testis
C0392536|ICD9CM|HT|638|Failed attempted abortion
C0392548|ICD9CM|HT|344.6|Cauda equina syndrome
C0392549|ICD9CM|HT|343|Infantile cerebral palsy
C0392549|ICD9CM|AB|343.9|Cerebral palsy NOS
C0392549|ICD9CM|PT|343.9|Infantile cerebral palsy, unspecified
C0392550|ICD9CM|AB|343.4|Infantile hemiplegia
C0392550|ICD9CM|PT|343.4|Infantile hemiplegia
C0392553|ICD9CM|PT|356.0|Hereditary peripheral neuropathy
C0392553|ICD9CM|AB|356.0|Hered periph neuropathy
C0392558|ICD9CM|PT|369.03|Better eye: near-total vision impairment; lesser eye: total vision impairment
C0392558|ICD9CM|AB|369.03|One eye-near tot/oth-tot
C0392559|ICD9CM|PT|369.05|Better eye: profound vision impairment; lesser eye: not further specified
C0392559|ICD9CM|AB|369.05|One eye-profound/oth-NOS
C0392560|ICD9CM|PT|369.06|Better eye: profound vision impairment; lesser eye: total vision impairment
C0392560|ICD9CM|AB|369.06|One eye-profound/oth-tot
C0392561|ICD9CM|PT|369.07|Better eye: profound vision impairment; lesser eye: near-total vision impairment
C0392561|ICD9CM|AB|369.07|One eye-prfnd/oth-nr tot
C0392562|ICD9CM|PT|369.11|Better eye: severe vision impairment; lesser eye: blind, not further specified
C0392562|ICD9CM|AB|369.11|1 eye-sev/oth-blind NOS
C0392563|ICD9CM|PT|369.12|Better eye: severe vision impairment; lesser eye: total vision impairment
C0392563|ICD9CM|AB|369.12|One eye-severe/oth-total
C0392564|ICD9CM|PT|369.13|Better eye: severe vision impairment; lesser eye: near-total vision impairment
C0392564|ICD9CM|AB|369.13|One eye-sev/oth-near tot
C0392565|ICD9CM|PT|369.14|Better eye: severe vision impairment; lesser eye: profound vision impairment
C0392565|ICD9CM|AB|369.14|One eye-sev/oth-prfnd
C0392566|ICD9CM|PT|369.15|Better eye: moderate vision impairment; lesser eye: blind, not further specified
C0392566|ICD9CM|AB|369.15|One eye-mod/oth-blind
C0392567|ICD9CM|PT|369.16|Better eye: moderate vision impairment; lesser eye: total vision impairment
C0392567|ICD9CM|AB|369.16|One eye-moderate/oth-tot
C0392568|ICD9CM|PT|369.17|Better eye: moderate vision impairment; lesser eye: near-total vision impairment
C0392568|ICD9CM|AB|369.17|One eye-mod/oth-near tot
C0392569|ICD9CM|PT|369.18|Better eye: moderate vision impairment; lesser eye: profound vision impairment
C0392569|ICD9CM|AB|369.18|One eye-mod/oth-profound
C0392570|ICD9CM|PT|369.21|Better eye: severe vision impairment; lesser eye; impairment not further specified
C0392570|ICD9CM|AB|369.21|One eye-severe/oth-NOS
C0392571|ICD9CM|PT|369.23|Better eye: moderate vision impairment; lesser eye: impairment not further specified
C0392571|ICD9CM|AB|369.23|One eye-moderate/oth-NOS
C0392572|ICD9CM|PT|369.24|Better eye: moderate vision impairment; lesser eye: severe vision impairment
C0392572|ICD9CM|AB|369.24|One eye-moderate/oth-sev
C0392573|ICD9CM|PT|369.62|One eye: total vision impairment; other eye: near-normal vision
C0392573|ICD9CM|AB|369.62|One eye-tot/oth-near nor
C0392574|ICD9CM|PT|369.63|One eye: total vision impairment; other eye: normal vision
C0392574|ICD9CM|AB|369.63|One eye-total/oth-normal
C0392575|ICD9CM|PT|369.64|One eye: near-total vision impairment; other eye: vision not specified
C0392575|ICD9CM|AB|369.64|One eye-near tot/oth-NOS
C0392576|ICD9CM|PT|369.65|One eye: near-total vision impairment; other eye: near-normal vision
C0392576|ICD9CM|AB|369.65|Near-tot imp/near-normal
C0392577|ICD9CM|PT|369.66|One eye: near-total vision impairment; other eye: normal vision
C0392577|ICD9CM|AB|369.66|Near-total impair/normal
C0392578|ICD9CM|PT|369.67|One eye: profound vision impairment; other eye: vision not specified
C0392578|ICD9CM|AB|369.60|Blindness, one eye
C0392578|ICD9CM|PT|369.60|Profound impairment, one eye, impairment level not further specified
C0392578|ICD9CM|AB|369.67|One eye-prfound/oth-unkn
C0392579|ICD9CM|PT|369.68|One eye: profound vision impairment; other eye: near-normal vision
C0392579|ICD9CM|AB|369.68|Profnd impair/near norm
C0392580|ICD9CM|PT|369.69|One eye: profound vision impairment; other eye: normal vision
C0392580|ICD9CM|AB|369.69|Profound impair/normal
C0392581|ICD9CM|PT|369.71|One eye: severe vision impairment; other eye: vision not specified
C0392581|ICD9CM|AB|369.71|One eye-severe/oth-unknw
C0392582|ICD9CM|PT|369.72|One eye: severe vision impairment; other eye: near-normal vision
C0392582|ICD9CM|AB|369.72|One eye-sev/oth-nr norm
C0392583|ICD9CM|PT|369.73|One eye: severe vision impairment; other eye: normal vision
C0392583|ICD9CM|AB|369.73|One eye-severe/oth-norm
C0392584|ICD9CM|PT|369.74|One eye: moderate vision impairment; other eye: vision not specified
C0392584|ICD9CM|AB|369.74|One eye-mod/other-unknwn
C0392585|ICD9CM|PT|369.75|One eye: moderate vision impairment; other eye: near-normal vision
C0392585|ICD9CM|AB|369.75|One eye-mod/oth-nr norm
C0392586|ICD9CM|PT|369.76|One eye: moderate vision impairment; other eye: normal vision
C0392586|ICD9CM|AB|369.76|One eye-mod/oth normal
C0392587|ICD9CM|AB|374.31|Paralytic ptosis
C0392587|ICD9CM|PT|374.31|Paralytic ptosis
C0392611|ICD9CM|PT|824.4|Bimalleolar fracture, closed
C0392611|ICD9CM|AB|824.4|Fx bimalleolar-closed
C0392617|ICD9CM|PT|997.61|Neuroma of amputation stump
C0392617|ICD9CM|AB|997.61|Neuroma amputation stump
C0392618|ICD9CM|HT|998.5|Postoperative infection
C0392622|ICD9CM|PT|982.1|Toxic effect of carbon tetrachloride
C0392622|ICD9CM|AB|982.1|Toxic eff carbon tetrach
C0392646|ICD9CM|PT|054.9|Herpes simplex without mention of complication
C0392646|ICD9CM|AB|054.9|Herpes simplex NOS
C0392650|ICD9CM|PT|055.9|Measles without mention of complication
C0392650|ICD9CM|AB|055.9|Measles uncomplicated
C0392663|ICD9CM|AB|125.0|Bancroftian filariasis
C0392663|ICD9CM|PT|125.0|Bancroftian filariasis
C0392682|ICD9CM|PT|796.2|Elevated blood pressure reading without diagnosis of hypertension
C0392682|ICD9CM|AB|796.2|Elev bl pres w/o hypertn
C0392702|ICD9CM|PT|781.0|Abnormal involuntary movements
C0392702|ICD9CM|AB|781.0|Abn involun movement NEC
C0392799|ICD9CM|PT|97.88|Removal of external immobilization device
C0392799|ICD9CM|AB|97.88|Remov ext immobilization
C0392801|ICD9CM|AB|83.94|Aspiration of bursa
C0392801|ICD9CM|PT|83.94|Aspiration of bursa
C0392807|ICD9CM|PT|84.07|Amputation through humerus
C0392807|ICD9CM|AB|84.07|Amputation thru humerus
C0392808|ICD9CM|PT|79.01|Closed reduction of fracture without internal fixation, humerus
C0392808|ICD9CM|AB|79.01|Closed fx reduct humerus
C0392829|ICD9CM|PT|35.91|Interatrial transposition of venous return
C0392829|ICD9CM|AB|35.91|Interat ven retrn transp
C0392832|ICD9CM|PT|35.04|Closed heart valvotomy, tricuspid valve
C0392832|ICD9CM|AB|35.04|Closed tricusp valvotomy
C0392852|ICD9CM|PT|64.96|Removal of internal prosthesis of penis
C0392852|ICD9CM|AB|64.96|Remove int penile prosth
C0392875|ICD9CM|PT|12.51|Goniopuncture without goniotomy
C0392875|ICD9CM|AB|12.51|Goniopuncture
C0392892|ICD9CM|AB|94.31|Psychoanalysis
C0392892|ICD9CM|PT|94.31|Psychoanalysis
C0393517|ICD9CM|PT|334.4|Cerebellar ataxia in diseases classified elsewhere
C0393517|ICD9CM|AB|334.4|Cerebel atax in oth dis
C0393570|ICD9CM|PT|331.6|Corticobasal degeneration
C0393570|ICD9CM|AB|331.6|Corticobasal degneration
C0393596|ICD9CM|PT|333.72|Acute dystonia due to drugs
C0393596|ICD9CM|AB|333.72|Acute dystonia d/t drugs
C0393647|ICD9CM|PT|331.7|Cerebral degeneration in diseases classified elsewhere
C0393647|ICD9CM|AB|331.7|Cereb degen in oth dis
C0393737|ICD9CM|PT|339.11|Episodic tension type headache
C0393737|ICD9CM|AB|339.11|Episdic tension headache
C0393738|ICD9CM|PT|339.12|Chronic tension type headache
C0393738|ICD9CM|AB|339.12|Chronic tension headache
C0393739|ICD9CM|PT|339.01|Episodic cluster headache
C0393739|ICD9CM|AB|339.01|Episodc cluster headache
C0393743|ICD9CM|PT|339.04|Chronic paroxysmal hemicrania
C0393743|ICD9CM|AB|339.04|Chr paroxysml hemicrania
C0393745|ICD9CM|PT|339.22|Chronic post-traumatic headache
C0393745|ICD9CM|AB|339.22|Chr post-trauma headache
C0393754|ICD9CM|PT|339.82|Headache associated with sexual activity
C0393754|ICD9CM|AB|339.82|Headache w sex activity
C0393770|ICD9CM|PT|327.31|Circadian rhythm sleep disorder, delayed sleep phase type
C0393770|ICD9CM|AB|327.31|Circadian rhy-delay slp
C0393772|ICD9CM|PT|327.34|Circadian rhythm sleep disorder, free-running type
C0393772|ICD9CM|AB|327.34|Circadian rhym-free run
C0393773|ICD9CM|PT|327.36|Circadian rhythm sleep disorder, shift work type
C0393773|ICD9CM|AB|327.36|Circadian rhy-shift work
C0393774|ICD9CM|AB|327.53|Sleep related bruxism
C0393774|ICD9CM|PT|327.53|Sleep related bruxism
C0393797|ICD9CM|PT|352.2|Other disorders of glossopharyngeal [9th] nerve
C0393797|ICD9CM|AB|352.2|Glossophar nerve dis NEC
C0393819|ICD9CM|PT|357.81|Chronic inflammatory demyelinating polyneuritis
C0393819|ICD9CM|AB|357.81|Chr inflam polyneuritis
C0393851|ICD9CM|PT|357.82|Critical illness polyneuropathy
C0393851|ICD9CM|AB|357.82|Crit illness neuropathy
C0393939|ICD9CM|PT|358.2|Toxic myoneural disorders
C0393939|ICD9CM|AB|358.2|Toxic myoneural disorder
C0394082|ICD9CM|HT|02.1|Repair of cerebral meninges
C0394158|ICD9CM|PT|02.93|Implantation or replacement of intracranial neurostimulator lead(s)
C0394158|ICD9CM|AB|02.93|Imp/repl brain stim lead
C0394208|ICD9CM|PT|02.42|Replacement of ventricular shunt
C0394208|ICD9CM|AB|02.42|Replace ventricle shunt
C0394374|ICD9CM|HT|44.0|Vagotomy
C0394374|ICD9CM|AB|44.00|Vagotomy NOS
C0394374|ICD9CM|PT|44.00|Vagotomy, not otherwise specified
C0394407|ICD9CM|PT|04.71|Hypoglossal-facial anastomosis
C0394407|ICD9CM|AB|04.71|Hypogloss-facial anastom
C0394646|ICD9CM|AB|94.24|Chemical shock therapy
C0394646|ICD9CM|PT|94.24|Chemical shock therapy
C0394932|ICD9CM|PT|05.32|Injection of neurolytic agent into sympathetic nerve
C0394932|ICD9CM|AB|05.32|Neurolyt injec-symp nrv
C0394996|ICD9CM|HT|303.0|Acute alcoholic intoxication
C0395020|ICD9CM|HT|08-16.99|OPERATIONS ON THE EYE
C0395087|ICD9CM|PT|16.31|Removal of ocular contents with synchronous implant into scleral shell
C0395087|ICD9CM|AB|16.31|Eye evisc w synch implan
C0395105|ICD9CM|PT|97.31|Removal of eye prosthesis
C0395105|ICD9CM|AB|97.31|Remove eye prosthesis
C0395166|ICD9CM|PT|08.24|Excision of major lesion of eyelid, full-thickness
C0395166|ICD9CM|AB|08.24|Exc maj les lid ful-thic
C0395208|ICD9CM|PT|08.02|Severing of blepharorrhaphy
C0395208|ICD9CM|AB|08.02|Blepharorrhaphy severing
C0395408|ICD9CM|PT|11.32|Excision of pterygium with corneal graft
C0395408|ICD9CM|AB|11.32|Pteryg exc w cornea grft
C0395450|ICD9CM|PT|12.87|Scleral reinforcement with graft
C0395450|ICD9CM|AB|12.87|Graft reinforce sclera
C0395490|ICD9CM|AB|12.73|Cyclophotocoagulation
C0395490|ICD9CM|PT|12.73|Cyclophotocoagulation
C0395536|ICD9CM|PT|13.8|Removal of implanted lens
C0395536|ICD9CM|AB|13.8|Implanted lens removal
C0395542|ICD9CM|HT|14.7|Operations on vitreous
C0395549|ICD9CM|PT|14.75|Injection of vitreous substitute
C0395549|ICD9CM|AB|14.75|Vitreous substitut injec
C0395567|ICD9CM|PT|14.55|Repair of retinal detachment with photocoagulation of unspecified type
C0395567|ICD9CM|AB|14.55|Detach ret photocoag NOS
C0395569|ICD9CM|PT|14.54|Repair of retinal detachment with laser photocoagulation
C0395569|ICD9CM|AB|14.54|Detach retina laser coag
C0395570|ICD9CM|PT|14.53|Repair of retinal detachment with xenon arc photocoagulation
C0395570|ICD9CM|AB|14.53|Detach retina xenon coag
C0395659|ICD9CM|PT|18.72|Reattachment of amputated ear
C0395659|ICD9CM|AB|18.72|Reattach amputated ear
C0395663|ICD9CM|PT|18.6|Reconstruction of external auditory canal
C0395663|ICD9CM|AB|18.6|Ext audit canal reconstr
C0395769|ICD9CM|PT|20.8|Operations on eustachian tube
C0395769|ICD9CM|AB|20.8|Eustachian tube ops
C0395839|ICD9CM|PT|380.51|Acquired stenosis of external ear canal secondary to trauma
C0395839|ICD9CM|AB|380.51|Stenosis ear d/t trauma
C0395841|ICD9CM|PT|380.52|Acquired stenosis of external ear canal secondary to surgery
C0395841|ICD9CM|AB|380.52|Stenosis ear d/t surgery
C0395842|ICD9CM|PT|380.53|Acquired stenosis of external ear canal secondary to inflammation
C0395842|ICD9CM|AB|380.53|Stenosis ear d/t inflam
C0395849|ICD9CM|PT|384.1|Chronic myringitis without mention of otitis media
C0395849|ICD9CM|AB|384.1|Chronic myringitis
C0395861|ICD9CM|PT|382.00|Acute suppurative otitis media without spontaneous rupture of eardrum
C0395861|ICD9CM|AB|382.00|Ac supp otitis media NOS
C0395862|ICD9CM|PT|382.01|Acute suppurative otitis media with spontaneous rupture of eardrum
C0395862|ICD9CM|AB|382.01|Ac supp OM w drum rupt
C0395863|ICD9CM|PT|381.02|Acute mucoid otitis media
C0395863|ICD9CM|AB|381.02|Ac mucoid otitis media
C0395865|ICD9CM|PT|381.03|Acute sanguinous otitis media
C0395865|ICD9CM|AB|381.03|Ac sanguin otitis media
C0395887|ICD9CM|HT|385.0|Tympanosclerosis
C0395887|ICD9CM|AB|385.00|Tympanosclerosis NOS
C0395887|ICD9CM|PT|385.00|Tympanosclerosis, unspecified as to involvement
C0395888|ICD9CM|PT|385.01|Tympanosclerosis involving tympanic membrane only
C0395888|ICD9CM|AB|385.01|Tympanoscl-tympanic memb
C0395889|ICD9CM|PT|385.02|Tympanosclerosis involving tympanic membrane and ear ossicles
C0395889|ICD9CM|AB|385.02|Tympnoscler-tymp/ossicle
C0395890|ICD9CM|PT|385.03|Tympanosclerosis involving tympanic membrane, ear ossicles, and middle ear
C0395890|ICD9CM|AB|385.03|Tympanoscler-all parts
C0395905|ICD9CM|AB|383.81|Postauricular fistula
C0395905|ICD9CM|PT|383.81|Postauricular fistula
C0395986|ICD9CM|PT|473.8|Other chronic sinusitis
C0395986|ICD9CM|AB|473.8|Chronic sinusitis NEC
C0396023|ICD9CM|AB|474.01|Chronic adenoiditis
C0396023|ICD9CM|PT|474.01|Chronic adenoiditis
C0396041|ICD9CM|PT|464.30|Acute epiglottitis without mention of obstruction
C0396041|ICD9CM|AB|464.30|Ac epiglottitis no obstr
C0396168|ICD9CM|PT|21.62|Fracture of the turbinates
C0396168|ICD9CM|AB|21.62|Turbinate fracture
C0396187|ICD9CM|PT|97.32|Removal of nasal packing
C0396187|ICD9CM|AB|97.32|Remove nasal packing
C0396200|ICD9CM|HT|22|Operations on nasal sinuses
C0396338|ICD9CM|PT|29.32|Pharyngeal diverticulectomy
C0396338|ICD9CM|AB|29.32|Pharyngeal diverticulec
C0396566|ICD9CM|AB|32.9|Other excision of lung
C0396566|ICD9CM|PT|32.9|Other excision of lung
C0396598|ICD9CM|PT|33.51|Unilateral lung transplantation
C0396598|ICD9CM|AB|33.51|Unilat lung transplant
C0396599|ICD9CM|PT|33.52|Bilateral lung transplantation
C0396599|ICD9CM|AB|33.52|Bilat lung transplant
C0396664|ICD9CM|HT|00.5|Other cardiovascular procedures
C0396814|ICD9CM|AB|38.22|Percutaneous angioscopy
C0396814|ICD9CM|PT|38.22|Percutaneous angioscopy
C0397314|ICD9CM|PT|35.53|Repair of ventricular septal defect with prosthesis, open technique
C0397314|ICD9CM|AB|35.53|Pros rep ventric def-opn
C0398053|ICD9CM|AB|39.31|Suture of artery
C0398053|ICD9CM|PT|39.31|Suture of artery
C0398341|ICD9CM|PT|99.76|Extracorporeal immunoadsorption
C0398341|ICD9CM|AB|99.76|Extracorp immunoabsorpt
C0398402|ICD9CM|PT|40.51|Radical excision of axillary lymph nodes
C0398402|ICD9CM|AB|40.51|Rad dissec axillary node
C0398404|ICD9CM|PT|40.52|Radical excision of periaortic lymph nodes
C0398404|ICD9CM|AB|40.52|Rad dissec periaort node
C0398530|ICD9CM|PT|41.09|Autologous bone marrow transplant with purging
C0398530|ICD9CM|AB|41.09|Auto bone mt w purging
C0398580|ICD9CM|PT|289.53|Neutropenic splenomegaly
C0398580|ICD9CM|AB|289.53|Neutropenic splenomegaly
C0398648|ICD9CM|PT|287.41|Posttransfusion purpura
C0398648|ICD9CM|AB|287.41|Posttransfusion purpura
C0398650|ICD9CM|PT|287.31|Immune thrombocytopenic purpura
C0398650|ICD9CM|AB|287.31|Immune thrombocyt purpra
C0398661|ICD9CM|PT|289.51|Chronic congestive splenomegaly
C0398661|ICD9CM|AB|289.51|Chr congest splenomegaly
C0398672|ICD9CM|PT|279.8|Other specified disorders involving the immune mechanism
C0398672|ICD9CM|AB|279.8|Immune mechanism dis NEC
C0399352|ICD9CM|AB|520.0|Anodontia
C0399352|ICD9CM|PT|520.0|Anodontia
C0399396|ICD9CM|PT|521.03|Dental caries extending into pulp
C0399396|ICD9CM|AB|521.03|Dental caries - pulp
C0399400|ICD9CM|PT|521.31|Erosion, limited to enamel
C0399400|ICD9CM|AB|521.31|Erosion-enamel
C0399408|ICD9CM|PT|522.3|Abnormal hard tissue formation in pulp
C0399408|ICD9CM|AB|522.3|Abn hard tiss-tooth pulp
C0399424|ICD9CM|AB|522.5|Periapical abscess
C0399424|ICD9CM|PT|522.5|Periapical abscess without sinus
C0399519|ICD9CM|AB|524.11|Maxillary asymmetry
C0399519|ICD9CM|PT|524.11|Anomalies of relationship of jaw to cranial base, maxillary asymmetry
C0399523|ICD9CM|PT|524.21|Malocclusion, Angle's class I
C0399523|ICD9CM|AB|524.21|Malocc- Angle's class I
C0399526|ICD9CM|PT|524.23|Malocclusion, Angle's class III
C0399526|ICD9CM|AB|524.23|Malocc-Angle's class III
C0399623|ICD9CM|PT|45.21|Transabdominal endoscopy of large intestine
C0399623|ICD9CM|AB|45.21|Transab lg bowel endosc
C0399857|ICD9CM|HT|46.9|Other operations on intestines
C0399857|ICD9CM|PT|46.99|Other operations on intestines
C0399857|ICD9CM|HT|46|Other operations on intestine
C0399857|ICD9CM|AB|46.99|Intestinal op NEC
C0399989|ICD9CM|AB|47.09|Other appendectomy
C0399989|ICD9CM|PT|47.09|Other appendectomy
C0400250|ICD9CM|PT|49.52|Posterior anal sphincterotomy
C0400250|ICD9CM|AB|49.52|Post sphincterotomy
C0400305|ICD9CM|PT|96.28|Manual reduction of enterostomy prolapse
C0400305|ICD9CM|AB|96.28|Manl reduct stoma prolap
C0400505|ICD9CM|PT|52.96|Anastomosis of pancreas
C0400505|ICD9CM|AB|52.96|Pancreatic anastomosis
C0400522|ICD9CM|PT|52.93|Endoscopic insertion of stent (tube) into pancreatic duct
C0400522|ICD9CM|AB|52.93|Endosc inser panc stent
C0400806|ICD9CM|PT|531.90|Gastric ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation, without mention of obstruction
C0400806|ICD9CM|AB|531.90|Stomach ulcer NOS
C0400806|ICD9CM|HT|531.9|Gastric ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation
C0400832|ICD9CM|PT|569.41|Ulcer of anus and rectum
C0400832|ICD9CM|AB|569.41|Rectal & anal ulcer
C0400853|ICD9CM|PT|777.2|Intestinal obstruction in newborn due to inspissated milk
C0400853|ICD9CM|AB|777.2|Intest obst-inspiss milk
C0400895|ICD9CM|AB|130.5|Toxoplasma hepatitis
C0400895|ICD9CM|PT|130.5|Hepatitis due to toxoplasmosis
C0400932|ICD9CM|PT|646.71|Liver and biliary tract disorders in pregnancy, delivered, with or without mention of antepartum condition
C0400932|ICD9CM|AB|646.71|Liver/bil trct disr-del
C0400985|ICD9CM|PT|574.00|Calculus of gallbladder with acute cholecystitis, without mention of obstruction
C0400985|ICD9CM|AB|574.00|Cholelith w ac cholecyst
C0401080|ICD9CM|PT|550.12|Inguinal hernia, with obstruction, without mention of gangrene, bilateral (not specified as recurrent)
C0401080|ICD9CM|AB|550.12|Bilat ing hernia w obst
C0401094|ICD9CM|PT|553.02|Femoral hernia without mention of obstruction or gangrene, bilateral (not specified as recurrent)
C0401094|ICD9CM|AB|553.02|Bilateral femoral hernia
C0401143|ICD9CM|PT|558.3|Allergic gastroenteritis and colitis
C0401143|ICD9CM|AB|558.3|Allrgic gastro & colitis
C0401161|ICD9CM|HT|55-59.99|OPERATIONS ON THE URINARY SYSTEM
C0401283|ICD9CM|AB|56.41|Partial ureterectomy
C0401283|ICD9CM|PT|56.41|Partial ureterectomy
C0401481|ICD9CM|PT|97.63|Removal of cystostomy tube
C0401481|ICD9CM|AB|97.63|Remov cystostomy tube
C0401640|ICD9CM|PT|60.11|Closed [percutaneous] [needle] biopsy of prostate
C0401640|ICD9CM|AB|60.11|Closed prostatic biopsy
C0403331|ICD9CM|PT|64.93|Division of penile adhesions
C0403331|ICD9CM|AB|64.93|Division of penile adhes
C0403334|ICD9CM|AB|99.95|Stretching of foreskin
C0403334|ICD9CM|PT|99.95|Stretching of foreskin
C0403529|ICD9CM|AB|446.21|Goodpasture's syndrome
C0403529|ICD9CM|PT|446.21|Goodpasture's syndrome
C0403645|ICD9CM|AB|596.4|Atony of bladder
C0403645|ICD9CM|PT|596.4|Atony of bladder
C0403673|ICD9CM|AB|608.87|Retrograde ejaculation
C0403673|ICD9CM|PT|608.87|Retrograde ejaculation
C0403696|ICD9CM|HT|598.0|Urethral stricture due to infection
C0403696|ICD9CM|PT|598.00|Urethral stricture due to unspecified infection
C0403696|ICD9CM|AB|598.00|Urethr strict:infect NOS
C0403698|ICD9CM|PT|598.1|Traumatic urethral stricture
C0403698|ICD9CM|AB|598.1|Traum urethral stricture
C0403719|ICD9CM|PT|274.11|Uric acid nephrolithiasis
C0403719|ICD9CM|AB|274.11|Uric acid nephrolithias
C0403853|ICD9CM|AB|71.62|Bilateral vulvectomy
C0403853|ICD9CM|PT|71.62|Bilateral vulvectomy
C0403929|ICD9CM|PT|70.4|Obliteration and total excision of vagina
C0403929|ICD9CM|AB|70.4|Vaginal obliteration
C0404009|ICD9CM|AB|70.12|Culdotomy
C0404009|ICD9CM|PT|70.12|Culdotomy
C0404050|ICD9CM|PT|67.0|Dilation of cervical canal
C0404050|ICD9CM|AB|67.0|Cervical canal dilation
C0404079|ICD9CM|HT|68.4|Total abdominal hysterectomy
C0404362|ICD9CM|PT|72.6|Forceps application to aftercoming head
C0404362|ICD9CM|AB|72.6|Forceps-aftercoming head
C0404458|ICD9CM|PT|614.4|Chronic or unspecified parametritis and pelvic cellulitis
C0404458|ICD9CM|AB|614.4|Chronic parametritis
C0404531|ICD9CM|AB|624.3|Hypertrophy of labia
C0404531|ICD9CM|PT|624.3|Hypertrophy of labia
C0404550|ICD9CM|PT|626.1|Scanty or infrequent menstruation
C0404550|ICD9CM|AB|626.1|Scanty menstruation
C0404572|ICD9CM|PT|628.0|Infertility, female, associated with anovulation
C0404572|ICD9CM|AB|628.0|Infertility-anovulation
C0404709|ICD9CM|HT|654.3|Retroverted and incarcerated gravid uterus
C0404725|ICD9CM|HT|648|Other current conditions in the mother classifiable elsewhere, but complicating pregnancy, childbirth, or the puerperium
C0404902|ICD9CM|PT|634.62|Spontaneous abortion, complicated by embolism, complete
C0404902|ICD9CM|AB|634.62|Spon abort w embol-comp
C0404903|ICD9CM|PT|634.52|Spontaneous abortion, complicated by shock, complete
C0404903|ICD9CM|AB|634.52|Spon abort w shock-comp
C0404905|ICD9CM|PT|634.32|Spontaneous abortion, complicated by renal failure, complete
C0404905|ICD9CM|AB|634.32|Spon ab w ren fail-comp
C0404919|ICD9CM|PT|634.61|Spontaneous abortion, complicated by embolism, incomplete
C0404919|ICD9CM|AB|634.61|Spon abort w embol-inc
C0404921|ICD9CM|PT|634.41|Spontaneous abortion, complicated by metabolic disorder, incomplete
C0404921|ICD9CM|AB|634.41|Spon ab w metab dis-inc
C0404922|ICD9CM|PT|634.31|Spontaneous abortion, complicated by renal failure, incomplete
C0404922|ICD9CM|AB|634.31|Spon ab w ren fail-inc
C0405011|ICD9CM|HT|653.7|Other fetal abnormality causing disproportion
C0405012|ICD9CM|HT|653.6|Hydrocephalic fetus causing disproportion
C0405034|ICD9CM|HT|658.9|Unspecified problem associated with amniotic cavity and membranes
C0405037|ICD9CM|PT|658.90|Unspecified problem associated with amniotic cavity and membranes, unspecified as to episode of care or not applicable
C0405037|ICD9CM|AB|658.90|Amniotic prob NOS-unspec
C0405072|ICD9CM|HT|646.4|Peripheral neuritis in pregnancy
C0405072|ICD9CM|PT|646.43|Peripheral neuritis in pregnancy, antepartum condition or complication
C0405072|ICD9CM|AB|646.43|Neuritis of preg-antepar
C0405080|ICD9CM|HT|643.1|Hyperemesis gravidarum with metabolic disturbance
C0405169|ICD9CM|HT|661.1|Secondary uterine inertia
C0405185|ICD9CM|HT|660.5|Locked twins
C0405189|ICD9CM|HT|659.1|Failed medical or unspecified induction of labor
C0405309|ICD9CM|PT|675.14|Abscess of breast associated with childbirth, postpartum condition or complication
C0405309|ICD9CM|AB|675.14|Breast abscess-postpart
C0405415|ICD9CM|AB|85.54|Bilateral breast implant
C0405415|ICD9CM|PT|85.54|Bilateral breast implant
C0405498|ICD9CM|HT|06|Operations on thyroid and parathyroid glands
C0405532|ICD9CM|PT|06.2|Unilateral thyroid lobectomy
C0405532|ICD9CM|AB|06.2|Unilat thyroid lobectomy
C0405540|ICD9CM|HT|06.5|Substernal thyroidectomy
C0405540|ICD9CM|PT|06.50|Substernal thyroidectomy, not otherwise specified
C0405540|ICD9CM|AB|06.50|Substern thyroidect NOS
C0405570|ICD9CM|HT|07.0|Exploration of adrenal field
C0405570|ICD9CM|PT|07.00|Exploration of adrenal field, not otherwise specified
C0405570|ICD9CM|AB|07.00|Adrenal exploration NOS
C0405578|ICD9CM|AB|253.0|Acromegaly and gigantism
C0405578|ICD9CM|PT|253.0|Acromegaly and gigantism
C0405580|ICD9CM|HT|255.4|Corticoadrenal insufficiency
C0405581|ICD9CM|HT|257|Testicular dysfunction
C0405581|ICD9CM|PT|257.9|Unspecified testicular dysfunction
C0405581|ICD9CM|AB|257.9|Testicular dysfunct NOS
C0405757|ICD9CM|PT|54.12|Reopening of recent laparotomy site
C0405757|ICD9CM|AB|54.12|Reopen recent lap site
C0405803|ICD9CM|PT|97.82|Removal of peritoneal drainage device
C0405803|ICD9CM|AB|97.82|Remov peritoneal drain
C0405808|ICD9CM|PT|54.51|Laparoscopic lysis of peritoneal adhesions
C0405808|ICD9CM|AB|54.51|Lap periton adhesiolysis
C0405902|ICD9CM|AB|34.26|Open mediastinal biopsy
C0405902|ICD9CM|PT|34.26|Open mediastinal biopsy
C0405910|ICD9CM|PT|34.79|Other repair of chest wall
C0405910|ICD9CM|AB|34.79|Other chest wall repair
C0405932|ICD9CM|PT|34.74|Repair of pectus deformity
C0405932|ICD9CM|AB|34.74|Pectus deformity repair
C0405992|ICD9CM|PT|34.20|Thoracoscopic pleural biopsy
C0405992|ICD9CM|AB|34.20|Thoracoscopic pleural bx
C0406047|ICD9CM|PT|686.9|Unspecified local infection of skin and subcutaneous tissue
C0406047|ICD9CM|AB|686.9|Local skin infection NOS
C0406078|ICD9CM|AB|682.4|Cellulitis of hand
C0406078|ICD9CM|PT|682.4|Cellulitis and abscess of hand, except fingers and thumb
C0406089|ICD9CM|PT|682.7|Cellulitis and abscess of foot, except toes
C0406089|ICD9CM|AB|682.7|Cellulitis of foot
C0406670|ICD9CM|HT|625.7|Vulvodynia
C0406670|ICD9CM|AB|625.70|Vulvodynia NOS
C0406670|ICD9CM|PT|625.70|Vulvodynia, unspecified
C0407093|ICD9CM|AB|83.12|Adductor tenotomy of hip
C0407093|ICD9CM|PT|83.12|Adductor tenotomy of hip
C0407183|ICD9CM|PT|83.93|Removal of skeletal muscle stimulator
C0407183|ICD9CM|AB|83.93|Remov skel musc stimulat
C0407232|ICD9CM|PT|79.19|Closed reduction of fracture with internal fixation, other specified bone
C0407232|ICD9CM|AB|79.19|Cl fx reduc-int fix NEC
C0407407|ICD9CM|PT|77.30|Other division of bone, unspecified site
C0407407|ICD9CM|HT|77.3|Other division of bone
C0407407|ICD9CM|AB|77.30|Other bone division NOS
C0407941|ICD9CM|AB|81.12|Triple arthrodesis
C0407941|ICD9CM|PT|81.12|Triple arthrodesis
C0408314|ICD9CM|AB|81.73|Total wrist replacement
C0408314|ICD9CM|PT|81.73|Total wrist replacement
C0408839|ICD9CM|AB|84.06|Disarticulation of elbow
C0408839|ICD9CM|PT|84.06|Disarticulation of elbow
C0408884|ICD9CM|HT|84.2|Reattachment of extremity
C0408885|ICD9CM|AB|84.24|Upper arm reattachment
C0408885|ICD9CM|PT|84.24|Upper arm reattachment
C0408894|ICD9CM|AB|84.22|Finger reattachment
C0408894|ICD9CM|PT|84.22|Finger reattachment
C0408900|ICD9CM|AB|84.26|Foot reattachment
C0408900|ICD9CM|PT|84.26|Foot reattachment
C0409209|ICD9CM|AB|716.93|Arthropathy NOS-forearm
C0409209|ICD9CM|PT|716.93|Arthropathy, unspecified, forearm
C0409215|ICD9CM|PT|716.89|Other specified arthropathy, multiple sites
C0409215|ICD9CM|AB|716.89|Arthropathy NEC-mult
C0409216|ICD9CM|PT|716.88|Other specified arthropathy, other specified sites
C0409216|ICD9CM|AB|716.88|Arthropathy NEC-oth site
C0409217|ICD9CM|PT|716.87|Other specified arthropathy, ankle and foot
C0409217|ICD9CM|AB|716.87|Arthropathy NEC-ankle
C0409218|ICD9CM|PT|716.86|Other specified arthropathy, lower leg
C0409218|ICD9CM|AB|716.86|Arthropathy NEC-l/leg
C0409219|ICD9CM|PT|716.85|Other specified arthropathy, pelvic region and thigh
C0409219|ICD9CM|AB|716.85|Arthropathy NEC-pelvis
C0409220|ICD9CM|PT|716.84|Other specified arthropathy, hand
C0409220|ICD9CM|AB|716.84|Arthropathy NEC-hand
C0409221|ICD9CM|PT|716.83|Other specified arthropathy, forearm
C0409221|ICD9CM|AB|716.83|Arthropathy NEC-forearm
C0409222|ICD9CM|PT|716.82|Other specified arthropathy, upper arm
C0409222|ICD9CM|AB|716.82|Arthropathy NEC-up/arm
C0409223|ICD9CM|PT|716.81|Other specified arthropathy, shoulder region
C0409223|ICD9CM|AB|716.81|Arthropathy NEC-shlder
C0409225|ICD9CM|PT|716.68|Unspecified monoarthritis, other specified sites
C0409225|ICD9CM|AB|716.68|Monoarthrit NOS-oth site
C0409226|ICD9CM|PT|716.67|Unspecified monoarthritis, ankle and foot
C0409226|ICD9CM|AB|716.67|Monoarthritis NOS-ankle
C0409227|ICD9CM|PT|716.66|Unspecified monoarthritis, lower leg
C0409227|ICD9CM|AB|716.66|Monoarthritis NOS-l/leg
C0409228|ICD9CM|PT|716.65|Unspecified monoarthritis, pelvic region and thigh
C0409228|ICD9CM|AB|716.65|Monoarthritis NOS-pelvis
C0409229|ICD9CM|PT|716.64|Unspecified monoarthritis, hand
C0409229|ICD9CM|AB|716.64|Monoarthritis NOS-hand
C0409230|ICD9CM|PT|716.63|Unspecified monoarthritis, forearm
C0409230|ICD9CM|AB|716.63|Monoarthrit NOS-forearm
C0409231|ICD9CM|PT|716.62|Unspecified monoarthritis, upper arm
C0409231|ICD9CM|AB|716.62|Monoarthritis NOS-up/arm
C0409232|ICD9CM|PT|716.61|Unspecified monoarthritis, shoulder region
C0409232|ICD9CM|AB|716.61|Monoarthritis NOS-shlder
C0409243|ICD9CM|PT|716.39|Climacteric arthritis, multiple sites
C0409243|ICD9CM|AB|716.39|Climact arthritis-mult
C0409244|ICD9CM|PT|716.38|Climacteric arthritis, other specified sites
C0409244|ICD9CM|AB|716.38|Climact arthritis NEC
C0409246|ICD9CM|PT|716.36|Climacteric arthritis, lower leg
C0409246|ICD9CM|AB|716.36|Climact arthritis-l/leg
C0409247|ICD9CM|PT|716.35|Climacteric arthritis, pelvic region and thigh
C0409247|ICD9CM|AB|716.35|Climact arthritis-pelvis
C0409248|ICD9CM|PT|716.34|Climacteric arthritis, hand
C0409248|ICD9CM|AB|716.34|Climact arthritis-hand
C0409249|ICD9CM|PT|716.33|Climacteric arthritis, forearm
C0409249|ICD9CM|AB|716.33|Climact arthrit-forearm
C0409250|ICD9CM|PT|716.32|Climacteric arthritis, upper arm
C0409250|ICD9CM|AB|716.32|Climact arthritis-up/arm
C0409251|ICD9CM|PT|716.31|Climacteric arthritis, shoulder region
C0409251|ICD9CM|AB|716.31|Climact arthritis-shlder
C0409252|ICD9CM|PT|716.29|Allergic arthritis, multiple sites
C0409252|ICD9CM|AB|716.29|Allerg arthritis-mult
C0409253|ICD9CM|PT|716.28|Allergic arthritis, other specified sites
C0409253|ICD9CM|AB|716.28|Allerg arthritis NEC
C0409254|ICD9CM|PT|716.27|Allergic arthritis, ankle and foot
C0409254|ICD9CM|AB|716.27|Allerg arthritis-ankle
C0409255|ICD9CM|PT|716.26|Allergic arthritis, lower leg
C0409255|ICD9CM|AB|716.26|Allerg arthritis-l/leg
C0409256|ICD9CM|PT|716.25|Allergic arthritis, pelvic region and thigh
C0409256|ICD9CM|AB|716.25|Allerg arthritis-pelvis
C0409257|ICD9CM|PT|716.24|Allergic arthritis, hand
C0409257|ICD9CM|AB|716.24|Allerg arthritis-hand
C0409258|ICD9CM|PT|716.23|Allergic arthritis, forearm
C0409258|ICD9CM|AB|716.23|Allerg arthritis-forearm
C0409259|ICD9CM|PT|716.22|Allergic arthritis, upper arm
C0409259|ICD9CM|AB|716.22|Allerg arthritis-up/arm
C0409260|ICD9CM|PT|716.21|Allergic arthritis, shoulder region
C0409260|ICD9CM|AB|716.21|Allerg arthritis-shlder
C0409264|ICD9CM|PT|719.97|Unspecified disorder of joint, ankle and foot
C0409264|ICD9CM|AB|719.97|Joint dis NOS-ankle
C0409271|ICD9CM|PT|718.99|Unspecified derangement of joint, multiple sites
C0409271|ICD9CM|AB|718.99|Jt derangement NOS-mult
C0409272|ICD9CM|PT|718.98|Unspecified derangement of joint, other specified sites
C0409272|ICD9CM|AB|718.98|Jt derangment NOS-oth jt
C0409273|ICD9CM|PT|718.97|Unspecified derangement of joint, ankle and foot
C0409273|ICD9CM|AB|718.97|Jt derangement NOS-ankle
C0409274|ICD9CM|PT|718.95|Unspecified derangement of joint, pelvic region and thigh
C0409274|ICD9CM|AB|718.95|Jt derangment NOS-pelvis
C0409275|ICD9CM|PT|718.94|Unspecified derangement of joint, hand
C0409275|ICD9CM|AB|718.94|Jt derangement NOS-hand
C0409276|ICD9CM|PT|718.93|Unspecified derangement of joint, forearm
C0409276|ICD9CM|AB|718.93|Jt derangmnt NOS-forearm
C0409277|ICD9CM|PT|718.92|Unspecified derangement of joint, upper arm
C0409277|ICD9CM|AB|718.92|Jt derangment NOS-up/arm
C0409278|ICD9CM|PT|718.91|Unspecified derangement of joint, shoulder region
C0409278|ICD9CM|AB|718.91|Jt derangment NOS-shlder
C0409415|ICD9CM|PT|718.31|Recurrent dislocation of joint, shoulder region
C0409415|ICD9CM|AB|718.31|Recur dislocat-shlder
C0409531|ICD9CM|PT|711.48|Arthropathy associated with other bacterial diseases, other specified sites
C0409531|ICD9CM|AB|711.48|Bact arthritis NEC
C0409532|ICD9CM|PT|711.49|Arthropathy associated with other bacterial diseases, multiple sites
C0409532|ICD9CM|AB|711.49|Bact arthritis-mult
C0409533|ICD9CM|PT|711.47|Arthropathy associated with other bacterial diseases, ankle and foot
C0409533|ICD9CM|AB|711.47|Bact arthritis-ankle
C0409534|ICD9CM|PT|711.46|Arthropathy associated with other bacterial diseases, lower leg
C0409534|ICD9CM|AB|711.46|Bact arthritis-l/leg
C0409535|ICD9CM|PT|711.45|Arthropathy associated with other bacterial diseases, pelvic region and thigh
C0409535|ICD9CM|AB|711.45|Bact arthritis-pelvis
C0409536|ICD9CM|PT|711.44|Arthropathy associated with other bacterial diseases, hand
C0409536|ICD9CM|AB|711.44|Bact arthritis-hand
C0409537|ICD9CM|PT|711.43|Arthropathy associated with other bacterial diseases, forearm
C0409537|ICD9CM|AB|711.43|Bact arthritis-forearm
C0409538|ICD9CM|PT|711.42|Arthropathy associated with other bacterial diseases, upper arm
C0409538|ICD9CM|AB|711.42|Bact arthritis-up/arm
C0409539|ICD9CM|PT|711.41|Arthropathy associated with other bacterial diseases, shoulder region
C0409539|ICD9CM|AB|711.41|Bact arthritis-shlder
C0409540|ICD9CM|PT|711.08|Pyogenic arthritis, other specified sites
C0409540|ICD9CM|AB|711.08|Pyogen arthritis NEC
C0409544|ICD9CM|PT|711.05|Pyogenic arthritis, pelvic region and thigh
C0409544|ICD9CM|AB|711.05|Pyogen arthritis-pelvis
C0409548|ICD9CM|PT|711.58|Arthropathy associated with other viral diseases, other specified sites
C0409548|ICD9CM|AB|711.58|Viral arthritis NEC
C0409549|ICD9CM|PT|711.59|Arthropathy associated with other viral diseases, multiple sites
C0409549|ICD9CM|AB|711.59|Viral arthritis-mult
C0409550|ICD9CM|PT|711.57|Arthropathy associated with other viral diseases, ankle and foot
C0409550|ICD9CM|AB|711.57|Viral arthritis-ankle
C0409551|ICD9CM|PT|711.56|Arthropathy associated with other viral diseases, lower leg
C0409551|ICD9CM|AB|711.56|Viral arthritis-l/leg
C0409552|ICD9CM|PT|711.55|Arthropathy associated with other viral diseases, pelvic region and thigh
C0409552|ICD9CM|AB|711.55|Viral arthritis-pelvis
C0409554|ICD9CM|PT|711.53|Arthropathy associated with other viral diseases, forearm
C0409554|ICD9CM|AB|711.53|Viral arthritis-forearm
C0409555|ICD9CM|PT|711.52|Arthropathy associated with other viral diseases, upper arm
C0409555|ICD9CM|AB|711.52|Viral arthritis-up/arm
C0409556|ICD9CM|PT|711.51|Arthropathy associated with other viral diseases, shoulder region
C0409556|ICD9CM|AB|711.51|Viral arthritis-shlder
C0409559|ICD9CM|PT|711.68|Arthropathy associated with mycoses, other specified sites
C0409559|ICD9CM|AB|711.68|Mycotic arthritis NEC
C0409561|ICD9CM|PT|711.67|Arthropathy associated with mycoses, ankle and foot
C0409561|ICD9CM|AB|711.67|Mycotic arthritis-ankle
C0409562|ICD9CM|PT|711.66|Arthropathy associated with mycoses, lower leg
C0409562|ICD9CM|AB|711.66|Mycotic arthritis-l/leg
C0409563|ICD9CM|PT|711.65|Arthropathy associated with mycoses, pelvic region and thigh
C0409563|ICD9CM|AB|711.65|Mycotic arthritis-pelvis
C0409564|ICD9CM|PT|711.64|Arthropathy associated with mycoses, hand
C0409564|ICD9CM|AB|711.64|Mycotic arthritis-hand
C0409565|ICD9CM|PT|711.63|Arthropathy associated with mycoses, forearm
C0409565|ICD9CM|AB|711.63|Mycotic arthrit-forearm
C0409566|ICD9CM|PT|711.62|Arthropathy associated with mycoses, upper arm
C0409566|ICD9CM|AB|711.62|Mycotic arthritis-up/arm
C0409567|ICD9CM|PT|711.61|Arthropathy associated with mycoses, shoulder region
C0409567|ICD9CM|AB|711.61|Mycotic arthritis-shlder
C0409569|ICD9CM|PT|711.70|Arthropathy associated with helminthiasis, site unspecified
C0409569|ICD9CM|AB|711.70|Helminth arthrit-unspec
C0409570|ICD9CM|PT|711.78|Arthropathy associated with helminthiasis, other specified sites
C0409570|ICD9CM|AB|711.78|Helminth arthrit NEC
C0409571|ICD9CM|PT|711.79|Arthropathy associated with helminthiasis, multiple sites
C0409571|ICD9CM|AB|711.79|Helminth arthrit-mult
C0409572|ICD9CM|AB|711.77|Helminth arthrit-ankle
C0409572|ICD9CM|PT|711.77|Arthropathy associated with helminthiasis, ankle and foot
C0409573|ICD9CM|PT|711.76|Arthropathy associated with helminthiasis, lower leg
C0409573|ICD9CM|AB|711.76|Helminth arthrit-l/leg
C0409574|ICD9CM|PT|711.75|Arthropathy associated with helminthiasis, pelvic region and thigh
C0409574|ICD9CM|AB|711.75|Helminth arthrit-pelvis
C0409575|ICD9CM|PT|711.74|Arthropathy associated with helminthiasis, hand
C0409575|ICD9CM|AB|711.74|Helminth arthrit-hand
C0409576|ICD9CM|PT|711.73|Arthropathy associated with helminthiasis, forearm
C0409576|ICD9CM|AB|711.73|Helminth arthrit-forearm
C0409577|ICD9CM|PT|711.72|Arthropathy associated with helminthiasis, upper arm
C0409577|ICD9CM|AB|711.72|Helminth arthrit-up/arm
C0409658|ICD9CM|PT|719.38|Palindromic rheumatism, other specified sites
C0409658|ICD9CM|AB|719.38|Palindrom rheum-jt NEC
C0409659|ICD9CM|PT|719.37|Palindromic rheumatism, ankle and foot
C0409659|ICD9CM|AB|719.37|Palindrom rheum-ankle
C0409660|ICD9CM|PT|719.36|Palindromic rheumatism, lower leg
C0409660|ICD9CM|AB|719.36|Palindrom rheum-l/leg
C0409661|ICD9CM|PT|719.35|Palindromic rheumatism, pelvic region and thigh
C0409661|ICD9CM|AB|719.35|Palindrom rheum-pelvis
C0409662|ICD9CM|PT|719.33|Palindromic rheumatism, forearm
C0409662|ICD9CM|AB|719.33|Palindrom rheum-forearm
C0409663|ICD9CM|PT|719.32|Palindromic rheumatism, upper arm
C0409663|ICD9CM|AB|719.32|Palindrom rheum-up/arm
C0409667|ICD9CM|HT|714.3|Juvenile chronic polyarthritis
C0409684|ICD9CM|PT|711.28|Arthropathy in Behcet's syndrome, other specified sites
C0409684|ICD9CM|AB|711.28|Behcet arthritis NEC
C0409685|ICD9CM|PT|711.29|Arthropathy in Behcet's syndrome, multiple sites
C0409685|ICD9CM|AB|711.29|Behcet arthritis-mult
C0409686|ICD9CM|PT|711.27|Arthropathy in Behcet's syndrome, ankle and foot
C0409686|ICD9CM|AB|711.27|Behcet arthritis-ankle
C0409687|ICD9CM|PT|711.26|Arthropathy in Behcet's syndrome, lower leg
C0409687|ICD9CM|AB|711.26|Behcet arthritis-l/leg
C0409688|ICD9CM|PT|711.25|Arthropathy in Behcet's syndrome, pelvic region and thigh
C0409688|ICD9CM|AB|711.25|Behcet arthritis-pelvis
C0409689|ICD9CM|PT|711.24|Arthropathy in Behcet's syndrome, hand
C0409689|ICD9CM|AB|711.24|Behcet arthritis-hand
C0409690|ICD9CM|PT|711.23|Arthropathy in Behcet's syndrome, forearm
C0409690|ICD9CM|AB|711.23|Behcet arthritis-forearm
C0409691|ICD9CM|PT|711.22|Arthropathy in Behcet's syndrome, upper arm
C0409691|ICD9CM|AB|711.22|Behcet arthritis-up/arm
C0409692|ICD9CM|PT|711.21|Arthropathy in Behcet's syndrome, shoulder region
C0409692|ICD9CM|AB|711.21|Behcet arthritis-shlder
C0409729|ICD9CM|PT|713.0|Arthropathy associated with other endocrine and metabolic disorders
C0409729|ICD9CM|AB|713.0|Arthrop w endocr/met dis
C0409752|ICD9CM|PT|716.19|Traumatic arthropathy, multiple sites
C0409752|ICD9CM|AB|716.19|Traum arthropathy-mult
C0409753|ICD9CM|PT|716.18|Traumatic arthropathy, other specified sites
C0409753|ICD9CM|AB|716.18|Traum arthropathy NEC
C0409754|ICD9CM|PT|716.17|Traumatic arthropathy, ankle and foot
C0409754|ICD9CM|AB|716.17|Traum arthropathy-ankle
C0409755|ICD9CM|PT|716.16|Traumatic arthropathy, lower leg
C0409755|ICD9CM|AB|716.16|Traum arthropathy-l/leg
C0409756|ICD9CM|PT|716.15|Traumatic arthropathy, pelvic region and thigh
C0409756|ICD9CM|AB|716.15|Traum arthropathy-pelvis
C0409757|ICD9CM|PT|716.14|Traumatic arthropathy, hand
C0409757|ICD9CM|AB|716.14|Traum arthropathy-hand
C0409758|ICD9CM|PT|716.13|Traumatic arthropathy, forearm
C0409758|ICD9CM|AB|716.13|Traum arthropath-forearm
C0409759|ICD9CM|PT|716.12|Traumatic arthropathy, upper arm
C0409759|ICD9CM|AB|716.12|Traum arthropathy-up/arm
C0409760|ICD9CM|PT|716.11|Traumatic arthropathy, shoulder region
C0409760|ICD9CM|AB|716.11|Traum arthropathy-shlder
C0409765|ICD9CM|PT|719.28|Villonodular synovitis, other specified sites
C0409765|ICD9CM|AB|719.28|Villonod synovit-jt NEC
C0409774|ICD9CM|PT|719.26|Villonodular synovitis, lower leg
C0409774|ICD9CM|AB|719.26|Villonod synovit-l/leg
C0409775|ICD9CM|PT|719.25|Villonodular synovitis, pelvic region and thigh
C0409775|ICD9CM|AB|719.25|Villonod synovit-pelvis
C0409780|ICD9CM|PT|719.24|Villonodular synovitis, hand
C0409780|ICD9CM|AB|719.24|Villonod synovit-hand
C0409784|ICD9CM|PT|719.23|Villonodular synovitis, forearm
C0409784|ICD9CM|AB|719.23|Villonod synovit-forearm
C0409787|ICD9CM|PT|719.22|Villonodular synovitis, upper arm
C0409787|ICD9CM|AB|719.22|Villonod synovit-up/arm
C0409809|ICD9CM|PT|716.49|Transient arthropathy, multiple sites
C0409809|ICD9CM|AB|716.49|Trans arthropathy-mult
C0409810|ICD9CM|PT|716.48|Transient arthropathy, other specified sites
C0409810|ICD9CM|AB|716.48|Trans arthropathy NEC
C0409811|ICD9CM|PT|716.47|Transient arthropathy, ankle and foot
C0409811|ICD9CM|AB|716.47|Trans arthropathy-ankle
C0409812|ICD9CM|PT|716.46|Transient arthropathy, lower leg
C0409812|ICD9CM|AB|716.46|Trans arthropathy-l/leg
C0409813|ICD9CM|PT|716.45|Transient arthropathy, pelvic region and thigh
C0409813|ICD9CM|AB|716.45|Trans arthropathy-pelvis
C0409814|ICD9CM|PT|716.44|Transient arthropathy, hand
C0409814|ICD9CM|AB|716.44|Trans arthropathy-hand
C0409815|ICD9CM|PT|716.43|Transient arthropathy, forearm
C0409815|ICD9CM|AB|716.43|Trans arthropath-forearm
C0409816|ICD9CM|PT|716.42|Transient arthropathy, upper arm
C0409816|ICD9CM|AB|716.42|Trans arthropathy-up/arm
C0409843|ICD9CM|PT|712.95|Unspecified crystal arthropathy, pelvic region and thigh
C0409843|ICD9CM|AB|712.95|Cryst arthrop NOS-pelvis
C0409862|ICD9CM|PT|712.28|Chondrocalcinosis, due to pyrophosphate crystals, other specified sites
C0409862|ICD9CM|AB|712.28|Pyrophos cryst-site NEC
C0409863|ICD9CM|PT|712.29|Chondrocalcinosis, due to pyrophosphate crystals, multiple sites
C0409863|ICD9CM|AB|712.29|Pyrophos cryst-mult
C0409864|ICD9CM|PT|712.27|Chondrocalcinosis, due to pyrophosphate crystals, ankle and foot
C0409864|ICD9CM|AB|712.27|Pyrophosph cryst-ankle
C0409865|ICD9CM|PT|712.26|Chondrocalcinosis, due to pyrophosphate crystals, lower leg
C0409865|ICD9CM|AB|712.26|Pyrophosph cryst-l/leg
C0409867|ICD9CM|PT|712.25|Chondrocalcinosis, due to pyrophosphate crystals, pelvic region and thigh
C0409867|ICD9CM|AB|712.25|Pyrophosph cryst-pelvis
C0409868|ICD9CM|AB|712.24|Pyrophosph cryst-hand
C0409868|ICD9CM|PT|712.24|Chondrocalcinosis, due to pyrophosphate crystals, hand
C0409869|ICD9CM|PT|712.23|Chondrocalcinosis, due to pyrophosphate crystals, forearm
C0409869|ICD9CM|AB|712.23|Pyrophosph cryst-forearm
C0409870|ICD9CM|PT|712.22|Chondrocalcinosis, due to pyrophosphate crystals, upper arm
C0409870|ICD9CM|AB|712.22|Pyrophosph cryst-up/arm
C0409871|ICD9CM|PT|712.21|Chondrocalcinosis, due to pyrophosphate crystals, shoulder region
C0409871|ICD9CM|AB|712.21|Pyrophosph cryst-shlder
C0409873|ICD9CM|PT|712.18|Chondrocalcinosis, due to dicalcium phosphate crystals, other specified sites
C0409873|ICD9CM|AB|712.18|Dicalc phos cry-site NEC
C0409874|ICD9CM|PT|712.19|Chondrocalcinosis, due to dicalcium phosphate crystals, multiple sites
C0409874|ICD9CM|AB|712.19|Dicalc phos cryst-mult
C0409875|ICD9CM|PT|712.17|Chondrocalcinosis, due to dicalcium phosphate crystals, ankle and foot
C0409875|ICD9CM|AB|712.17|Dicalc phos cryst-ankle
C0409876|ICD9CM|PT|712.16|Chondrocalcinosis, due to dicalcium phosphate crystals, lower leg
C0409876|ICD9CM|AB|712.16|Dicalc phos cryst-l/leg
C0409877|ICD9CM|PT|712.15|Chondrocalcinosis, due to dicalcium phosphate crystals, pelvic region and thigh
C0409877|ICD9CM|AB|712.15|Dicalc phos cryst-pelvis
C0409878|ICD9CM|PT|712.14|Chondrocalcinosis, due to dicalcium phosphate crystals, hand
C0409878|ICD9CM|AB|712.14|Dicalc phos cryst-hand
C0409879|ICD9CM|PT|712.13|Chondrocalcinosis, due to dicalcium phosphate crystals, forearm
C0409879|ICD9CM|AB|712.13|Dicalc phos crys-forearm
C0409880|ICD9CM|PT|712.12|Chondrocalcinosis, due to dicalcium phosphate crystals, upper arm
C0409880|ICD9CM|AB|712.12|Dicalc phos cryst-up/arm
C0409881|ICD9CM|PT|712.11|Chondrocalcinosis, due to dicalcium phosphate crystals, shoulder region
C0409881|ICD9CM|AB|712.11|Dicalc phos cryst-shlder
C0409882|ICD9CM|PT|712.10|Chondrocalcinosis, due to dicalcium phosphate crystals, site unspecified
C0409882|ICD9CM|AB|712.10|Dicalc phos cryst-unspec
C0409886|ICD9CM|PT|712.38|Chondrocalcinosis, unspecified, other specified sites
C0409886|ICD9CM|AB|712.38|Chondrocalc NOS-oth site
C0409887|ICD9CM|PT|712.39|Chondrocalcinosis, unspecified, multiple sites
C0409887|ICD9CM|AB|712.39|Chondrocalcin NOS-mult
C0409888|ICD9CM|PT|712.37|Chondrocalcinosis, unspecified, ankle and foot
C0409888|ICD9CM|AB|712.37|Chondrocalcin NOS-ankle
C0409889|ICD9CM|PT|712.36|Chondrocalcinosis, unspecified, lower leg
C0409889|ICD9CM|AB|712.36|Chondrocalcin NOS-l/leg
C0409890|ICD9CM|PT|712.35|Chondrocalcinosis, unspecified, pelvic region and thigh
C0409890|ICD9CM|AB|712.35|Chondrocalcin NOS-pelvis
C0409891|ICD9CM|PT|712.34|Chondrocalcinosis, unspecified, hand
C0409891|ICD9CM|AB|712.34|Chondrocalcin NOS-hand
C0409892|ICD9CM|PT|712.33|Chondrocalcinosis, unspecified, forearm
C0409892|ICD9CM|AB|712.33|Chondrocalc NOS-forearm
C0409893|ICD9CM|PT|712.32|Chondrocalcinosis, unspecified, upper arm
C0409893|ICD9CM|AB|712.32|Chondrocalcin NOS-up/arm
C0409894|ICD9CM|PT|712.31|Chondrocalcinosis, unspecified, shoulder region
C0409894|ICD9CM|AB|712.31|Chondrocalcin NOS-shlder
C0409968|ICD9CM|PT|716.08|Kaschin-Beck disease, other specified sites
C0409968|ICD9CM|AB|716.08|Kaschin-beck dis NEC
C0409969|ICD9CM|PT|716.07|Kaschin-Beck disease, ankle and foot
C0409969|ICD9CM|AB|716.07|Kaschin-beck dis-ankle
C0409970|ICD9CM|PT|716.05|Kaschin-Beck disease, pelvic region and thigh
C0409970|ICD9CM|AB|716.05|Kaschin-beck dis-pelvis
C0409974|ICD9CM|AB|695.4|Lupus erythematosus
C0409974|ICD9CM|PT|695.4|Lupus erythematosus
C0410017|ICD9CM|PT|727.61|Complete rupture of rotator cuff
C0410017|ICD9CM|AB|727.61|Rotator cuff rupture
C0410224|ICD9CM|PT|359.29|Other specified myotonic disorder
C0410224|ICD9CM|AB|359.29|Myotonic disorder NEC
C0410318|ICD9CM|PT|730.79|Osteopathy resulting from poliomyelitis, multiple sites
C0410318|ICD9CM|AB|730.79|Polio osteopathy-mult
C0410319|ICD9CM|PT|730.78|Osteopathy resulting from poliomyelitis, other specified sites
C0410319|ICD9CM|AB|730.78|Polio osteopathy NEC
C0410320|ICD9CM|PT|730.77|Osteopathy resulting from poliomyelitis, ankle and foot
C0410320|ICD9CM|AB|730.77|Polio osteopathy-ankle
C0410321|ICD9CM|PT|730.76|Osteopathy resulting from poliomyelitis, lower leg
C0410321|ICD9CM|AB|730.76|Polio osteopathy-l/leg
C0410322|ICD9CM|PT|730.75|Osteopathy resulting from poliomyelitis, pelvic region and thigh
C0410322|ICD9CM|AB|730.75|Polio osteopathy-pelvis
C0410323|ICD9CM|AB|730.74|Polio osteopathy-hand
C0410323|ICD9CM|PT|730.74|Osteopathy resulting from poliomyelitis, hand
C0410324|ICD9CM|AB|730.73|Polio osteopathy-forearm
C0410324|ICD9CM|PT|730.73|Osteopathy resulting from poliomyelitis, forearm
C0410325|ICD9CM|PT|730.72|Osteopathy resulting from poliomyelitis, upper arm
C0410325|ICD9CM|AB|730.72|Polio osteopathy-up/arm
C0410326|ICD9CM|PT|730.71|Osteopathy resulting from poliomyelitis, shoulder region
C0410326|ICD9CM|AB|730.71|Polio osteopathy-shlder
C0410331|ICD9CM|PT|718.08|Articular cartilage disorder, other specified sites
C0410331|ICD9CM|AB|718.08|Artic cartil dis-jt NEC
C0410332|ICD9CM|PT|718.05|Articular cartilage disorder, pelvic region and thigh
C0410332|ICD9CM|AB|718.05|Artic cartil dis-pelvis
C0410376|ICD9CM|PT|730.28|Unspecified osteomyelitis, other specified sites
C0410376|ICD9CM|AB|730.28|Osteomyelit NOS-oth site
C0410385|ICD9CM|PT|730.08|Acute osteomyelitis, other specified sites
C0410385|ICD9CM|AB|730.08|Ac osteomyelitis NEC
C0410417|ICD9CM|PT|730.18|Chronic osteomyelitis, other specified sites
C0410417|ICD9CM|AB|730.18|Chr osteomyelit NEC
C0410420|ICD9CM|PT|730.15|Chronic osteomyelitis, pelvic region and thigh
C0410420|ICD9CM|AB|730.15|Chr osteomyelit-pelvis
C0410434|ICD9CM|PT|730.38|Periostitis, without mention of osteomyelitis, other specified sites
C0410434|ICD9CM|AB|730.38|Periostitis NEC
C0410435|ICD9CM|PT|730.35|Periostitis, without mention of osteomyelitis, pelvic region and thigh
C0410435|ICD9CM|AB|730.35|Periostitis-pelvis
C0410436|ICD9CM|PT|730.31|Periostitis, without mention of osteomyelitis, shoulder region
C0410436|ICD9CM|AB|730.31|Periostitis-shlder
C0410437|ICD9CM|PT|730.30|Periostitis, without mention of osteomyelitis, site unspecified
C0410437|ICD9CM|AB|730.30|Periostitis-unspec
C0410502|ICD9CM|PT|732.1|Juvenile osteochondrosis of hip and pelvis
C0410502|ICD9CM|AB|732.1|Juv osteochondros pelvis
C0410632|ICD9CM|HT|722.3|Schmorl's nodes
C0410632|ICD9CM|AB|722.30|Schmorl's nodes NOS
C0410632|ICD9CM|PT|722.30|Schmorl's nodes, unspecified region
C0410693|ICD9CM|PT|737.8|Other curvatures of spine
C0410693|ICD9CM|AB|737.8|Curvature of spine NEC
C0410740|ICD9CM|PT|736.20|Unspecified deformity of finger
C0410740|ICD9CM|AB|736.20|Acq finger deformity NOS
C0410779|ICD9CM|AB|735.3|Hallux malleus
C0410779|ICD9CM|PT|735.3|Hallux malleus
C0410807|ICD9CM|PT|996.42|Dislocation of prosthetic joint
C0410807|ICD9CM|AB|996.42|Dislocate prosthetic jt
C0411063|ICD9CM|PT|767.4|Injury to spine and spinal cord due to birth trauma
C0411063|ICD9CM|AB|767.4|Spinal cord inj at birth
C0411160|ICD9CM|PT|761.1|Premature rupture of membranes affecting fetus or newborn
C0411160|ICD9CM|AB|761.1|Premat rupt memb aff NB
C0411164|ICD9CM|PT|761.4|Ectopic pregnancy affecting fetus or newborn
C0411164|ICD9CM|AB|761.4|Ectopic pregnancy aff NB
C0411169|ICD9CM|PT|761.5|Multiple pregnancy affecting fetus or newborn
C0411169|ICD9CM|AB|761.5|Mult pregnancy aff NB
C0411175|ICD9CM|PT|760.9|Unspecified maternal condition affecting fetus or newborn
C0411175|ICD9CM|AB|760.9|Maternal cond NOS aff NB
C0411176|ICD9CM|PT|760.0|Maternal hypertensive disorders affecting fetus or newborn
C0411176|ICD9CM|AB|760.0|Matern hyperten aff NB
C0411178|ICD9CM|PT|760.2|Maternal infections affecting fetus or newborn
C0411178|ICD9CM|AB|760.2|Maternal infec aff NB
C0411268|ICD9CM|PT|007.3|Intestinal trichomoniasis
C0411268|ICD9CM|AB|007.3|Intest trichomoniasis
C0411279|ICD9CM|PT|126.9|Ancylostomiasis and necatoriasis, unspecified
C0411279|ICD9CM|AB|126.9|Ancylostomiasis NOS
C0411279|ICD9CM|HT|126|Ancylostomiasis and necatoriasis
C0411665|ICD9CM|AB|18.01|Piercing of ear lobe
C0411665|ICD9CM|PT|18.01|Piercing of ear lobe
C0412048|ICD9CM|PT|88.46|Arteriography of placenta
C0412048|ICD9CM|AB|88.46|Contrast placentogram
C0412112|ICD9CM|AB|87.63|Small bowel series
C0412112|ICD9CM|PT|87.63|Small bowel series
C0412201|ICD9CM|PT|87.38|Sinogram of chest wall
C0412201|ICD9CM|AB|87.38|Chest wall sinogram
C0412375|ICD9CM|PT|92.16|Scan of lymphatic system
C0412375|ICD9CM|AB|92.16|Lymphatic system scan
C0412412|ICD9CM|PT|92.03|Renal scan and radioisotope function study
C0412412|ICD9CM|AB|92.03|Renal scan/isotope funct
C0412512|ICD9CM|AB|95.13|Ultrasound study of eye
C0412512|ICD9CM|PT|95.13|Ultrasound study of eye
C0412527|ICD9CM|PT|88.77|Diagnostic ultrasound of peripheral vascular system
C0412527|ICD9CM|AB|88.77|Dx ultrasound-vascular
C0412620|ICD9CM|PT|88.01|Computerized axial tomography of abdomen
C0412620|ICD9CM|AB|88.01|C.A.T. scan of abdomen
C0412623|ICD9CM|PT|87.71|Computerized axial tomography of kidney
C0412623|ICD9CM|AB|87.71|C.A.T. scan of kidney
C0412675|ICD9CM|PT|88.91|Magnetic resonance imaging of brain and brain stem
C0412675|ICD9CM|AB|88.91|Mri of brain & brainstem
C0412755|ICD9CM|HT|88|Other diagnostic radiology and related techniques
C0412836|ICD9CM|PT|963.1|Poisoning by antineoplastic and immunosuppressive drugs
C0412836|ICD9CM|AB|963.1|Pois-antineopl/immunosup
C0412842|ICD9CM|PT|964.0|Poisoning by iron and its compounds
C0412842|ICD9CM|AB|964.0|Poisoning-iron/compounds
C0412845|ICD9CM|PT|964.4|Poisoning by fibrinolysis-affecting drugs
C0412845|ICD9CM|AB|964.4|Poison-fibrinolysis agnt
C0412862|ICD9CM|PT|969.4|Poisoning by benzodiazepine-based tranquilizers
C0412862|ICD9CM|AB|969.4|Pois-benzodiazepine tran
C0412869|ICD9CM|PT|970.89|Poisoning by other central nervous system stimulants
C0412869|ICD9CM|AB|970.89|Poison-CNS stimulant NEC
C0412870|ICD9CM|PT|971.1|Poisoning by parasympatholytics (anticholinergics and antimuscarinics) and spasmolytics
C0412870|ICD9CM|AB|971.1|Pois-parasympatholytics
C0412873|ICD9CM|PT|972.0|Poisoning by cardiac rhythm regulators
C0412873|ICD9CM|AB|972.0|Pois-card rhythm regulat
C0412909|ICD9CM|HT|977|Poisoning by other and unspecified drugs and medicinal substances
C0412915|ICD9CM|PT|978.1|Poisoning by typhoid and paratyphoid vaccine
C0412915|ICD9CM|AB|978.1|Pois-typh/paratyph vacc
C0412916|ICD9CM|PT|978.6|Poisoning by pertussis vaccine, including combinations with a pertussis component
C0412916|ICD9CM|AB|978.6|Pois-pertussis vaccine
C0412917|ICD9CM|PT|978.9|Poisoning by mixed bacterial vaccines, except combinations with a pertussis component
C0412917|ICD9CM|AB|978.9|Pois-mix bacter vaccines
C0412928|ICD9CM|HT|966|Poisoning by anticonvulsants and anti-Parkinsonism drugs
C0412954|ICD9CM|PT|982.3|Toxic effect of other chlorinated hydrocarbon solvents
C0412954|ICD9CM|AB|982.3|Tx ef cl-hydcarb slv NEC
C0412991|ICD9CM|PT|985.2|Toxic effect of manganese and its compounds
C0412991|ICD9CM|AB|985.2|Toxic effect manganese
C0412992|ICD9CM|PT|985.3|Toxic effect of beryllium and its compounds
C0412992|ICD9CM|AB|985.3|Toxic effect beryllium
C0412994|ICD9CM|PT|985.5|Toxic effect of cadmium and its compounds
C0412994|ICD9CM|AB|985.5|Toxic effect cadmium
C0413000|ICD9CM|HT|987|Toxic effect of other gases, fumes, or vapors
C0413004|ICD9CM|PT|987.1|Toxic effect of other hydrocarbon gas
C0413004|ICD9CM|AB|987.1|Tox ef hydrocarb gas NEC
C0413005|ICD9CM|PT|987.0|Toxic effect of liquefied petroleum gases
C0413005|ICD9CM|AB|987.0|Toxic eff liq petrol gas
C0413040|ICD9CM|PT|989.3|Toxic effect of organophosphate and carbamate
C0413040|ICD9CM|AB|989.3|Tox eff organphos/carbam
C0413252|ICD9CM|AB|991.6|Hypothermia
C0413252|ICD9CM|PT|991.6|Hypothermia
C0413443|ICD9CM|PT|E930.0|Penicillins causing adverse effects in therapeutic use
C0413443|ICD9CM|AB|E930.0|Adv eff penicillins
C0413512|ICD9CM|PT|E931.6|Anthelmintics causing adverse effects in therapeutic use
C0413512|ICD9CM|AB|E931.6|Adv eff anthelmintics
C0413956|ICD9CM|PT|E943.9|Unspecified agent primarily affecting the gastrointestinal system causing adverse effects in therapeutic use
C0413956|ICD9CM|HT|E943|Agents primarily affecting gastrointestinal system causing adverse effects in therapeutic use
C0413956|ICD9CM|AB|E943.9|Adv eff GI agent NOS
C0414020|ICD9CM|PT|E945.0|Oxytocic agents causing adverse effects in therapeutic use
C0414020|ICD9CM|AB|E945.0|Adv eff oxytocic agents
C0414040|ICD9CM|PT|E945.6|Anti-common cold drugs causing adverse effects in therapeutic use
C0414040|ICD9CM|AB|E945.6|Adv eff anti-common cold
C0414053|ICD9CM|PT|E946.2|Local astringents and local detergents causing adverse effects in therapeutic use
C0414053|ICD9CM|AB|E946.2|Adv eff local astringent
C0414054|ICD9CM|PT|E946.3|Emollients, demulcents, and protectants causing adverse effects in therapeutic use
C0414054|ICD9CM|AB|E946.3|Adv eff emollient/demulc
C0414055|ICD9CM|PT|E946.4|Keratolytics, keratoplastics, other hair treatment drugs and preparations causing adverse effects in therapeutic use
C0414055|ICD9CM|AB|E946.4|Adv eff hair/scalp prep
C0414085|ICD9CM|HT|E800-E807.9|RAILWAY ACCIDENTS
C0414085|ICD9CM|HT|E807|Railway accident of unspecified nature
C0414276|ICD9CM|HT|E804|Fall in, on, or from railway train
C0414277|ICD9CM|PT|E804.9|Fall in, on, or from railway train injuring unspecified person
C0414277|ICD9CM|AB|E804.9|Fall from train-pers NOS
C0414278|ICD9CM|PT|E804.8|Fall in, on, or from railway train injuring other specified person
C0414278|ICD9CM|AB|E804.8|Fall from train-pers NEC
C0414279|ICD9CM|PT|E804.3|Fall in, on, or from railway train injuring pedal cyclist
C0414279|ICD9CM|AB|E804.3|Fall from train-ped cycl
C0414280|ICD9CM|PT|E804.2|Fall in, on, or from railway train injuring pedestrian
C0414280|ICD9CM|AB|E804.2|Fall from train-pedest
C0414282|ICD9CM|PT|E804.0|Fall in, on, or from railway train injuring railway employee
C0414282|ICD9CM|AB|E804.0|Fall on/from train-empl
C0414302|ICD9CM|HT|E805|Hit by rolling stock
C0414364|ICD9CM|PT|E829.8|Other road vehicle accidents injuring other specified person
C0414364|ICD9CM|AB|E829.8|Oth rd veh acc-pers NEC
C0414438|ICD9CM|PT|E810.9|Motor vehicle traffic accident involving collision with train injuring unspecified person
C0414438|ICD9CM|HT|E810|Motor vehicle traffic accident involving collision with train
C0414438|ICD9CM|AB|E810.9|Mv-train coll-pers NOS
C0414439|ICD9CM|PT|E810.8|Motor vehicle traffic accident involving collision with train injuring other specified person
C0414439|ICD9CM|AB|E810.8|Mv-train coll-pers NEC
C0414440|ICD9CM|PT|E810.7|Motor vehicle traffic accident involving collision with train injuring pedestrian
C0414440|ICD9CM|AB|E810.7|Mv-train coll-pedest
C0414441|ICD9CM|PT|E810.6|Motor vehicle traffic accident involving collision with train injuring pedal cyclist
C0414441|ICD9CM|AB|E810.6|Mv-train coll-ped cycl
C0414471|ICD9CM|PT|E813.9|Motor vehicle traffic accident involving collision with other vehicle injuring unspecified person
C0414471|ICD9CM|AB|E813.9|Mv-oth veh coll-pers NOS
C0414494|ICD9CM|PT|E811.7|Motor vehicle traffic accident involving re-entrant collision with another motor vehicle injuring pedestrian
C0414494|ICD9CM|AB|E811.7|Reentrant coll-pedest
C0414733|ICD9CM|PT|E816.9|Motor vehicle traffic accident due to loss of control, without collision on the highway, injuring unspecified person
C0414733|ICD9CM|AB|E816.9|Loss control mv-pers NOS
C0414734|ICD9CM|PT|E816.8|Motor vehicle traffic accident due to loss of control, without collision on the highway, injuring other specified person
C0414734|ICD9CM|AB|E816.8|Loss control mv-pers NEC
C0414735|ICD9CM|PT|E816.7|Motor vehicle traffic accident due to loss of control, without collision on the highway, injuring pedestrian
C0414735|ICD9CM|AB|E816.7|Loss control mv-pedest
C0414736|ICD9CM|PT|E816.6|Motor vehicle traffic accident due to loss of control, without collision on the highway, injuring pedal cyclist
C0414736|ICD9CM|AB|E816.6|Loss control mv-ped cycl
C0414740|ICD9CM|PT|E816.2|Motor vehicle traffic accident due to loss of control, without collision on the highway, injuring motorcyclist
C0414740|ICD9CM|AB|E816.2|Loss control mv-mocycl
C0415270|ICD9CM|HT|E820|Nontraffic accident involving motor-driven snow vehicle
C0415505|ICD9CM|PT|E826.3|Pedal cycle accident injuring occupant of animal-drawn vehicle
C0415505|ICD9CM|AB|E826.3|Ped cyc acc-occ anim veh
C0415658|ICD9CM|PT|E828.2|Accident involving animal being ridden injuring rider of animal
C0415658|ICD9CM|AB|E828.2|Ridden animal acc-rider
C0415659|ICD9CM|PT|E828.0|Accident involving animal being ridden injuring pedestrian
C0415659|ICD9CM|AB|E828.0|Ridden animal acc-pedest
C0416143|ICD9CM|HT|E841|Accident to powered aircraft, other and unspecified
C0416348|ICD9CM|PT|E842.7|Accident to unpowered aircraft injuring parachutist (military) (other)
C0416348|ICD9CM|AB|E842.7|Unpow aircrf acc-chutist
C0416598|ICD9CM|PT|E850.6|Accidental poisoning by antirheumatics (antiphlogistics)
C0416598|ICD9CM|AB|E850.6|Acc poison-antirheumatic
C0416665|ICD9CM|PT|E855.3|Accidental poisoning by parasympathomimetics [cholinergics]
C0416665|ICD9CM|AB|E855.3|Acc poison-cholinergics
C0416674|ICD9CM|PT|E855.5|Accidental poisoning by sympathomimetics [adrenergics]
C0416674|ICD9CM|AB|E855.5|Acc poison-adrenergics
C0416678|ICD9CM|PT|E855.6|Accidental poisoning by sympatholytics [antiadrenergics]
C0416678|ICD9CM|AB|E855.6|Acc poisn-sympatholytics
C0416707|ICD9CM|PT|E861.3|Accidental poisoning by other cleansing and polishing agents
C0416707|ICD9CM|AB|E861.3|Acc poison-cleanser NEC
C0416786|ICD9CM|PT|E865.0|Accidental poisoning by meat
C0416786|ICD9CM|AB|E865.0|Acc poison-meat
C0416882|ICD9CM|PT|E862.1|Accidental poisoning by petroleum fuels and cleaners
C0416882|ICD9CM|AB|E862.1|Acc poisn-petroleum fuel
C0416973|ICD9CM|PT|E869.3|Accidental poisoning by lacrimogenic gas [tear gas]
C0416973|ICD9CM|AB|E869.3|Acc poison-tear gas
C0416980|ICD9CM|PT|E888.8|Other fall
C0416980|ICD9CM|AB|E888.8|Fall NEC
C0417007|ICD9CM|HT|E886|Fall on same level from collision, pushing, or shoving, by or with other person
C0417080|ICD9CM|PT|E896|Accident caused by controlled fire in other and unspecified building or structure
C0417080|ICD9CM|AB|E896|Burn acc in bldg NEC
C0417090|ICD9CM|PT|E891.8|Other accident resulting from conflagration in other and unspecified building or structure
C0417090|ICD9CM|AB|E891.8|Fire in bldg-accid NEC
C0417282|ICD9CM|PT|E890.1|Fumes from combustion of polyvinylchloride [pvc] and similar material in conflagration in private dwelling
C0417282|ICD9CM|AB|E890.1|Priv dwel fire-pvc fumes
C0417413|ICD9CM|PT|E893.9|Accident caused by ignition of clothing by unspecified source
C0417413|ICD9CM|AB|E893.9|Clothing fire NOS
C0417424|ICD9CM|PT|E893.0|Accident caused by ignition of clothing from controlled fire in private dwelling
C0417424|ICD9CM|AB|E893.0|Clothing fire-priv dwell
C0417496|ICD9CM|PT|E898.0|Accident caused by burning bedclothes
C0417496|ICD9CM|AB|E898.0|Burning bedclothes
C0417584|ICD9CM|PT|E904.9|Accident due to privation, unqualified
C0417584|ICD9CM|AB|E904.9|Privation NOS
C0417614|ICD9CM|PT|E909.0|Earthquakes
C0417614|ICD9CM|AB|E909.0|Acc d/t earthquakes
C0417672|ICD9CM|PT|E904.1|Accident due to lack of food
C0417672|ICD9CM|AB|E904.1|Lack of food
C0417673|ICD9CM|PT|E904.2|Accident due to lack of water
C0417673|ICD9CM|AB|E904.2|Lack of water
C0417758|ICD9CM|HT|E906|Other injury caused by animals
C0417794|ICD9CM|PT|E910.1|Accidental drowning and submersion while engaged in other sport or recreational activity with diving equipment
C0417794|ICD9CM|AB|E910.1|Skin/scuba diving acc
C0418343|ICD9CM|PT|E968.4|Assault by criminal neglect
C0418343|ICD9CM|AB|E968.4|Assault-criminal neglect
C0418380|ICD9CM|PT|E965.6|Assault by gasoline bomb
C0418380|ICD9CM|AB|E965.6|Assault-gasoline bomb
C0418384|ICD9CM|PT|E966|Assault by cutting and piercing instrument
C0418384|ICD9CM|AB|E966|Assault-cutting instr
C0418414|ICD9CM|PT|E968.7|Assault by human bite
C0418414|ICD9CM|AB|E968.7|Human bite - assault
C0418456|ICD9CM|AB|E969|Late effect assault
C0418456|ICD9CM|PT|E969|Late effects of injury purposely inflicted by other person
C0418479|ICD9CM|PT|E974|Injury due to legal intervention by cutting and piercing instrument
C0418479|ICD9CM|AB|E974|Legal interven-cut instr
C0418593|ICD9CM|PT|E876.9|Unspecified misadventure during medical care
C0418593|ICD9CM|AB|E876.9|Medical misadventure NOS
C0418624|ICD9CM|PT|E873.6|Nonadministration of necessary drug or medicinal substance
C0418624|ICD9CM|AB|E873.6|Nonadmin necess medicine
C0418626|ICD9CM|PT|E873.5|Inappropriate [too hot or too cold] temperature in local application and packing
C0418626|ICD9CM|AB|E873.5|Wrng temp in applic/pack
C0418696|ICD9CM|PT|E878.4|Other restorative surgery causing abnormal patient reaction, or later complication, without mention of misadventure at time of operation
C0418696|ICD9CM|AB|E878.4|Abn react-plast surg NEC
C0418697|ICD9CM|PT|E878.5|Amputation of limb(s) causing abnormal patient reaction, or later complication, without mention of misadventure at time of operation
C0418697|ICD9CM|AB|E878.5|Abn react-limb amputat
C0418710|ICD9CM|HT|E996|Injury due to war operations by nuclear weapons
C0418717|ICD9CM|AB|E993.9|War inj:explosion NOS
C0418717|ICD9CM|PT|E993.9|Injury due to war operations by unspecified explosion
C0418930|ICD9CM|PT|93.76|Training in use of lead dog for the blind
C0418930|ICD9CM|AB|93.76|Training in lead dog use
C0419069|ICD9CM|PT|99.11|Injection of Rh immune globulin
C0419069|ICD9CM|AB|99.11|Inject rh immune globul
C0419270|ICD9CM|PT|95.32|Prescription, fitting, and dispensing of contact lens
C0419270|ICD9CM|AB|95.32|Perscr/fit/disp contacts
C0419377|ICD9CM|PT|V27.4|Outcome of delivery, twins, both stillborn
C0419377|ICD9CM|AB|V27.4|Deliver-twins, both sb
C0419585|ICD9CM|PT|V73.3|Screening examination for rubella
C0419585|ICD9CM|AB|V73.3|Screening for rubella
C0420007|ICD9CM|AB|V74.2|Screening for leprosy
C0420007|ICD9CM|PT|V74.2|Screening examination for leprosy (Hansen's disease)
C0420015|ICD9CM|AB|V75.2|Screen for leishmaniasis
C0420015|ICD9CM|PT|V75.2|Screening examination for leishmaniasis
C0420019|ICD9CM|PT|V76.89|Special screening for other malignant neoplasms
C0420019|ICD9CM|AB|V76.89|Screen neoplasm NEC
C0420201|ICD9CM|PT|89.62|Central venous pressure monitoring
C0420201|ICD9CM|AB|89.62|Cvp monitoring
C0420585|ICD9CM|PT|V63.1|Medical services in home not available
C0420585|ICD9CM|AB|V63.1|No medical serv in home
C0423124|ICD9CM|AB|374.87|Dermatochalasis
C0423124|ICD9CM|PT|374.87|Dermatochalasis
C0423665|ICD9CM|AB|719.44|Joint pain-hand
C0423665|ICD9CM|PT|719.44|Pain in joint, hand
C0423729|ICD9CM|AB|786.52|Painful respiration
C0423729|ICD9CM|PT|786.52|Painful respiration
C0424000|ICD9CM|AB|V62.84|Suicidal ideation
C0424000|ICD9CM|PT|V62.84|Suicidal ideation
C0424605|ICD9CM|PT|315.9|Unspecified delay in development
C0424605|ICD9CM|AB|315.9|Development delay NOS
C0424641|ICD9CM|AB|781.91|Loss of height
C0424641|ICD9CM|PT|781.91|Loss of height
C0424813|ICD9CM|PT|376.33|Orbital edema or congestion
C0424813|ICD9CM|AB|376.33|Orbital edema
C0426066|ICD9CM|HT|652.0|Unstable lie of fetus
C0426187|ICD9CM|HT|652.5|High fetal head at term
C0426365|ICD9CM|PT|788.65|Straining on urination
C0426365|ICD9CM|AB|788.65|Straining on urination
C0426636|ICD9CM|PT|787.63|Fecal urgency
C0426636|ICD9CM|AB|787.63|Fecal urgency
C0427055|ICD9CM|AB|438.83|Facial weakness
C0427055|ICD9CM|AB|781.94|Facial weakness
C0427055|ICD9CM|PT|781.94|Facial weakness
C0427055|ICD9CM|PT|438.83|Other late effects of cerebrovascular disease, facial weakness
C0428908|ICD9CM|PT|427.81|Sinoatrial node dysfunction
C0428908|ICD9CM|AB|427.81|Sinoatrial node dysfunct
C0430458|ICD9CM|PT|89.41|Cardiovascular stress test using treadmill
C0430458|ICD9CM|AB|89.41|Treadmill stress test
C0430459|ICD9CM|PT|89.43|Cardiovascular stress test using bicycle ergometer
C0430459|ICD9CM|AB|89.43|Bicycle ergometer test
C0430520|ICD9CM|PT|89.42|Masters' two-step stress test
C0430520|ICD9CM|AB|89.42|Masters' 2-step test
C0431319|ICD9CM|PT|741.03|Spina bifida with hydrocephalus, lumbar region
C0431319|ICD9CM|AB|741.03|Spin bif w hydrceph-lumb
C0431320|ICD9CM|PT|741.02|Spina bifida with hydrocephalus, dorsal (thoracic) region
C0431320|ICD9CM|AB|741.02|Spin bif w hydrceph-dors
C0431321|ICD9CM|PT|741.01|Spina bifida with hydrocephalus, cervical region
C0431321|ICD9CM|AB|741.01|Spin bif w hydrceph-cerv
C0431467|ICD9CM|PT|744.02|Other anomalies of external ear with impairment of hearing
C0431467|ICD9CM|AB|744.02|Ex ear anm NEC-impr hear
C0431468|ICD9CM|AB|744.03|Middle ear anomaly NEC
C0431468|ICD9CM|PT|744.03|Anomaly of middle ear, except ossicles
C0431479|ICD9CM|PT|744.29|Other specified anomalies of ear
C0431479|ICD9CM|AB|744.29|Ear anomalies NEC
C0431491|ICD9CM|PT|744.49|Other branchial cleft cyst or fistula; preauricular sinus
C0431491|ICD9CM|AB|744.49|Branchial cleft anom NEC
C0431510|ICD9CM|PT|748.3|Other anomalies of larynx, trachea, and bronchus
C0431510|ICD9CM|AB|748.3|Laryngotrach anomaly NEC
C0431553|ICD9CM|HT|750.2|Other specified congenital anomalies of mouth and pharynx
C0431614|ICD9CM|PT|752.89|Other specified anomalies of genital organs
C0431614|ICD9CM|HT|752.8|Other specified congenital anomalies of genital organs
C0431614|ICD9CM|AB|752.89|Genital organ anom NEC
C0431635|ICD9CM|PT|752.39|Other anomalies of uterus
C0431635|ICD9CM|HT|752.3|Other congenital anomalies of uterus
C0431635|ICD9CM|AB|752.39|Anomalies of uterus NEC
C0431668|ICD9CM|AB|752.65|Hidden penis
C0431668|ICD9CM|PT|752.65|Hidden penis
C0431681|ICD9CM|HT|753.2|Obstructive defects of renal pelvis and ureter, congenital
C0431681|ICD9CM|PT|753.20|Unspecified obstructive defect of renal pelvis and ureter
C0431681|ICD9CM|AB|753.20|Obs dfct ren plv&urt NOS
C0431705|ICD9CM|PT|753.19|Other specified cystic kidney disease
C0431705|ICD9CM|AB|753.19|Cystic kidney diseas NEC
C0431725|ICD9CM|PT|753.4|Other specified anomalies of ureter
C0431725|ICD9CM|AB|753.4|Ureteral anomaly NEC
C0431741|ICD9CM|AB|753.7|Anomalies of urachus
C0431741|ICD9CM|PT|753.7|Anomalies of urachus
C0431826|ICD9CM|PT|755.21|Transverse deficiency of upper limb
C0431826|ICD9CM|AB|755.21|Transverse defic arm
C0431943|ICD9CM|PT|755.60|Unspecified anomaly of lower limb
C0431943|ICD9CM|AB|755.60|Lower limb anomaly NOS
C0431946|ICD9CM|HT|754.4|Congenital genu recurvatum and bowing of long bones of leg
C0432018|ICD9CM|PT|755.66|Other anomalies of toes
C0432018|ICD9CM|AB|755.66|Anomalies of toes NEC
C0432068|ICD9CM|PT|754.0|Congenital musculoskeletal deformities of skull, face, and jaw
C0432068|ICD9CM|AB|754.0|Cong skull/face/jaw def
C0432133|ICD9CM|PT|756.3|Other anomalies of ribs and sternum
C0432133|ICD9CM|AB|756.3|Rib & sternum anomal NEC
C0432138|ICD9CM|PT|756.19|Other anomalies of spine
C0432138|ICD9CM|AB|756.19|Anomaly of spine NEC
C0432162|ICD9CM|PT|756.11|Spondylolysis, lumbosacral region
C0432162|ICD9CM|AB|756.11|Lumbosacr spondylolysis
C0432333|ICD9CM|AB|757.2|Dermatoglyphic anomalies
C0432333|ICD9CM|PT|757.2|Dermatoglyphic anomalies
C0432340|ICD9CM|PT|757.4|Specified anomalies of hair
C0432340|ICD9CM|AB|757.4|Hair anomalies NEC
C0432351|ICD9CM|PT|757.5|Specified anomalies of nails
C0432351|ICD9CM|AB|757.5|Nail anomalies NEC
C0432354|ICD9CM|PT|757.6|Specified congenital anomalies of breast
C0432354|ICD9CM|AB|757.6|Cong breast anomaly NEC
C0432378|ICD9CM|PT|759.2|Anomalies of other endocrine glands
C0432378|ICD9CM|AB|759.2|Endocrine anomaly NEC
C0432487|ICD9CM|PT|238.77|Post-transplant lymphoproliferative disorder (PTLD)
C0432487|ICD9CM|AB|238.77|Post tp lymphprolif dis
C0432520|ICD9CM|PT|140.1|Malignant neoplasm of lower lip, vermilion border
C0432520|ICD9CM|AB|140.1|Mal neo lower vermilion
C0432534|ICD9CM|PT|201.08|Hodgkin's paragranuloma, lymph nodes of multiple sites
C0432534|ICD9CM|AB|201.08|Hodgkins paragran mult
C0432538|ICD9CM|PT|202.31|Malignant histiocytosis, lymph nodes of head, face, and neck
C0432538|ICD9CM|AB|202.31|Mal histiocytosis head
C0432539|ICD9CM|PT|202.32|Malignant histiocytosis, intrathoracic lymph nodes
C0432539|ICD9CM|AB|202.32|Mal histiocytosis thorax
C0432540|ICD9CM|PT|202.33|Malignant histiocytosis, intra-abdominal lymph nodes
C0432540|ICD9CM|AB|202.33|Mal histiocytosis abdom
C0432541|ICD9CM|PT|202.34|Malignant histiocytosis, lymph nodes of axilla and upper limb
C0432541|ICD9CM|AB|202.34|Mal histiocytosis axilla
C0432542|ICD9CM|PT|202.35|Malignant histiocytosis, lymph nodes of inguinal region and lower limb
C0432542|ICD9CM|AB|202.35|Mal histiocytosis inguin
C0432543|ICD9CM|PT|202.36|Malignant histiocytosis, intrapelvic lymph nodes
C0432543|ICD9CM|AB|202.36|Mal histiocytosis pelvic
C0432544|ICD9CM|PT|202.37|Malignant histiocytosis, spleen
C0432544|ICD9CM|AB|202.37|Mal histiocytosis spleen
C0432545|ICD9CM|PT|202.38|Malignant histiocytosis, lymph nodes of multiple sites
C0432545|ICD9CM|AB|202.38|Mal histiocytosis mult
C0432547|ICD9CM|PT|202.51|Letterer-siwe disease, lymph nodes of head, face, and neck
C0432547|ICD9CM|AB|202.51|Letterer-siwe dis head
C0432548|ICD9CM|PT|202.52|Letterer-siwe disease, intrathoracic lymph nodes
C0432548|ICD9CM|AB|202.52|Letterer-siwe dis thorax
C0432549|ICD9CM|PT|202.53|Letterer-siwe disease, intra-abdominal lymph nodes
C0432549|ICD9CM|AB|202.53|Letterer-siwe dis abdom
C0432550|ICD9CM|PT|202.54|Letterer-siwe disease, lymph nodes of axilla and upper limb
C0432550|ICD9CM|AB|202.54|Letterer-siwe dis axilla
C0432551|ICD9CM|PT|202.55|Letterer-siwe disease, lymph nodes of inguinal region and lower limb
C0432551|ICD9CM|AB|202.55|Letterer-siwe dis inguin
C0432552|ICD9CM|PT|202.56|Letterer-siwe disease, intrapelvic lymph nodes
C0432552|ICD9CM|AB|202.56|Letterer-siwe dis pelvic
C0432553|ICD9CM|PT|202.57|Letterer-siwe disease, spleen
C0432553|ICD9CM|AB|202.57|Letterer-siwe dis spleen
C0432554|ICD9CM|PT|202.58|Letterer-siwe disease, lymph nodes of multiple sites
C0432554|ICD9CM|AB|202.58|Letterer-siwe dis mult
C0432579|ICD9CM|PT|140.3|Malignant neoplasm of upper lip, inner aspect
C0432579|ICD9CM|AB|140.3|Mal neo upper lip, inner
C0432581|ICD9CM|PT|143.1|Malignant neoplasm of lower gum
C0432581|ICD9CM|AB|143.1|Malig neo lower gum
C0432721|ICD9CM|HT|914|Superficial injury of hand(s) except finger(s) alone
C0432762|ICD9CM|AB|923.10|Contusion of forearm
C0432762|ICD9CM|PT|923.10|Contusion of forearm
C0432763|ICD9CM|AB|923.11|Contusion of elbow
C0432763|ICD9CM|PT|923.11|Contusion of elbow
C0432769|ICD9CM|AB|923.20|Contusion of hand(s)
C0432769|ICD9CM|PT|923.20|Contusion of hand(s)
C0432773|ICD9CM|AB|923.3|Contusion of finger
C0432773|ICD9CM|PT|923.3|Contusion of finger
C0432869|ICD9CM|PT|917.0|Abrasion or friction burn of foot and toe(s), without mention of infection
C0432869|ICD9CM|AB|917.0|Abrasion foot & toe
C0432873|ICD9CM|PT|917.1|Abrasion or friction burn of foot and toe(s), infected
C0432873|ICD9CM|AB|917.1|Abrasion foot/toe-infec
C0432918|ICD9CM|PT|917.2|Blister of foot and toe(s), without mention of infection
C0432918|ICD9CM|AB|917.2|Blister foot & toe
C0432922|ICD9CM|PT|917.3|Blister of foot and toe(s), infected
C0432922|ICD9CM|AB|917.3|Blister foot & toe-infec
C0432959|ICD9CM|HT|880|Open wound of shoulder and upper arm
C0433039|ICD9CM|PT|917.4|Insect bite, nonvenomous, of foot and toe(s), without mention of infection
C0433039|ICD9CM|AB|917.4|Insect bite foot/toe
C0433050|ICD9CM|PT|917.5|Insect bite, nonvenomous, of foot and toe(s), infected
C0433050|ICD9CM|AB|917.5|Insect bite foot/toe-inf
C0433193|ICD9CM|HT|943|Burn of upper limb, except wrist and hand
C0433205|ICD9CM|HT|944|Burn of wrist(s) and hand(s)
C0433217|ICD9CM|PT|947.4|Burn of vagina and uterus
C0433217|ICD9CM|AB|947.4|Burn of vagina & uterus
C0433219|ICD9CM|HT|948|Burns classified according to extent of body surface involved
C0433307|ICD9CM|PT|941.14|Erythema [first degree] of chin
C0433307|ICD9CM|AB|941.14|1st deg burn chin
C0433333|ICD9CM|PT|944.16|Erythema [first degree] of back of hand
C0433333|ICD9CM|AB|944.16|1 deg burn back of hand
C0433353|ICD9CM|HT|942.2|Blisters with epidermal loss due to burn [second degree] of trunk
C0433361|ICD9CM|PT|944.20|Blisters, epidermal loss [second degree] of hand, unspecified site
C0433361|ICD9CM|AB|944.20|2nd deg burn hand NOS
C0433480|ICD9CM|PT|942.31|Full-thickness skin loss [third degree,not otherwise specified] of breast
C0433480|ICD9CM|AB|942.31|3rd deg burn breast
C0433482|ICD9CM|PT|942.33|Full-thickness skin loss [third degree, not otherwise specified] of abdominal wall
C0433482|ICD9CM|AB|942.33|3rd deg burn abdomn wall
C0433625|ICD9CM|PT|895.1|Traumatic amputation of toe(s) (complete) (partial), complicated
C0433625|ICD9CM|AB|895.1|Amputation toe-complicat
C0433638|ICD9CM|PT|885.0|Traumatic amputation of thumb (complete)(partial), without mention of complication
C0433638|ICD9CM|AB|885.0|Amputation thumb
C0433686|ICD9CM|PT|939.1|Foreign body in uterus, any part
C0433686|ICD9CM|AB|939.1|Foreign body uterus
C0433815|ICD9CM|PT|851.00|Cortex (cerebral) contusion without mention of open intracranial wound, unspecified state of consciousness
C0433815|ICD9CM|AB|851.00|Cerebral cortx contusion
C0433816|ICD9CM|PT|851.01|Cortex (cerebral) contusion without mention of open intracranial wound, with no loss of consciousness
C0433816|ICD9CM|AB|851.01|Cortex contusion-no coma
C0433821|ICD9CM|PT|851.06|Cortex (cerebral) contusion without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0433821|ICD9CM|AB|851.06|Cortex contus-coma NOS
C0433845|ICD9CM|PT|851.35|Cortex (cerebral) laceration with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0433845|ICD9CM|AB|851.35|Opn cortex lac-deep coma
C0433846|ICD9CM|HT|851.2|Cortex (cerebral) laceration without mention of open intracranial wound
C0433847|ICD9CM|PT|851.20|Cortex (cerebral) laceration without mention of open intracranial wound, unspecified state of consciousness
C0433847|ICD9CM|AB|851.20|Cerebral cortex lacerat
C0433848|ICD9CM|PT|851.21|Cortex (cerebral) laceration without mention of open intracranial wound, with no loss of consciousness
C0433848|ICD9CM|AB|851.21|Cortex lacerat w/o coma
C0433853|ICD9CM|PT|851.26|Cortex (cerebral) laceration without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0433853|ICD9CM|AB|851.26|Cortex lacerat-coma NOS
C0433854|ICD9CM|PT|851.29|Cortex (cerebral) laceration without mention of open intracranial wound, with concussion, unspecified
C0433854|ICD9CM|AB|851.29|Cortex lacerat-concuss
C0433857|ICD9CM|HT|954|Injury to other nerve(s) of trunk, excluding shoulder and pelvic girdles
C0433858|ICD9CM|HT|952.0|Cervical spinal cord injury without evidence of spinal bone injury
C0433976|ICD9CM|PT|871.0|Ocular laceration without prolapse of intraocular tissue
C0433976|ICD9CM|AB|871.0|Ocular lac w/o prolapse
C0433980|ICD9CM|PT|870.1|Laceration of eyelid, full-thickness, not involving lacrimal passages
C0433980|ICD9CM|AB|870.1|Full-thicknes lac eyelid
C0433981|ICD9CM|PT|870.2|Laceration of eyelid involving lacrimal passages
C0433981|ICD9CM|AB|870.2|Lac eyelid inv lacrm pas
C0434058|ICD9CM|PT|863.59|Other injury to colon or rectum, with open wound into cavity
C0434058|ICD9CM|AB|863.59|Colon injury NEC-open
C0434062|ICD9CM|PT|863.49|Other injury to colon or rectum, without mention of open wound into cavity
C0434062|ICD9CM|AB|863.49|Colon injury NEC-closed
C0434143|ICD9CM|PT|878.2|Open wound of scrotum and testes, without mention of complication
C0434143|ICD9CM|AB|878.2|Opn wound scrotum/testes
C0434195|ICD9CM|PT|903.1|Injury to brachial blood vessels
C0434195|ICD9CM|AB|903.1|Injury brachial vessels
C0434291|ICD9CM|PT|957.1|Injury to other specified nerve(s)
C0434291|ICD9CM|AB|957.1|Injury to nerve NEC
C0434322|ICD9CM|PT|840.4|Rotator cuff (capsule) sprain
C0434322|ICD9CM|AB|840.4|Sprain rotator cuff
C0434411|ICD9CM|HT|848.4|Sternum sprain
C0434411|ICD9CM|AB|848.40|Sprain of sternum NOS
C0434411|ICD9CM|PT|848.40|Sprain of sternum, unspecified site
C0434473|ICD9CM|PT|846.1|Sprain of sacroiliac ligament
C0434473|ICD9CM|AB|846.1|Sprain sacroiliac
C0434483|ICD9CM|AB|843.1|Sprain ischiocapsular
C0434483|ICD9CM|PT|843.1|Ischiocapsular (ligament) sprain
C0434579|ICD9CM|HT|831.0|Closed dislocation of shoulder
C0434583|ICD9CM|HT|831.1|Open dislocation of shoulder
C0434585|ICD9CM|PT|831.11|Open anterior dislocation of humerus
C0434585|ICD9CM|AB|831.11|Ant disloc humerus-open
C0434587|ICD9CM|PT|831.13|Open inferior dislocation of humerus
C0434587|ICD9CM|AB|831.13|Infer disloc humerus-opn
C0434599|ICD9CM|HT|832.0|Closed dislocation of elbow
C0434601|ICD9CM|PT|832.11|Open anterior dislocation of elbow
C0434601|ICD9CM|AB|832.11|Ant disloc elbow-open
C0434602|ICD9CM|PT|832.12|Open posterior dislocation of elbow
C0434602|ICD9CM|AB|832.12|Post disloc elbow-open
C0434603|ICD9CM|PT|832.13|Open medial dislocation of elbow
C0434603|ICD9CM|AB|832.13|Med disloc elbow-open
C0434604|ICD9CM|PT|832.14|Open lateral dislocation of elbow
C0434604|ICD9CM|AB|832.14|Lat dislocat elbow-open
C0434608|ICD9CM|HT|832.1|Open dislocation of elbow
C0434608|ICD9CM|PT|832.10|Open dislocation of elbow, unspecified
C0434608|ICD9CM|AB|832.10|Dislocat elbow NOS-open
C0434619|ICD9CM|HT|833.1|Open dislocation of wrist
C0434663|ICD9CM|PT|835.11|Open posterior dislocation of hip
C0434663|ICD9CM|AB|835.11|Posterior disloc hip-opn
C0434666|ICD9CM|HT|835.1|Open dislocation of hip
C0434685|ICD9CM|PT|836.3|Dislocation of patella, closed
C0434685|ICD9CM|AB|836.3|Dislocat patella-closed
C0434691|ICD9CM|HT|837|Dislocation of ankle
C0434692|ICD9CM|PT|837.0|Closed dislocation of ankle
C0434692|ICD9CM|AB|837.0|Dislocation ankle-closed
C0434696|ICD9CM|HT|838.0|Closed dislocation of foot
C0434707|ICD9CM|HT|838.1|Open dislocation of foot
C0434714|ICD9CM|PT|838.13|Open dislocation of tarsometatarsal (joint)
C0434714|ICD9CM|AB|838.13|Disl tarsometatarsal-opn
C0434715|ICD9CM|PT|838.12|Open dislocation of midtarsal (joint)
C0434715|ICD9CM|AB|838.12|Disloc midtarsal-open
C0434992|ICD9CM|PT|717.41|Bucket handle tear of lateral meniscus
C0434992|ICD9CM|AB|717.41|Old bucket tear lat men
C0435003|ICD9CM|AB|840.2|Sprain coracohumeral
C0435003|ICD9CM|PT|840.2|Coracohumeral (ligament) sprain
C0435005|ICD9CM|PT|841.3|Ulnohumeral (joint) sprain
C0435005|ICD9CM|AB|841.3|Sprain ulnohumeral
C0435018|ICD9CM|PT|844.3|Sprain of tibiofibular (joint) (ligament) superior, of knee
C0435018|ICD9CM|AB|844.3|Sprain super tibiofibula
C0435019|ICD9CM|PT|848.5|Sprain of pelvic
C0435019|ICD9CM|AB|848.5|Sprain of pelvis
C0435271|ICD9CM|HT|801.0|Closed fracture of base of skull without mention of intracranial injury
C0435334|ICD9CM|PT|802.25|Closed fracture of mandible, angle of jaw
C0435334|ICD9CM|AB|802.25|Fx angle of jaw-closed
C0435335|ICD9CM|PT|802.28|Closed fracture of mandible, body, other and unspecified
C0435335|ICD9CM|AB|802.28|Fx mandible body NEC-cl
C0435337|ICD9CM|PT|802.35|Open fracture of mandible, angle of jaw
C0435337|ICD9CM|AB|802.35|Fx angle of jaw-open
C0435338|ICD9CM|PT|802.38|Open fracture of mandible, body, other and unspecified
C0435338|ICD9CM|AB|802.38|Fx mandible body NEC-opn
C0435349|ICD9CM|HT|806|Fracture of vertebral column with spinal cord injury
C0435397|ICD9CM|PT|806.01|Closed fracture of C1-C4 level with complete lesion of cord
C0435397|ICD9CM|AB|806.01|C1-c4 fx-cl/com cord les
C0435403|ICD9CM|PT|806.06|Closed fracture of C5-C7 level with complete lesion of cord
C0435403|ICD9CM|AB|806.06|C5-c7 fx-cl/com cord les
C0435410|ICD9CM|PT|806.11|Open fracture of C1-C4 level with complete lesion of cord
C0435410|ICD9CM|AB|806.11|C1-c4 fx-op/com cord les
C0435416|ICD9CM|PT|806.16|Open fracture of C5-C7 level with complete lesion of cord
C0435416|ICD9CM|AB|806.16|C5-c7 fx-op/com cord les
C0435439|ICD9CM|PT|806.21|Closed fracture of T1-T6 level with complete lesion of cord
C0435439|ICD9CM|AB|806.21|T1-t6 fx-cl/com cord les
C0435445|ICD9CM|PT|806.26|Closed fracture of T7-T12 level with complete lesion of cord
C0435445|ICD9CM|AB|806.26|T7-t12 fx-cl/com crd les
C0435452|ICD9CM|PT|806.31|Open fracture of T1-T6 level with complete lesion of cord
C0435452|ICD9CM|AB|806.31|T1-t6 fx-op/com cord les
C0435457|ICD9CM|PT|806.36|Open fracture of T7-T12 level with complete lesion of cord
C0435457|ICD9CM|AB|806.36|T7-t12 fx-op/com crd les
C0435484|ICD9CM|PT|806.5|Open fracture of lumbar spine with spinal cord injury
C0435484|ICD9CM|AB|806.5|Opn lumbar fx w cord inj
C0435521|ICD9CM|PT|810.01|Closed fracture of sternal end of clavicle
C0435521|ICD9CM|AB|810.01|Fx clavicl, stern end-cl
C0435522|ICD9CM|PT|810.03|Closed fracture of acromial end of clavicle
C0435522|ICD9CM|AB|810.03|Fx clavicl, acrom end-cl
C0435523|ICD9CM|PT|810.11|Open fracture of sternal end of clavicle
C0435523|ICD9CM|AB|810.11|Fx clavic, stern end-opn
C0435524|ICD9CM|PT|810.13|Open fracture of acromial end of clavicle
C0435524|ICD9CM|AB|810.13|Fx clavic, acrom end-opn
C0435525|ICD9CM|PT|811.02|Closed fracture of coracoid process of scapula
C0435525|ICD9CM|AB|811.02|Fx scapul, corac proc-cl
C0435532|ICD9CM|PT|812.02|Closed fracture of anatomical neck of humerus
C0435532|ICD9CM|AB|812.02|Fx anatom nck humerus-cl
C0435533|ICD9CM|PT|812.03|Closed fracture of greater tuberosity of humerus
C0435533|ICD9CM|AB|812.03|Fx gr tuberos humerus-cl
C0435539|ICD9CM|PT|812.12|Open fracture of anatomical neck of humerus
C0435539|ICD9CM|AB|812.12|Fx anat neck humerus-opn
C0435540|ICD9CM|PT|812.13|Open fracture of greater tuberosity of humerus
C0435540|ICD9CM|AB|812.13|Fx gr tuberos humer-open
C0435552|ICD9CM|PT|812.42|Closed fracture of lateral condyle of humerus
C0435552|ICD9CM|AB|812.42|Fx humer, lat condyl-cl
C0435553|ICD9CM|PT|812.43|Closed fracture of medial condyle of humerus
C0435553|ICD9CM|AB|812.43|Fx humer, med condyl-cl
C0435563|ICD9CM|PT|812.52|Open fracture of lateral condyle of humerus
C0435563|ICD9CM|AB|812.52|Fx humer, lat condyl-opn
C0435564|ICD9CM|PT|812.53|Open fracture of medial condyle of humerus
C0435564|ICD9CM|AB|812.53|Fx humer, med condyl-opn
C0435569|ICD9CM|PT|812.41|Closed supracondylar fracture of humerus
C0435569|ICD9CM|AB|812.41|Suprcondyl fx humerus-cl
C0435570|ICD9CM|PT|812.51|Open supracondylar fracture of humerus
C0435570|ICD9CM|AB|812.51|Supracondyl fx humer-opn
C0435603|ICD9CM|PT|813.02|Closed fracture of coronoid process of ulna
C0435603|ICD9CM|AB|813.02|Fx coronoid proc ulna-cl
C0435623|ICD9CM|HT|813.0|Fracture of upper end of radius and ulna, closed
C0435623|ICD9CM|PT|813.08|Closed fracture of radius with ulna, upper end [any part]
C0435623|ICD9CM|AB|813.08|Fx up radius w ulna-clos
C0435633|ICD9CM|PT|814.02|Closed fracture of lunate [semilunar] bone of wrist
C0435633|ICD9CM|AB|814.02|Fx lunate, wrist-closed
C0435634|ICD9CM|PT|814.06|Closed fracture of trapezoid bone [smaller multangular] of wrist
C0435634|ICD9CM|AB|814.06|Fx trapezoid bone-closed
C0435638|ICD9CM|PT|814.12|Open fracture of lunate [semilunar] bone of wrist
C0435638|ICD9CM|AB|814.12|Fx lunate, wrist-open
C0435639|ICD9CM|PT|814.16|Open fracture of trapezoid bone [smaller multangular] of wrist
C0435639|ICD9CM|AB|814.16|Fx trapezoid bone-open
C0435644|ICD9CM|PT|814.01|Closed fracture of navicular [scaphoid] bone of wrist
C0435644|ICD9CM|AB|814.01|Fx navicular, wrist-clos
C0435650|ICD9CM|PT|814.11|Open fracture of navicular [scaphoid] bone of wrist
C0435650|ICD9CM|AB|814.11|Fx navicular, wrist-open
C0435656|ICD9CM|PT|815.19|Open fracture of multiple sites of metacarpus
C0435656|ICD9CM|AB|815.19|Mult fx metacarpus-open
C0435669|ICD9CM|PT|815.09|Closed fracture of multiple sites of metacarpus
C0435669|ICD9CM|AB|815.09|Mult fx metacarpus-close
C0435750|ICD9CM|HT|807.0|Closed fracture of rib(s)
C0435750|ICD9CM|AB|807.00|Fracture rib NOS-closed
C0435750|ICD9CM|PT|807.00|Closed fracture of rib(s), unspecified
C0435751|ICD9CM|HT|807.1|Open fracture of rib(s)
C0435751|ICD9CM|AB|807.10|Fracture rib NOS-open
C0435751|ICD9CM|PT|807.10|Open fracture of rib(s), unspecified
C0435771|ICD9CM|PT|808.51|Open fracture of ilium
C0435771|ICD9CM|AB|808.51|Fracture of ilium-open
C0435830|ICD9CM|PT|820.22|Closed fracture of subtrochanteric section of neck of femur
C0435830|ICD9CM|AB|820.22|Subtrochanteric fx-close
C0435834|ICD9CM|PT|820.32|Open fracture of subtrochanteric section of neck of femur
C0435834|ICD9CM|AB|820.32|Subtrochanteric fx-open
C0435844|ICD9CM|PT|821.23|Closed supracondylar fracture of femur
C0435844|ICD9CM|AB|821.23|Supracondyl fx femur-cl
C0435845|ICD9CM|PT|821.33|Open supracondylar fracture of femur
C0435845|ICD9CM|AB|821.33|Supracondyl fx femur-opn
C0435876|ICD9CM|PT|823.11|Open fracture of upper end of fibula alone
C0435876|ICD9CM|AB|823.11|Fx upper end fibula-open
C0435890|ICD9CM|PT|824.0|Fracture of medial malleolus, closed
C0435890|ICD9CM|AB|824.0|Fx medial malleolus-clos
C0435891|ICD9CM|PT|824.1|Fracture of medial malleolus, open
C0435891|ICD9CM|AB|824.1|Fx medial malleolus-open
C0435892|ICD9CM|PT|824.2|Fracture of lateral malleolus, closed
C0435892|ICD9CM|AB|824.2|Fx lateral malleolus-cl
C0435898|ICD9CM|PT|823.01|Closed fracture of upper end of fibula alone
C0435898|ICD9CM|AB|823.01|Fx upper end fibula-clos
C0435900|ICD9CM|PT|824.3|Fracture of lateral malleolus, open
C0435900|ICD9CM|AB|824.3|Fx lateral malleolus-opn
C0435903|ICD9CM|HT|823.0|Fracture of upper end of tibia and fibula, closed
C0435903|ICD9CM|PT|823.02|Closed fracture of upper end of fibula with tibia
C0435903|ICD9CM|AB|823.02|Fx up tibia w fibula-cl
C0435905|ICD9CM|HT|823.1|Fracture of upper end of tibia and fibula, open
C0435905|ICD9CM|PT|823.12|Open fracture of upper end of fibula with tibia
C0435905|ICD9CM|AB|823.12|Fx up tibia w fibula-opn
C0435920|ICD9CM|PT|825.34|Open fracture of cuneiform, foot
C0435920|ICD9CM|AB|825.34|Fx cuneiform, foot-open
C0435924|ICD9CM|PT|825.24|Closed fracture of cuneiform, foot
C0435924|ICD9CM|AB|825.24|Fx cuneiform, foot-clos
C0435940|ICD9CM|PT|825.22|Closed fracture of navicular [scaphoid], foot
C0435940|ICD9CM|AB|825.22|Fx navicular, foot-clos
C0435941|ICD9CM|PT|825.32|Open fracture of navicular [scaphoid], foot
C0435941|ICD9CM|AB|825.32|Fx navicular, foot-open
C0435944|ICD9CM|PT|825.25|Closed fracture of metatarsal bone(s)
C0435944|ICD9CM|AB|825.25|Fx metatarsal-closed
C0435950|ICD9CM|PT|825.35|Open fracture of metatarsal bone(s)
C0435950|ICD9CM|AB|825.35|Fx metatarsal-open
C0436055|ICD9CM|PT|959.11|Other injury of chest wall
C0436055|ICD9CM|AB|959.11|Injury of chest wall NEC
C0436064|ICD9CM|PT|959.14|Other injury of external genitals
C0436064|ICD9CM|AB|959.14|Inj external genital NEC
C0436099|ICD9CM|PT|905.2|Late effect of fracture of upper extremities
C0436099|ICD9CM|AB|905.2|Late effect arm fx
C0436114|ICD9CM|PT|909.1|Late effect of toxic effects of nonmedical substances
C0436114|ICD9CM|AB|909.1|Late eff nonmed substanc
C0436115|ICD9CM|HT|909|Late effects of other and unspecified external causes
C0438413|ICD9CM|PT|194.6|Malignant neoplasm of aortic body and other paraganglia
C0438413|ICD9CM|AB|194.6|Mal neo paraganglia NEC
C0438624|ICD9CM|AB|921.9|Contusion of eye NOS
C0438624|ICD9CM|PT|921.9|Unspecified contusion of eye
C0438699|ICD9CM|AB|748.5|Agenesis of lung
C0438699|ICD9CM|PT|748.5|Agenesis, hypoplasia, and dysplasia of lung
C0438989|ICD9CM|AB|V41.2|Problems with hearing
C0438989|ICD9CM|PT|V41.2|Problems with hearing
C0439001|ICD9CM|HT|743.5|Congenital anomalies of posterior segment
C0439002|ICD9CM|PT|756.81|Absence of muscle and tendon
C0439002|ICD9CM|AB|756.81|Absence of muscle/tendon
C0441655|ICD9CM|HT|E001-E030.9|ACTIVITY
C0451636|ICD9CM|PT|V22.2|Pregnant state, incidental
C0451636|ICD9CM|AB|V22.2|Preg state, incidental
C0451639|ICD9CM|HT|289|Other diseases of blood and blood-forming organs
C0451640|ICD9CM|PT|732.8|Other specified forms of osteochondropathy
C0451640|ICD9CM|AB|732.8|Osteochondropathy NEC
C0451984|ICD9CM|HT|929|Crushing injury of multiple and unspecified sites
C0451998|ICD9CM|PT|692.76|Sunburn of second degree
C0451998|ICD9CM|AB|692.76|2nd degree sunburn
C0452001|ICD9CM|PT|692.77|Sunburn of third degree
C0452001|ICD9CM|AB|692.77|3rd degree sunburn
C0452136|ICD9CM|PT|389.06|Conductive hearing loss, bilateral
C0452136|ICD9CM|AB|389.06|Condctv hear loss, bilat
C0452138|ICD9CM|PT|389.18|Sensorineural hearing loss, bilateral
C0452138|ICD9CM|AB|389.18|Sensonrl hear loss,bilat
C0452153|ICD9CM|PT|389.22|Mixed hearing loss, bilateral
C0452153|ICD9CM|AB|389.22|Mixed hearing loss,bilat
C0452240|ICD9CM|HT|93.1|Physical therapy exercises
C0454060|ICD9CM|AB|92.21|Superficial radiation
C0454060|ICD9CM|PT|92.21|Superficial radiation
C0454077|ICD9CM|PT|92.25|Teleradiotherapy using electrons
C0454077|ICD9CM|AB|92.25|Electron teleradiotherap
C0454533|ICD9CM|PT|438.14|Late effects of cerebrovascular disease, fluency disorder
C0454533|ICD9CM|AB|438.14|Late eff CV-fluency dis
C0455204|ICD9CM|AB|V62.85|Homicidal ideation
C0455204|ICD9CM|PT|V62.85|Homicidal ideation
C0455397|ICD9CM|PT|V19.11|Family history of glaucoma
C0455397|ICD9CM|AB|V19.11|Family history glaucoma
C0455422|ICD9CM|PT|V18.61|Family history of polycystic kidney
C0455422|ICD9CM|AB|V18.61|Fam hx-polycystic kidney
C0455701|ICD9CM|PT|V73.6|Screening examination for trachoma
C0455701|ICD9CM|AB|V73.6|Screening for trachoma
C0455970|ICD9CM|AB|63.71|Ligation of vas deferens
C0455970|ICD9CM|PT|63.71|Ligation of vas deferens
C0455988|ICD9CM|PT|778.0|Hydrops fetalis not due to isoimmunization
C0455988|ICD9CM|AB|778.0|Hydrops fetalis no isoim
C0455990|ICD9CM|PT|773.3|Hydrops fetalis due to isoimmunization
C0455990|ICD9CM|AB|773.3|Hydrops fetalis:isoimm
C0456017|ICD9CM|PT|770.7|Chronic respiratory disease arising in the perinatal period
C0456017|ICD9CM|AB|770.7|Perinatal chr resp dis
C0456089|ICD9CM|PT|768.6|Mild or moderate birth asphyxia
C0456089|ICD9CM|AB|768.6|Mild/mod birth asphyxia
C0456582|ICD9CM|PT|96.53|Irrigation of nasal passages
C0456582|ICD9CM|AB|96.53|Irrigation of nasal pass
C0472692|ICD9CM|PT|457.0|Postmastectomy lymphedema syndrome
C0472692|ICD9CM|AB|457.0|Postmastect lymphedema
C0472702|ICD9CM|HT|285|Other and unspecified anemias
C0472777|ICD9CM|AB|282.47|Hgb E-beta thalassemia
C0472777|ICD9CM|PT|282.47|Hemoglobin E-beta thalassemia
C0472948|ICD9CM|PT|42.01|Incision of esophageal web
C0472948|ICD9CM|AB|42.01|Esophageal web incision
C0473237|ICD9CM|PT|599.71|Gross hematuria
C0473237|ICD9CM|AB|599.71|Gross hematuria
C0473333|ICD9CM|AB|647.14|Gonorrhea-postpartum
C0473333|ICD9CM|PT|647.14|Gonorrhea of mother, complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication
C0473384|ICD9CM|PT|646.12|Edema or excessive weight gain in pregnancy, without mention of hypertension, delivered, with mention of postpartum complication
C0473384|ICD9CM|AB|646.12|Edema in preg-del w p/p
C0473388|ICD9CM|HT|644.1|Other threatened labor
C0473390|ICD9CM|HT|644.0|Threatened premature labor
C0473461|ICD9CM|AB|661.91|Abnormal labor NOS-deliv
C0473461|ICD9CM|PT|661.91|Unspecified abnormality of labor, delivered, with or without mention of antepartum condition
C0473462|ICD9CM|HT|661|Abnormality of forces of labor
C0473472|ICD9CM|HT|661.3|Precipitate labor
C0473485|ICD9CM|HT|669.0|Maternal distress
C0473508|ICD9CM|HT|666.2|Delayed and secondary postpartum hemorrhage
C0473508|ICD9CM|PT|666.20|Delayed and secondary postpartum hemorrhage, unspecified as to episode of care or not applicable
C0473508|ICD9CM|AB|666.24|Delay p/part hem-postpar
C0473508|ICD9CM|AB|666.20|Delay p/part hem-unspec
C0473508|ICD9CM|PT|666.24|Delayed and secondary postpartum hemorrhage, postpartum condition or complication
C0473719|ICD9CM|PT|719.18|Hemarthrosis, other specified sites
C0473719|ICD9CM|AB|719.18|Hemarthrosis-jt NEC
C0473748|ICD9CM|PT|715.15|Osteoarthrosis, localized, primary, pelvic region and thigh
C0473748|ICD9CM|AB|715.15|Loc prim osteoart-pelvis
C0473754|ICD9CM|HT|715.2|Osteoarthrosis, localized, secondary
C0473789|ICD9CM|PT|772.3|Umbilical hemorrhage after birth
C0473789|ICD9CM|AB|772.3|Post-birth umbil hemorr
C0473800|ICD9CM|HT|772|Fetal and neonatal hemorrhage
C0473833|ICD9CM|HT|763|Fetus or newborn affected by other complications of labor and delivery
C0473867|ICD9CM|PT|761.7|Malpresentation before labor affecting fetus or newborn
C0473867|ICD9CM|AB|761.7|Antepart malpres aff NB
C0473878|ICD9CM|PT|123.0|Taenia solium infection, intestinal form
C0473878|ICD9CM|AB|123.0|Taenia solium intestine
C0473975|ICD9CM|PT|968.2|Poisoning by other gaseous anesthetics
C0473975|ICD9CM|AB|968.2|Poison-gas anesthet NEC
C0474019|ICD9CM|PT|E938.5|Surface and infiltration anesthetics causing adverse effects in therapeutic use
C0474019|ICD9CM|AB|E938.5|Adv eff topic/infil anes
C0474035|ICD9CM|PT|E943.5|Antidiarrheal drugs causing adverse effects in therapeutic use
C0474035|ICD9CM|AB|E943.5|Adv eff antidiarrhea agt
C0474334|ICD9CM|PT|362.85|Retinal nerve fiber bundle defects
C0474334|ICD9CM|AB|362.85|Retinal nerv fiber defec
C0474442|ICD9CM|PT|371.24|Corneal edema due to wearing of contact lenses
C0474442|ICD9CM|AB|371.24|Edema d/t contact lens
C0474873|ICD9CM|AB|753.23|Congenital ureterocele
C0474873|ICD9CM|PT|753.23|Congenital ureterocele
C0474962|ICD9CM|PT|140.0|Malignant neoplasm of upper lip, vermilion border
C0474962|ICD9CM|AB|140.0|Mal neo upper vermilion
C0474963|ICD9CM|PT|141.5|Malignant neoplasm of junctional zone of tongue
C0474963|ICD9CM|AB|141.5|Mal neo tongue junction
C0474971|ICD9CM|PT|140.5|Malignant neoplasm of lip, unspecified, inner aspect
C0474971|ICD9CM|AB|140.5|Mal neo lip, inner NOS
C0475036|ICD9CM|PT|853.09|Other and unspecified intracranial hemorrhage following injury without mention of open intracranial wound, with concussion, unspecified
C0475036|ICD9CM|AB|853.09|Brain hem NEC-concussion
C0475045|ICD9CM|PT|853.19|Other and unspecified intracranial hemorrhage following injury with open intracranial wound, with concussion, unspecified
C0475045|ICD9CM|AB|853.19|Brain hem opn-concussion
C0475534|ICD9CM|PT|285.22|Anemia in neoplastic disease
C0475534|ICD9CM|AB|285.22|Anemia in neoplastic dis
C0475686|ICD9CM|PT|V10.60|Personal history of leukemia, unspecified
C0475686|ICD9CM|AB|V10.60|Hx of leukemia NOS
C0475713|ICD9CM|PT|770.3|Pulmonary hemorrhage
C0475713|ICD9CM|AB|770.3|NB pulmonary hemorrhage
C0476206|ICD9CM|AB|780.4|Dizziness and giddiness
C0476206|ICD9CM|PT|780.4|Dizziness and giddiness
C0476228|ICD9CM|PT|782.2|Localized superficial swelling, mass, or lump
C0476228|ICD9CM|AB|782.2|Local suprficial swellng
C0476232|ICD9CM|AB|782.4|Jaundice NOS
C0476232|ICD9CM|PT|782.4|Jaundice, unspecified, not of newborn
C0476235|ICD9CM|HT|783|Symptoms concerning nutrition, metabolism, and development
C0476241|ICD9CM|AB|783.42|Delayed milestones
C0476241|ICD9CM|PT|783.42|Delayed milestones
C0476247|ICD9CM|HT|784|Symptoms involving head and neck
C0476271|ICD9CM|HT|786|Symptoms involving respiratory system and other chest symptoms
C0476293|ICD9CM|HT|788|Symptoms involving urinary system
C0476310|ICD9CM|HT|789.3|Abdominal or pelvic swelling, mass, or lump
C0476319|ICD9CM|HT|790|Nonspecific findings on examination of blood
C0476338|ICD9CM|HT|791|Nonspecific findings on examination of urine
C0476346|ICD9CM|PT|792.1|Nonspecific abnormal findings in stool contents
C0476346|ICD9CM|AB|792.1|Abn find-stool contents
C0476359|ICD9CM|PT|793.0|Nonspecific (abnormal) findings on radiological and other examination of skull and head
C0476359|ICD9CM|AB|793.0|Nonsp abn fd-skull/head
C0476365|ICD9CM|HT|793.1|Nonspecific abnormal findings on radiological and other examination of lung field
C0476376|ICD9CM|PT|793.5|Nonspecific (abnormal) findings on radiological and other examination of genitourinary organs
C0476376|ICD9CM|AB|793.5|Nonsp abn find-gu organs
C0476388|ICD9CM|HT|794|Nonspecific abnormal results of function studies
C0476389|ICD9CM|HT|794.0|Nonspecific abnormal results of function study of brain and central nervous system
C0476389|ICD9CM|PT|794.00|Abnormal function study of brain and central nervous system, unspecified
C0476389|ICD9CM|AB|794.00|Abn cns funct study NOS
C0476391|ICD9CM|PT|794.01|Nonspecific abnormal echoencephalogram
C0476391|ICD9CM|AB|794.01|Abnorm echoencephalogram
C0476396|ICD9CM|PT|794.11|Nonspecific abnormal retinal function studies
C0476396|ICD9CM|AB|794.11|Abn retinal funct study
C0476402|ICD9CM|PT|794.16|Nonspecific abnormal vestibular function studies
C0476402|ICD9CM|AB|794.16|Abn vestibular func stud
C0476403|ICD9CM|PT|794.17|Nonspecific abnormal electromyogram [EMG]
C0476403|ICD9CM|AB|794.17|Abnorm electromyogram
C0476405|ICD9CM|PT|794.2|Nonspecific abnormal results of pulmonary function study
C0476405|ICD9CM|AB|794.2|Abn pulmonary func study
C0476409|ICD9CM|HT|794.3|Nonspecific abnormal results of function study, cardiovascular
C0476409|ICD9CM|PT|794.30|Abnormal cardiovascular function study, unspecified
C0476409|ICD9CM|AB|794.30|Abn cardiovasc study NOS
C0476414|ICD9CM|PT|794.5|Nonspecific abnormal results of function study of thyroid
C0476414|ICD9CM|AB|794.5|Abn thyroid funct study
C0476431|ICD9CM|PT|795.2|Nonspecific abnormal findings on chromosomal analysis
C0476431|ICD9CM|AB|795.2|Abn chromosomal analysis
C0476454|ICD9CM|PT|796.3|Nonspecific low blood pressure reading
C0476454|ICD9CM|AB|796.3|Low blood press reading
C0476465|ICD9CM|PT|799.9|Other unknown and unspecified cause of morbidity and mortality
C0476465|ICD9CM|AB|799.9|Unkn cause morb/mort NEC
C0476475|ICD9CM|HT|705.2|Focal hyperhidrosis
C0476476|ICD9CM|PT|780.8|Generalized hyperhidrosis
C0476476|ICD9CM|AB|780.8|Generalizd hyperhidrosis
C0476478|ICD9CM|PT|799.25|Demoralization and apathy
C0476478|ICD9CM|AB|799.25|Demoralization & apathy
C0476550|ICD9CM|PT|V08|Asymptomatic human immunodeficiency virus [HIV] infection status
C0476550|ICD9CM|AB|V08|Asymp hiv infectn status
C0476555|ICD9CM|PT|V05.3|Need for prophylactic vaccination and inoculation against viral hepatitis
C0476555|ICD9CM|AB|V05.3|Need prphyl vc vrl hepat
C0476556|ICD9CM|PT|V05.2|Need for prophylactic vaccination and inoculation against leishmaniasis
C0476556|ICD9CM|AB|V05.2|Vaccin for leishmaniasis
C0476560|ICD9CM|AB|V61.41|Alcoholism in family
C0476560|ICD9CM|PT|V61.41|Alcoholism in family
C0476582|ICD9CM|AB|V46.3|Wheelchair dependence
C0476582|ICD9CM|PT|V46.3|Wheelchair dependence
C0476658|ICD9CM|HT|V58.1|Encounter for antineoplastic chemotherapy and immunotherapy
C0476664|ICD9CM|PT|V64.09|Vaccination not carried out for other reason
C0476664|ICD9CM|AB|V64.09|No vaccination NEC
C0476665|ICD9CM|PT|V64.00|Vaccination not carried out, unspecified reason
C0476665|ICD9CM|AB|V64.00|No vaccination NOS
C0476681|ICD9CM|PT|V65.44|Human immunodeficiency virus (HIV) counseling
C0476681|ICD9CM|AB|V65.44|Hiv counseling
C0476700|ICD9CM|HT|V45.7|Acquired absence of organ
C0476705|ICD9CM|PT|V45.73|Acquired absence of kidney
C0476705|ICD9CM|AB|V45.73|Acquired absence kidney
C0476706|ICD9CM|PT|V45.77|Acquired absence of organ, genital organs
C0476706|ICD9CM|AB|V45.77|Acq absnce genital organ
C0476707|ICD9CM|PT|V20.0|Health supervision of foundling
C0476707|ICD9CM|AB|V20.0|Foundling health care
C0477306|ICD9CM|PT|282.49|Other thalassemia
C0477306|ICD9CM|AB|282.49|Thalassemia NEC
C0477317|ICD9CM|PT|287.39|Other primary thrombocytopenia
C0477317|ICD9CM|AB|287.39|Prim thrombocytopen NEC
C0477318|ICD9CM|PT|288.8|Other specified disease of white blood cells
C0477318|ICD9CM|AB|288.8|Wbc disease NEC
C0477341|ICD9CM|HT|323.0|Encephalitis, myelitis, and encephalomyelitis in viral diseases classified elsewhere
C0477355|ICD9CM|PT|333.90|Unspecified extrapyramidal disease and abnormal movement disorder
C0477355|ICD9CM|AB|333.90|Extrapyramidal dis NOS
C0477373|ICD9CM|HT|346.8|Other forms of migraine
C0477374|ICD9CM|HT|339.8|Other specified headache syndromes
C0477458|ICD9CM|AB|389.8|Hearing loss NEC
C0477458|ICD9CM|PT|389.8|Other specified forms of hearing loss
C0477492|ICD9CM|PT|695.19|Other erythema multiforme
C0477492|ICD9CM|AB|695.19|Erythema multiforme NEC
C0477572|ICD9CM|PT|735.4|Other hammer toe (acquired)
C0477572|ICD9CM|AB|735.4|Other hammer toe
C0477573|ICD9CM|PT|735.8|Other acquired deformities of toe
C0477573|ICD9CM|AB|735.8|Acq deformity of toe NEC
C0477758|ICD9CM|PT|599.89|Other specified disorders of urinary tract
C0477758|ICD9CM|AB|599.89|Oth spcf dsdr urnry trct
C0477784|ICD9CM|PT|622.8|Other specified noninflammatory disorders of cervix
C0477784|ICD9CM|AB|622.8|Noninflam dis cervix NEC
C0477810|ICD9CM|HT|639|Complications following abortion or ectopic and molar pregnancies
C0477810|ICD9CM|PT|639.9|Unspecified complication following abortion or ectopic and molar pregnancy
C0477810|ICD9CM|AB|639.9|Postabortion compl NOS
C0477814|ICD9CM|PT|671.83|Other venous complications of pregnancy and the puerperium, antepartum condition or complication
C0477814|ICD9CM|AB|671.83|Venous compl NEC-antepar
C0477835|ICD9CM|HT|656.7|Other placental conditions affecting management of mother
C0477838|ICD9CM|HT|661.2|Other and unspecified uterine inertia
C0477838|ICD9CM|PT|661.20|Other and unspecified uterine inertia, unspecified as to episode of care or not applicable
C0477838|ICD9CM|AB|661.20|Uterine inertia NEC-unsp
C0477869|ICD9CM|PT|671.84|Other venous complications of pregnancy and the puerperium, postpartum condition or complication
C0477869|ICD9CM|AB|671.84|Venous compl NEC-postpar
C0477876|ICD9CM|HT|647.6|Other viral diseases complicating pregnancy, childbirth, or the puerperium
C0477887|ICD9CM|PT|762.2|Other and unspecified morphological and functional abnormalities of placenta affecting fetus or newborn
C0477887|ICD9CM|AB|762.2|Abn plac NEC/NOS aff NB
C0477888|ICD9CM|PT|762.5|Other compression of umbilical cord affecting fetus or newborn
C0477888|ICD9CM|AB|762.5|Oth umbil cord compress
C0477889|ICD9CM|PT|762.6|Other and unspecified conditions of umbilical cord affecting fetus or newborn
C0477889|ICD9CM|AB|762.6|Umbil cond NEC aff NB
C0477891|ICD9CM|PT|763.1|Other malpresentation, malposition, and disproportion during labor and delivery affecting fetus or newborn
C0477891|ICD9CM|AB|763.1|Malpos/dispro NEC aff NB
C0477897|ICD9CM|PT|766.1|Other "heavy-for-dates" infants
C0477897|ICD9CM|AB|766.1|Heavy-for-date infan NEC
C0477903|ICD9CM|PT|767.8|Other specified birth trauma
C0477903|ICD9CM|AB|767.8|Birth trauma NEC
C0477914|ICD9CM|AB|770.82|Other apnea of newborn
C0477914|ICD9CM|PT|770.82|Other apnea of newborn
C0477961|ICD9CM|PT|778.8|Other specified conditions involving the integument of fetus and newborn
C0477961|ICD9CM|AB|778.8|NB integument cond NEC
C0477972|ICD9CM|PT|742.4|Other specified congenital anomalies of brain
C0477972|ICD9CM|AB|742.4|Brain anomaly NEC
C0477973|ICD9CM|HT|741.0|Spina bifida with hydrocephalus
C0477973|ICD9CM|PT|741.00|Spina bifida with hydrocephalus, unspecified region
C0477973|ICD9CM|AB|741.00|Spin bif w hydroceph NOS
C0477975|ICD9CM|HT|742.5|Other specified congenital anomalies of spinal cord
C0477975|ICD9CM|PT|742.59|Other specified congenital anomalies of spinal cord
C0477975|ICD9CM|AB|742.59|Spinal cord anomaly NEC
C0477976|ICD9CM|PT|742.8|Other specified congenital anomalies of nervous system
C0477976|ICD9CM|AB|742.8|Nervous system anom NEC
C0477986|ICD9CM|PT|743.8|Other specified anomalies of eye
C0477986|ICD9CM|AB|743.8|Eye anomalies NEC
C0477990|ICD9CM|HT|744.2|Other specified congenital anomalies of ear
C0477992|ICD9CM|HT|744.8|Other specified congenital anomalies of face and neck
C0477992|ICD9CM|PT|744.89|Other specified congenital anomalies of face and neck
C0477992|ICD9CM|AB|744.89|Cong face/neck anom NEC
C0477996|ICD9CM|PT|746.09|Other congenital anomalies of pulmonary valve
C0477996|ICD9CM|AB|746.09|Pulmonary valve anom NEC
C0477999|ICD9CM|HT|746.8|Other specified congenital anomalies of heart
C0477999|ICD9CM|PT|746.89|Other specified congenital anomalies of heart
C0477999|ICD9CM|AB|746.89|Cong heart anomaly NEC
C0478000|ICD9CM|HT|747.2|Other congenital anomalies of aorta
C0478000|ICD9CM|PT|747.29|Other anomalies of aorta
C0478000|ICD9CM|AB|747.29|Cong anom of aorta NEC
C0478008|ICD9CM|HT|747.8|Other specified congenital anomalies of circulatory system
C0478008|ICD9CM|PT|747.89|Other specified anomalies of circulatory system
C0478008|ICD9CM|AB|747.89|Circulatory anomaly NEC
C0478013|ICD9CM|PT|747.9|Unspecified anomaly of circulatory system
C0478013|ICD9CM|AB|747.9|Circulatory anomaly NOS
C0478014|ICD9CM|PT|748.1|Other anomalies of nose
C0478014|ICD9CM|AB|748.1|Nose anomaly NEC
C0478018|ICD9CM|PT|748.69|Other congenital anomalies of lung
C0478018|ICD9CM|HT|748.6|Congenital other anomalies of lung
C0478018|ICD9CM|AB|748.69|Lung anomaly NEC
C0478019|ICD9CM|PT|748.8|Other specified anomalies of respiratory system
C0478019|ICD9CM|AB|748.8|Respiratory anomaly NEC
C0478024|ICD9CM|HT|750.1|Other congenital anomalies of tongue
C0478024|ICD9CM|PT|750.19|Other congenital anomalies of tongue
C0478024|ICD9CM|AB|750.19|Tongue anomaly NEC
C0478039|ICD9CM|PT|751.8|Other specified anomalies of digestive system
C0478039|ICD9CM|AB|751.8|Anom digestive syst NEC
C0478043|ICD9CM|PT|752.19|Other anomalies of fallopian tubes and broad ligaments
C0478043|ICD9CM|AB|752.19|Tubal/broad lig anom NEC
C0478056|ICD9CM|PT|753.29|Other obstructive defects of renal pelvis and ureter
C0478056|ICD9CM|AB|753.29|Obst def ren plv&urt NEC
C0478058|ICD9CM|PT|753.3|Other specified anomalies of kidney
C0478058|ICD9CM|AB|753.3|Kidney anomaly NEC
C0478070|ICD9CM|HT|755.5|Other congenital anomalies of upper limb, including shoulder girdle
C0478070|ICD9CM|PT|755.59|Other anomalies of upper limb, including shoulder girdle
C0478070|ICD9CM|AB|755.59|Upper limb anomaly NEC
C0478071|ICD9CM|HT|755.6|Other congenital anomalies of lower limb, including pelvic girdle
C0478071|ICD9CM|PT|755.69|Other anomalies of lower limb, including pelvic girdle
C0478071|ICD9CM|AB|755.69|Lower limb anomaly NEC
C0478080|ICD9CM|PT|756.9|Other and unspecified anomalies of musculoskeletal system
C0478080|ICD9CM|AB|756.9|Musculoskel anom NEC/NOS
C0478090|ICD9CM|PT|757.8|Other specified anomalies of the integument
C0478090|ICD9CM|AB|757.8|Oth integument anomalies
C0478095|ICD9CM|HT|759.8|Other specified anomalies
C0478095|ICD9CM|PT|759.89|Other specified congenital anomalies
C0478095|ICD9CM|AB|759.89|Specfied cong anomal NEC
C0478100|ICD9CM|PT|758.39|Other autosomal deletions
C0478100|ICD9CM|AB|758.39|Autosomal deletions NEC
C0478140|ICD9CM|PT|799.29|Other signs and symptoms involving emotional state
C0478140|ICD9CM|AB|799.29|Emotional state sym NEC
C0478144|ICD9CM|HT|784.5|Other speech disturbance
C0478145|ICD9CM|HT|784.6|Other symbolic dysfunction
C0478145|ICD9CM|PT|784.69|Other symbolic dysfunction
C0478145|ICD9CM|AB|784.69|Symbolic dysfunction NEC
C0478148|ICD9CM|PT|338.29|Other chronic pain
C0478148|ICD9CM|AB|338.29|Chronic pain NEC
C0478205|ICD9CM|HT|951|Injury to other cranial nerve(s)
C0478263|ICD9CM|HT|867|Injury to pelvic organs
C0478269|ICD9CM|PT|912.8|Other and unspecified superficial injury of shoulder and upper arm, without mention of infection
C0478269|ICD9CM|AB|912.8|Superf inj shldr/arm NEC
C0478347|ICD9CM|PT|897.4|Traumatic amputation of leg(s) (complete) (partial), unilateral, level not specified, without mention of complication
C0478347|ICD9CM|AB|897.4|Amputat leg, unilat NOS
C0478453|ICD9CM|PT|975.8|Poisoning by other and unspecified respiratory drugs
C0478453|ICD9CM|AB|975.8|Pois-respir drug NEC/NOS
C0478483|ICD9CM|AB|999.59|Other serum reaction
C0478483|ICD9CM|PT|999.59|Other serum reaction
C0478550|ICD9CM|PT|V03.89|Other specified vaccination
C0478550|ICD9CM|AB|V03.89|Nd other specf vacnation
C0478559|ICD9CM|HT|V26.8|Other specified procreative management
C0478576|ICD9CM|PT|V53.09|Fitting and adjustment of other devices related to nervous system and special senses
C0478576|ICD9CM|AB|V53.09|Adj nerv syst device NEC
C0478581|ICD9CM|PT|V56.8|Encounter for other dialysis
C0478581|ICD9CM|AB|V56.8|Dialysis encounter, NEC
C0478874|ICD9CM|PT|E884.9|Other accidental fall from one level to another
C0478874|ICD9CM|HT|E884|Other accidental falls from one level to another
C0478874|ICD9CM|AB|E884.9|Fall-1 level to oth NEC
C0479196|ICD9CM|AB|E906.1|Rat bite
C0479196|ICD9CM|PT|E906.1|Rat bite
C0480040|ICD9CM|PT|E854.1|Accidental poisoning by psychodysleptics [hallucinogens]
C0480040|ICD9CM|AB|E854.1|Acc poison-hallucinogens
C0480073|ICD9CM|PT|E860.9|Accidental poisoning by unspecified alcohol
C0480073|ICD9CM|AB|E860.9|Acc poison-alcohol NOS
C0480147|ICD9CM|PT|E903|Accident caused by travel and motion
C0480147|ICD9CM|AB|E903|Travel and motion
C0480620|ICD9CM|PT|E965.4|Assault by other and unspecified firearm
C0480620|ICD9CM|AB|E965.4|Assault-firearm NEC
C0480686|ICD9CM|PT|E968.1|Assault by pushing from a high place
C0480686|ICD9CM|AB|E968.1|Asslt-push from hi place
C0481115|ICD9CM|PT|E930.1|Antifungal antibiotics causing adverse effects in therapeutic use
C0481115|ICD9CM|AB|E930.1|Adv eff antifung antbiot
C0481138|ICD9CM|PT|E935.6|Antirheumatics [antiphlogistics] causing adverse effects in therapeutic use
C0481138|ICD9CM|AB|E935.6|Adv eff antirheumatics
C0481142|ICD9CM|HT|E936|Anticonvulsants and anti-Parkinsonism drugs causing adverse effects in therapeutic use
C0481147|ICD9CM|PT|E936.4|Anti-parkinsonism drugs causing adverse effects in therapeutic use
C0481147|ICD9CM|AB|E936.4|Adv eff anti-parkinson
C0481188|ICD9CM|PT|E942.2|Antilipemic and antiarteriosclerotic drugs causing adverse effects in therapeutic use
C0481188|ICD9CM|AB|E942.2|Adv eff antilipemics
C0481197|ICD9CM|PT|E944.2|Carbonic acid anhydrase inhibitors causing adverse effects in therapeutic use
C0481197|ICD9CM|AB|E944.2|Adv eff acetazolamide
C0481202|ICD9CM|PT|E945.2|Skeletal muscle relaxants causing adverse effects in therapeutic use
C0481202|ICD9CM|AB|E945.2|Adv eff skelet musc relx
C0481222|ICD9CM|PT|E870.0|Accidental cut, puncture, perforation or hemorrhage during surgical operation
C0481222|ICD9CM|AB|E870.0|Acc cut/hem in surgery
C0481232|ICD9CM|PT|E871.1|Foreign object left in body during infusion or transfusion
C0481232|ICD9CM|AB|E871.1|Postinfusion foreign bdy
C0481233|ICD9CM|PT|E871.2|Foreign object left in body during kidney dialysis or other perfusion
C0481233|ICD9CM|AB|E871.2|Postperfusion forgn body
C0481234|ICD9CM|PT|E871.3|Foreign object left in body during injection or vaccination
C0481234|ICD9CM|AB|E871.3|Postinjection forgn body
C0481235|ICD9CM|PT|E871.4|Foreign object left in body during endoscopic examination
C0481235|ICD9CM|AB|E871.4|Postendoscopy forgn body
C0481236|ICD9CM|PT|E871.6|Foreign object left in body during heart catheterization
C0481236|ICD9CM|AB|E871.6|FB post heart catheter
C0481237|ICD9CM|PT|E871.5|Foreign object left in body during aspiration of fluid or tissue, puncture, and catheterization
C0481237|ICD9CM|AB|E871.5|Postcatheter forgn body
C0481246|ICD9CM|PT|E873.0|Excessive amount of blood or other fluid during transfusion or infusion
C0481246|ICD9CM|AB|E873.0|Excess fluid in infusion
C0481247|ICD9CM|PT|E873.1|Incorrect dilution of fluid during infusion
C0481247|ICD9CM|AB|E873.1|Incor dilut infusn fluid
C0481248|ICD9CM|PT|E873.2|Overdose of radiation in therapy
C0481248|ICD9CM|AB|E873.2|Therap radiation overdos
C0481253|ICD9CM|PT|E875.0|Contaminated substance transfused or infused
C0481253|ICD9CM|AB|E875.0|Contaminated transfusion
C0481254|ICD9CM|PT|E875.1|Contaminated substance injected or used for vaccination
C0481254|ICD9CM|AB|E875.1|Contaminated injection
C0481259|ICD9CM|PT|E876.2|Failure in suture and ligature during surgical operation
C0481259|ICD9CM|AB|E876.2|Failure in suture
C0481263|ICD9CM|HT|E870-E876.9|MISADVENTURES TO PATIENTS DURING SURGICAL AND MEDICAL CARE
C0481350|ICD9CM|PT|E879.5|Insertion of gastric or duodenal sound as the cause of abnormal reaction of patient, or of later complication, without mention of misadventure of time of procedure
C0481350|ICD9CM|AB|E879.5|Abn react-gastric sound
C0481354|ICD9CM|PT|E929.0|Late effects of motor vehicle accident
C0481354|ICD9CM|AB|E929.0|Late eff motor vehic acc
C0481355|ICD9CM|PT|E929.1|Late effects of other transport accident
C0481355|ICD9CM|AB|E929.1|Late eff transport acc
C0481358|ICD9CM|PT|E959|Late effects of self-inflicted injury
C0481358|ICD9CM|AB|E959|Late eff of self-injury
C0481360|ICD9CM|PT|E989|Late effects of injury, undetermined whether accidentally or purposely inflicted
C0481360|ICD9CM|AB|E989|Late eff inj-undet circ
C0481367|ICD9CM|PT|E977|Late effects of injuries due to legal intervention
C0481367|ICD9CM|AB|E977|Late eff-legal intervent
C0481368|ICD9CM|PT|E999.0|Late effect of injury due to war operations
C0481368|ICD9CM|AB|E999.0|Late effect, war injury
C0481434|ICD9CM|PT|V02.2|Carrier or suspected carrier of amebiasis
C0481434|ICD9CM|AB|V02.2|Amebiasis carrier
C0481436|ICD9CM|PT|V02.7|Carrier or suspected carrier of gonorrhea
C0481436|ICD9CM|AB|V02.7|Gonorrhea carrier
C0481459|ICD9CM|PT|V27.2|Outcome of delivery, twins, both liveborn
C0481459|ICD9CM|AB|V27.2|Deliver-twins, both live
C0481466|ICD9CM|PT|V27.3|Outcome of delivery, twins, one liveborn and one stillborn
C0481466|ICD9CM|AB|V27.3|Del-twins, 1 nb, 1 sb
C0481487|ICD9CM|PT|V43.5|Bladder replaced by other means
C0481487|ICD9CM|AB|V43.5|Bladder replacement NEC
C0481496|ICD9CM|AB|V45.11|Renal dialysis status
C0481496|ICD9CM|PT|V45.11|Renal dialysis status
C0481514|ICD9CM|HT|V61.4|Health problems within family
C0481522|ICD9CM|PT|V66.3|Convalescence following psychotherapy and other treatment for mental disorder
C0481522|ICD9CM|AB|V66.3|Mental dis convalescence
C0481525|ICD9CM|PT|V67.4|Follow-up examination, following treatment of healed fracture
C0481525|ICD9CM|AB|V67.4|FU exam treatd healed fx
C0481551|ICD9CM|HT|V02|Carrier or suspected carrier of infectious diseases
C0481651|ICD9CM|PT|V23.49|Pregnancy with other poor obstetric history
C0481651|ICD9CM|AB|V23.49|Preg w poor obs hx NEC
C0481671|ICD9CM|PT|V27.7|Outcome of delivery, other multiple birth, all stillborn
C0481671|ICD9CM|AB|V27.7|Del-mult birth, all sb
C0481686|ICD9CM|PT|V30.2|Single liveborn, born outside hospital and not hospitalized
C0481686|ICD9CM|AB|V30.2|Single liveborn-nonhosp
C0481689|ICD9CM|HT|V31|Twin birth, mate liveborn
C0481706|ICD9CM|PT|V41.6|Problems with swallowing and mastication
C0481706|ICD9CM|AB|V41.6|Problem w swallowing
C0481749|ICD9CM|PT|V52.3|Fitting and adjustment of dental prosthetic device
C0481749|ICD9CM|AB|V52.3|Fitting dental prosthes
C0481768|ICD9CM|PT|V53.8|Fitting and adjustment of wheelchair
C0481768|ICD9CM|AB|V53.8|Adjustment of wheelchair
C0481797|ICD9CM|HT|V61|Other family circumstances
C0481798|ICD9CM|HT|V61.0|Family disruption
C0481799|ICD9CM|AB|V61.8|Family circumstances NEC
C0481799|ICD9CM|PT|V61.8|Other specified family circumstances
C0481845|ICD9CM|PT|V70.3|Other general medical examination for administrative purposes
C0481845|ICD9CM|AB|V70.3|Med exam NEC-admin purp
C0481850|ICD9CM|PT|V29.8|Observation for other specified suspected conditions
C0481850|ICD9CM|HT|V71.8|Observation and evaluation for other specified suspected conditions
C0481850|ICD9CM|PT|V71.89|Observation and evaluation for other specified suspected conditions
C0481850|ICD9CM|AB|V71.89|Observ-suspect cond NEC
C0481850|ICD9CM|AB|V29.8|NB obsrv oth suspct cond
C0481870|ICD9CM|PT|V75.3|Screening examination for trypanosomiasis
C0481870|ICD9CM|AB|V75.3|Screen-trypanosomiasis
C0481873|ICD9CM|PT|V76.0|Special screening for malignant neoplasms of respiratory organs
C0481873|ICD9CM|AB|V76.0|Screen mal neop-resp org
C0489951|ICD9CM|HT|008.4|Intestinal infection due to other specified bacteria
C0489951|ICD9CM|PT|008.49|Intestinal infection due to other organisms
C0489951|ICD9CM|AB|008.49|Bacterial enteritis NEC
C0489952|MTH|PN|NOCODE|Intestinal infection due to other organism, NEC in ICD9CM
C0489952|ICD9CM|AB|008.8|Viral enteritis NOS
C0489952|ICD9CM|PT|008.8|Intestinal infection due to other organism, not elsewhere classified
C0489954|ICD9CM|PT|070.9|Unspecified viral hepatitis without mention of hepatic coma
C0489954|ICD9CM|AB|070.9|Viral hepat NOS w/o coma
C0489955|ICD9CM|PT|242.10|Toxic uninodular goiter without mention of thyrotoxic crisis or storm
C0489955|ICD9CM|AB|242.10|Tox uninod goit no cris
C0489958|ICD9CM|AB|392.9|Rheumatic chorea NOS
C0489958|ICD9CM|PT|392.9|Rheumatic chorea without mention of heart involvement
C0489959|ICD9CM|AB|398.0|Rheumatic myocarditis
C0489959|ICD9CM|PT|398.0|Rheumatic myocarditis
C0489962|ICD9CM|PT|532.90|Duodenal ulcer, unspecified as acute or chronic, without hemorrhage or perforation, without mention of obstruction
C0489962|ICD9CM|AB|532.90|Duodenal ulcer NOS
C0489966|ICD9CM|PT|574.51|Calculus of bile duct without mention of cholecystitis, with obstruction
C0489966|ICD9CM|AB|574.51|Choledochlith NOS w obst
C0489967|ICD9CM|AB|596.52|Low bladder compliance
C0489967|ICD9CM|PT|596.52|Low bladder compliance
C0489969|ICD9CM|PT|719.98|Unspecified disorder of joint, other specified sites
C0489969|ICD9CM|AB|719.98|Joint dis NOS-oth jt
C0489970|ICD9CM|PT|743.32|Congenital cortical and zonular cataract
C0489970|ICD9CM|AB|743.32|Cortical/zonular catarac
C0489974|ICD9CM|PT|996.94|Complications of reattached upper extremity, other and unspecified
C0489974|ICD9CM|AB|996.94|Compl reattached arm NEC
C0489976|ICD9CM|AB|49.91|Incision of anal septum
C0489976|ICD9CM|PT|49.91|Incision of anal septum
C0489977|ICD9CM|PT|66.51|Removal of both fallopian tubes at same operative episode
C0489977|ICD9CM|AB|66.51|Remove both fallop tubes
C0489980|ICD9CM|PT|031.2|Disseminated due to other mycobacteria
C0489980|ICD9CM|AB|031.2|DMAC bacteremia
C0489981|ICD9CM|PT|038.19|Other staphylococcal septicemia
C0489981|ICD9CM|AB|038.19|Staphylcocc septicem NEC
C0489982|ICD9CM|PT|275.49|Other disorders of calcium metabolism
C0489982|ICD9CM|AB|275.49|Dis calcium metablsm NEC
C0489983|ICD9CM|PT|438.0|Late effects of cerebrovascular disease, cognitive deficits
C0489983|ICD9CM|AB|438.0|Late ef CV dis-cognf def
C0489984|ICD9CM|HT|438.1|Speech and language deficits as late effect of cerebrovascular disease
C0489984|ICD9CM|PT|438.10|Late effects of cerebrovascular disease, speech and language deficit, unspecified
C0489984|ICD9CM|AB|438.10|Late ef-spch/lng def NOS
C0489985|ICD9CM|PT|438.11|Late effects of cerebrovascular disease, aphasia
C0489985|ICD9CM|AB|438.11|Late eff CV dis-aphasia
C0489986|ICD9CM|PT|438.12|Late effects of cerebrovascular disease, dysphasia
C0489986|ICD9CM|AB|438.12|Late eff CV dis-dysphsia
C0489987|ICD9CM|PT|438.19|Late effects of cerebrovascular disease, other speech and language deficits
C0489987|ICD9CM|AB|438.19|Late ef-spch/lang df NEC
C0489988|ICD9CM|HT|438.2|Hemiplegia/hemiparesis as late effect of cerebrovascular disease
C0489989|ICD9CM|PT|438.20|Late effects of cerebrovascular disease, hemiplegia affecting unspecified side
C0489989|ICD9CM|AB|438.20|Late ef-hemplga side NOS
C0489990|ICD9CM|PT|438.21|Late effects of cerebrovascular disease, hemiplegia affecting dominant side
C0489990|ICD9CM|AB|438.21|Late ef-hemplga dom side
C0489991|ICD9CM|PT|438.22|Late effects of cerebrovascular disease, hemiplegia affecting nondominant side
C0489991|ICD9CM|AB|438.22|Late ef-hemiplga non-dom
C0489992|ICD9CM|HT|438.3|Monoplegia of upper limb as late effect of cerebrovascular disease
C0489993|ICD9CM|PT|438.30|Late effects of cerebrovascular disease, monoplegia of upper limb affecting unspecified side
C0489993|ICD9CM|AB|438.30|Late ef-mplga up lmb NOS
C0489994|ICD9CM|PT|438.31|Late effects of cerebrovascular disease, monoplegia of upper limb affecting dominant side
C0489994|ICD9CM|AB|438.31|Late ef-mplga up lmb dom
C0489995|ICD9CM|PT|438.32|Late effects of cerebrovascular disease, monoplegia of upper limb affecting nondominant side
C0489995|ICD9CM|AB|438.32|Lt ef-mplga uplmb nondom
C0489996|ICD9CM|HT|438.4|Monoplegia of lower limb as late effect of cerebrovascular disease
C0489997|ICD9CM|PT|438.40|Late effects of cerebrovascular disease, monoplegia of lower limb affecting unspecified side
C0489997|ICD9CM|AB|438.40|Lte ef-mplga low lmb NOS
C0489998|ICD9CM|PT|438.41|Late effects of cerebrovascular disease, monoplegia of lower limb affecting dominant side
C0489998|ICD9CM|AB|438.41|Lte ef-mplga low lmb dom
C0489999|ICD9CM|PT|438.42|Late effects of cerebrovascular disease, monoplegia of lower limb affecting nondominant side
C0489999|ICD9CM|AB|438.42|Lt ef-mplga lowlmb nondm
C0490000|ICD9CM|HT|438.5|Other paralytic syndrome as late effect of cerebrovascular disease
C0490001|ICD9CM|PT|438.50|Late effects of cerebrovascular disease, other paralytic syndrome affecting unspecified side
C0490001|ICD9CM|AB|438.50|Lt ef oth paral side NOS
C0490002|ICD9CM|PT|438.51|Late effects of cerebrovascular disease, other paralytic syndrome affecting dominant side
C0490002|ICD9CM|AB|438.51|Lt ef oth paral dom side
C0490003|ICD9CM|PT|438.52|Late effects of cerebrovascular disease, other paralytic syndrome affecting nondominant side
C0490003|ICD9CM|AB|438.52|Lt ef oth parals non-dom
C0490004|ICD9CM|HT|438.8|Other late effects of cerebrovascular disease
C0490004|ICD9CM|PT|438.89|Other late effects of cerebrovascular disease
C0490004|ICD9CM|AB|438.89|Late effect CV dis NEC
C0490005|ICD9CM|PT|438.81|Other late effects of cerebrovascular disease, apraxia
C0490005|ICD9CM|AB|438.81|Late eff CV dis-apraxia
C0490006|ICD9CM|PT|438.82|Other late effects of cerebrovascular disease, dysphagia
C0490006|ICD9CM|AB|438.82|Late ef CV dis dysphagia
C0490007|ICD9CM|PT|458.8|Other specified hypotension
C0490007|ICD9CM|AB|458.8|Hypotension NEC
C0490008|ICD9CM|HT|655.7|Decreased fetal movements, affecting management of mother
C0490009|ICD9CM|PT|686.09|Other pyoderma
C0490009|ICD9CM|AB|686.09|Pyoderma NEC
C0490010|ICD9CM|PT|756.79|Other congenital anomalies of abdominal wall
C0490010|ICD9CM|AB|756.79|Congn anoml abd wall NEC
C0490011|ICD9CM|PT|780.39|Other convulsions
C0490011|ICD9CM|AB|780.39|Convulsions NEC
C0490012|ICD9CM|PT|796.5|Abnormal finding on antenatal screening
C0490012|ICD9CM|AB|796.5|Abn find antenatl screen
C0490013|ICD9CM|PT|V02.69|Other viral hepatitis carrier
C0490013|ICD9CM|AB|V02.69|Viral hep carrier NEC
C0490014|ICD9CM|PT|V12.41|Personal history of benign neoplasm of the brain
C0490014|ICD9CM|AB|V12.41|Hx benign neoplasm brain
C0490015|ICD9CM|PT|V12.49|Personal history of other disorders of nervous system and sense organs
C0490015|ICD9CM|AB|V12.49|Hx nerv sys/snse org NEC
C0490017|ICD9CM|PT|V16.41|Family history of malignant neoplasm of ovary
C0490017|ICD9CM|AB|V16.41|Fm hx ovary malignancy
C0490019|ICD9CM|PT|V16.43|Family history of malignant neoplasm of testis
C0490019|ICD9CM|AB|V16.43|Fm hx testis malig
C0490020|ICD9CM|PT|V16.49|Family history of malignant neoplasm of other genital organs
C0490020|ICD9CM|AB|V16.49|Fm hx genital malig NEC
C0490021|ICD9CM|PT|V28.6|Antenatal screening for Streptococcus B
C0490021|ICD9CM|AB|V28.6|Antenatal screen strep b
C0490022|ICD9CM|PT|V42.82|Peripheral stem cells replaced by transplant
C0490022|ICD9CM|AB|V42.82|Trspl sts-perip stm cell
C0490023|ICD9CM|HT|V42.8|Other specified organ or tissue replaced by transplant
C0490023|ICD9CM|PT|V42.89|Other specified organ or tissue replaced by transplant
C0490023|ICD9CM|AB|V42.89|Trnspl status organ NEC
C0490024|ICD9CM|AB|V45.61|Cataract extract status
C0490024|ICD9CM|PT|V45.61|Cataract extraction status
C0490025|ICD9CM|PT|V45.69|Other states following surgery of eye and adnexa
C0490025|ICD9CM|AB|V45.69|Post-proc st eye/adn NEC
C0490025|ICD9CM|HT|V45.6|States following surgery of eye and adnexa
C0490027|ICD9CM|PT|V45.72|Acquired absence of intestine (large) (small)
C0490027|ICD9CM|AB|V45.72|Acquire absnce intestine
C0490028|ICD9CM|PT|V53.01|Fitting and adjustment of cerebral ventricular (communicating) shunt
C0490028|ICD9CM|AB|V53.01|Adj cerebral vent shunt
C0490029|ICD9CM|PT|V53.02|Fitting and adjustment of neuropacemaker (brain) (peripheral nerve) (spinal cord)
C0490029|ICD9CM|AB|V53.02|Adjust neuropacemaker
C0490030|ICD9CM|HT|V64.4|Closed surgical procedure converted to open procedure
C0490031|ICD9CM|PT|V76.10|Breast screening, unspecified
C0490031|ICD9CM|AB|V76.10|Scrn mal neo breast NOS
C0490032|ICD9CM|PT|V76.11|Screening mammogram for high-risk patient
C0490032|ICD9CM|AB|V76.11|Screen mammogram hi risk
C0490033|ICD9CM|PT|V76.12|Other screening mammogram
C0490033|ICD9CM|AB|V76.12|Screen mammogram NEC
C0490034|ICD9CM|PT|V76.19|Other screening breast examination
C0490034|ICD9CM|AB|V76.19|Scrn mal neo breast NEC
C0490035|ICD9CM|PT|E922.4|Accident caused by air gun
C0490035|ICD9CM|AB|E922.4|Accident - air gun
C0490036|ICD9CM|PT|E955.6|Suicide and self-inflicted injury by air gun
C0490036|ICD9CM|AB|E955.6|Self inflict acc-air gun
C0490037|ICD9CM|PT|E968.6|Assault by air gun
C0490037|ICD9CM|AB|E968.6|Assault - air gun
C0490038|ICD9CM|PT|E985.6|Injury by air gun, undetermined whether accidental or purposely inflicted
C0490038|ICD9CM|AB|E985.6|Undetrmine accid-air gun
C0490039|ICD9CM|PT|041.04|Streptococcus infection in conditions classified elsewhere and of unspecified site, streptococcus, group D [Enterococcus]
C0490039|ICD9CM|AB|041.04|Enterococcus group d
C0490040|ICD9CM|HT|474.0|Chronic tonsillitis and adenoiditis
C0490040|ICD9CM|PT|474.02|Chronic tonsillitis and adenoiditis
C0490040|ICD9CM|AB|474.02|Chronic tonsils&adenoids
C0490041|ICD9CM|HT|959.0|Other and unspecified injury to head, face, and neck
C0490042|ICD9CM|HT|E922|Accident caused by firearm, and air gun missile
C0490043|ICD9CM|HT|E955|Suicide and self-inflicted injury by firearms, air guns, and explosives
C0490044|ICD9CM|HT|E985|Injury by firearms, air guns and explosives, undetermined whether accidentally or purposely inflicted
C0490045|ICD9CM|PT|59.12|Laparoscopic lysis of perivesical adhesions
C0490045|ICD9CM|AB|59.12|Lap lys perivesureth adh
C0490048|ICD9CM|PT|593.70|Vesicoureteral reflux unspecified or without reflux nephropathy
C0490048|ICD9CM|AB|593.70|Vescouretrl rflux unspcf
C0490049|ICD9CM|PT|647.21|Other venereal diseases of mother, complicating pregnancy, childbirth, or the puerperium, delivered, with or without mention of antepartum condition
C0490049|ICD9CM|AB|647.21|Other vd-delivered
C0490050|ICD9CM|PT|647.22|Other venereal diseases of mother, complicating pregnancy, childbirth, or the puerperium, delivered, with mention of postpartum complication
C0490050|ICD9CM|AB|647.22|Other vd-delivered w p/p
C0490051|ICD9CM|PT|664.14|Second-degree perineal laceration, postpartum condition or complication
C0490051|ICD9CM|AB|664.14|Del w 2 deg lac-postpart
C0490052|ICD9CM|AB|696.1|Other psoriasis
C0490052|ICD9CM|PT|696.1|Other psoriasis
C0490053|ICD9CM|PT|755.29|Longitudinal deficiency, phalanges, complete or partial
C0490053|ICD9CM|AB|755.29|Longitud defic phalanges
C0490054|ICD9CM|PT|755.39|Longitudinal deficiency, phalanges, complete or partial
C0490054|ICD9CM|AB|755.39|Longitud defic phalanges
C0490055|ICD9CM|PT|872.69|Open wound of other and multiple sites of ear, without mention of complication
C0490055|ICD9CM|AB|872.69|Open wound of ear NEC
C0490056|ICD9CM|PT|872.79|Open wound of other and multiple sites of ear, complicated
C0490056|ICD9CM|AB|872.79|Open wound ear NEC-compl
C0490057|ICD9CM|PT|873.49|Open wound of other and multiple sites of face, without mention of complication
C0490057|ICD9CM|AB|873.49|Open wound of face NEC
C0490058|ICD9CM|PT|873.59|Open wound of other and multiple sites of face, complicated
C0490058|ICD9CM|AB|873.59|Open wnd face NEC-compl
C0490059|ICD9CM|PT|873.69|Open wound of other and multiple sites of mouth, without mention of complication
C0490059|ICD9CM|AB|873.69|Open wound mouth NEC
C0490060|ICD9CM|PT|873.79|Open wound of other and multiple sites of mouth, complicated
C0490060|ICD9CM|AB|873.79|Open wnd mouth NOS-compl
C0490064|ICD9CM|PT|V29.9|Observation for unspecified suspected conditions
C0490064|ICD9CM|AB|V29.9|NB obsrv unsp suspct cnd
C0490065|ICD9CM|PT|V71.9|Observation for unspecified suspected condition
C0490065|ICD9CM|AB|V71.9|Observ-suspect cond NOS
C0490066|ICD9CM|AB|V72.2|Dental examination
C0490066|ICD9CM|PT|V72.2|Dental examination
C0490068|ICD9CM|PT|75.94|Immediate postpartum manual replacement of inverted uterus
C0490068|ICD9CM|AB|75.94|Man replac invert uterus
C0490069|ICD9CM|PT|83.83|Tendon pulley reconstruction other than hand
C0490069|ICD9CM|AB|83.83|Tendon pulley reconstruc
C0494024|ICD9CM|PT|008.09|Intestinal infection due to other intestinal E. coli infections
C0494024|ICD9CM|AB|008.09|Int inf e coli spcf NEC
C0494025|ICD9CM|PT|008.45|Intestinal infection due to Clostridium difficile
C0494025|ICD9CM|AB|008.45|Int inf clstrdium dfcile
C0494040|ICD9CM|AB|023.3|Brucella canis
C0494040|ICD9CM|PT|023.3|Brucella canis
C0494126|ICD9CM|HT|128|Other and unspecified helminthiases
C0494158|ICD9CM|PT|189.0|Malignant neoplasm of kidney, except pelvis
C0494158|ICD9CM|AB|189.0|Malig neopl kidney
C0494164|ICD9CM|PT|197.4|Secondary malignant neoplasm of small intestine including duodenum
C0494164|ICD9CM|AB|197.4|Sec malig neo sm bowel
C0494165|ICD9CM|PT|197.7|Malignant neoplasm of liver, secondary
C0494165|ICD9CM|AB|197.7|Second malig neo liver
C0494350|ICD9CM|PT|277.09|Cystic fibrosis with other manifestations
C0494350|ICD9CM|AB|277.09|Cystic fibrosis NEC
C0494362|ICD9CM|HT|277.8|Other specified disorders of metabolism
C0494362|ICD9CM|PT|277.89|Other specified disorders of metabolism
C0494362|ICD9CM|AB|277.89|Metabolism disorder NEC
C0494432|ICD9CM|PT|312.4|Mixed disturbance of conduct and emotions
C0494432|ICD9CM|AB|312.4|Mix dis conduct/emotion
C0494479|ICD9CM|HT|339|Other headache syndromes
C0494479|ICD9CM|PT|339.89|Other headache syndromes
C0494479|ICD9CM|HT|339-339.99|OTHER HEADACHE SYNDROMES
C0494479|ICD9CM|AB|339.89|Headache syndrome NEC
C0494553|ICD9CM|HT|380.3|Noninfectious disorders of pinna
C0494574|ICD9CM|PT|403.90|Hypertensive chronic kidney disease, unspecified, with chronic kidney disease stage I through stage IV, or unspecified
C0494574|ICD9CM|AB|403.90|Hy kid NOS w cr kid I-IV
C0494576|ICD9CM|PT|404.93|Hypertensive heart and chronic kidney disease, unspecified, with heart failure and chronic kidney disease stage V or end stage renal disease
C0494576|ICD9CM|AB|404.93|Hyp ht/kd NOS st V w hf
C0494580|ICD9CM|PT|410.70|Subendocardial infarction, episode of care unspecified
C0494580|ICD9CM|AB|410.70|Subendo infarct, unspec
C0494620|ICD9CM|PT|444.21|Arterial embolism and thrombosis of upper extremity
C0494620|ICD9CM|AB|444.21|Upper extremity embolism
C0494657|ICD9CM|HT|478.3|Paralysis of vocal cords or larynx
C0494675|ICD9CM|PT|507.1|Pneumonitis due to inhalation of oils and essences
C0494675|ICD9CM|AB|507.1|Oil/essence pneumonitis
C0494723|ICD9CM|HT|531.6|Chronic or unspecified gastric ulcer with hemorrhage and perforation
C0494726|ICD9CM|HT|532.6|Chronic or unspecified duodenal ulcer with hemorrhage and perforation
C0494730|ICD9CM|HT|533.4|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage
C0494731|ICD9CM|HT|533.5|Chronic or unspecified peptic ulcer of unspecified site with perforation
C0494732|ICD9CM|HT|533.6|Chronic or unspecified peptic ulcer of unspecified site with hemorrhage and perforation
C0494735|ICD9CM|HT|534.6|Chronic or unspecified gastrojejunal ulcer with hemorrhage and perforation
C0494736|ICD9CM|HT|534.9|Gastrojejunal ulcer, unspecified as acute or chronic, without mention of hemorrhage or perforation
C0494741|ICD9CM|PT|537.9|Unspecified disorder of stomach and duodenum
C0494741|ICD9CM|AB|537.9|Gastroduodenal dis NOS
C0494752|ICD9CM|PT|553.3|Diaphragmatic hernia without mention of obstruction or gangrene
C0494752|ICD9CM|AB|553.3|Diaphragmatic hernia
C0494776|ICD9CM|HT|564.8|Other specified functional disorders of intestine
C0494831|ICD9CM|AB|691.8|Other atopic dermatitis
C0494831|ICD9CM|PT|691.8|Other atopic dermatitis and related conditions
C0494843|ICD9CM|PT|693.1|Dermatitis due to food taken internally
C0494843|ICD9CM|AB|693.1|Dermat d/t food ingest
C0495094|ICD9CM|PT|620.4|Prolapse or hernia of ovary and fallopian tube
C0495094|ICD9CM|AB|620.4|Prolapse of ovary & tube
C0495106|ICD9CM|AB|624.01|Vulvar intraeph neopl I
C0495106|ICD9CM|PT|624.01|Vulvar intraepithelial neoplasia I [VIN I]
C0495107|ICD9CM|AB|624.02|Vulvr intraepth neopl II
C0495107|ICD9CM|PT|624.02|Vulvar intraepithelial neoplasia II [VIN II]
C0495168|ICD9CM|PT|639.1|Delayed or excessive hemorrhage following abortion or ectopic and molar pregnancies
C0495168|ICD9CM|AB|639.1|Postabortion hemorrhage
C0495169|ICD9CM|PT|639.6|Embolism following abortion or ectopic and molar pregnancies
C0495169|ICD9CM|AB|639.6|Postabortion embolism
C0495170|ICD9CM|PT|639.5|Shock following abortion or ectopic and molar pregnancies
C0495170|ICD9CM|AB|639.5|Postabortion shock
C0495172|ICD9CM|PT|639.4|Metabolic disorders following abortion or ectopic and molar pregnancies
C0495172|ICD9CM|AB|639.4|Postabort metabolic dis
C0495173|ICD9CM|PT|639.2|Damage to pelvic organs and tissues following abortion or ectopic and molar pregnancies
C0495173|ICD9CM|AB|639.2|Postabort pelvic damage
C0495184|ICD9CM|PT|671.93|Unspecified venous complication of pregnancy and the puerperium, antepartum condition or complication
C0495184|ICD9CM|AB|671.93|Venous compl NOS-antepar
C0495246|ICD9CM|HT|658.2|Delayed delivery after spontaneous or unspecified rupture of membranes
C0495255|ICD9CM|HT|661.4|Hypertonic, incoordinate, or prolonged uterine contractions
C0495263|ICD9CM|HT|660.7|Failed forceps or vacuum extractor, unspecified
C0495270|ICD9CM|HT|663.5|Vasa previa complicating labor and delivery
C0495270|ICD9CM|AB|663.50|Vasa previa-unspecified
C0495270|ICD9CM|PT|663.50|Vasa previa complicating labor and delivery, unspecified as to episode of care or not applicable
C0495289|ICD9CM|PT|671.24|Superficial thrombophlebitis complicating pregnancy and the puerperium, postpartum condition or complication
C0495289|ICD9CM|AB|671.24|Thrombophlebit-postpart
C0495308|ICD9CM|HT|647.2|Other venereal diseases in the mother complicating pregnancy, childbirth, or the puerperium
C0495310|ICD9CM|HT|647.8|Other specified infectious and parasitic diseases complicating pregnancy, childbirth, or the puerperium
C0495350|ICD9CM|PT|763.9|Unspecified complication of labor and delivery affecting fetus or newborn
C0495350|ICD9CM|AB|763.9|Compl deliv NOS aff NB
C0495351|ICD9CM|PT|763.5|Maternal anesthesia and analgesia affecting fetus or newborn
C0495351|ICD9CM|AB|763.5|Mat anesth/analg aff NB
C0495447|ICD9CM|PT|775.5|Other transitory neonatal electrolyte disturbances
C0495447|ICD9CM|AB|775.5|Neonatal dehydration
C0495615|ICD9CM|PT|756.0|Anomalies of skull and face bones
C0495615|ICD9CM|AB|756.0|Anomal skull/face bones
C0495689|ICD9CM|PT|781.1|Disturbances of sensation of smell and taste
C0495689|ICD9CM|AB|781.1|Smell & taste disturb
C0495691|ICD9CM|HT|799.2|Signs and symptoms involving emotional state
C0495795|ICD9CM|HT|794.1|Nonspecific abnormal results of function study of peripheral nervous system and special senses
C0495833|ICD9CM|PT|901.1|Injury to innominate and subclavian arteries
C0495833|ICD9CM|AB|901.1|Inj innomin/subclav art
C0495858|ICD9CM|PT|880.09|Open wound of multiple sites of shoulder and upper arm, without mention of complication
C0495858|ICD9CM|AB|880.09|Mult open wound shoulder
C0496029|ICD9CM|HT|941.0|Burn of face, head, and neck, unspecified degree
C0496137|ICD9CM|HT|996|Complications peculiar to certain specified procedures
C0496180|ICD9CM|PT|909.0|Late effect of poisoning due to drug, medicinal or biological substance
C0496180|ICD9CM|AB|909.0|Late eff drug poisoning
C0496530|ICD9CM|PT|E871.7|Foreign object left in body during removal of catheter or packing
C0496530|ICD9CM|AB|E871.7|FB post-catheter removal
C0496542|ICD9CM|PT|E878.3|Surgical operation with formation of external stoma causing abnormal patient reaction, or later complication, without mention of misadventure at time of operation
C0496542|ICD9CM|AB|E878.3|Abn react-external stoma
C0496613|ICD9CM|AB|V03.3|Vaccin for plague
C0496613|ICD9CM|PT|V03.3|Need for prophylactic vaccination and inoculation against plague
C0496614|ICD9CM|PT|V03.4|Need for prophylactic vaccination and inoculation against tularemia
C0496614|ICD9CM|AB|V03.4|Vaccin for tularemia
C0496615|ICD9CM|PT|V03.7|Need for prophylactic vaccination and inoculation against tetanus toxoid alone
C0496615|ICD9CM|AB|V03.7|Tetanus toxoid inoculat
C0496621|ICD9CM|PT|V04.4|Need for prophylactic vaccination and inoculation against yellow fever
C0496621|ICD9CM|AB|V04.4|Vaccin for yellow fever
C0496634|ICD9CM|PT|V06.4|Need for prophylactic vaccination and inoculation against measles-mumps-rubella (MMR)
C0496634|ICD9CM|AB|V06.4|Vac-measle-mumps-rubella
C0496640|ICD9CM|HT|V26.4|General counseling and advice on procreative management
C0496648|ICD9CM|PT|V28.1|Antenatal screening for raised alpha-fetoprotein levels in amniotic fluid
C0496648|ICD9CM|AB|V28.1|Screen-alphafetoprotein
C0496656|ICD9CM|HT|V33.0|Twin, unspecified, born in hospital
C0496662|ICD9CM|PT|V24.0|Postpartum care and examination immediately after delivery
C0496662|ICD9CM|AB|V24.0|Postpart care after del
C0496668|ICD9CM|PT|V53.90|Fitting and adjustment, unspecified device
C0496668|ICD9CM|AB|V53.90|Fit/adjust device NOS
C0496682|ICD9CM|AB|V62.0|Unemployment
C0496682|ICD9CM|PT|V62.0|Unemployment
C0496703|ICD9CM|AB|V65.2|Person feigning illness
C0496703|ICD9CM|PT|V65.2|Person feigning illness
C0496709|ICD9CM|PT|V19.0|Family history of blindness or visual loss
C0496709|ICD9CM|AB|V19.0|Family hx-blindness
C0496716|ICD9CM|HT|V18.5|Family history of digestive disorders
C0496723|ICD9CM|HT|V12.4|Personal history of disorders of nervous system and sense organs
C0496723|ICD9CM|PT|V12.40|Personal history of unspecified disorder of nervous system and sense organs
C0496723|ICD9CM|AB|V12.40|Hx nerv sys/snse org NOS
C0496750|ICD9CM|PT|V45.2|Presence of cerebrospinal fluid drainage device
C0496750|ICD9CM|AB|V45.2|Ventricular shunt status
C0496755|ICD9CM|PT|141.2|Malignant neoplasm of tip and lateral border of tongue
C0496755|ICD9CM|AB|141.2|Mal neo tip/lat tongue
C0496758|ICD9CM|PT|144.1|Malignant neoplasm of lateral portion of floor of mouth
C0496758|ICD9CM|AB|144.1|Mal neo lat floor mouth
C0496763|ICD9CM|HT|142|Malignant neoplasm of major salivary glands
C0496765|ICD9CM|PT|146.4|Malignant neoplasm of anterior aspect of epiglottis
C0496765|ICD9CM|AB|146.4|Mal neo ant epiglottis
C0496769|ICD9CM|PT|148.0|Malignant neoplasm of postcricoid region of hypopharynx
C0496769|ICD9CM|AB|148.0|Mal neo postcricoid
C0496770|ICD9CM|PT|148.3|Malignant neoplasm of posterior hypopharyngeal wall
C0496770|ICD9CM|AB|148.3|Mal neo post hypopharynx
C0496773|ICD9CM|PT|150.0|Malignant neoplasm of cervical esophagus
C0496773|ICD9CM|AB|150.0|Mal neo cervical esophag
C0496775|ICD9CM|PT|150.2|Malignant neoplasm of abdominal esophagus
C0496775|ICD9CM|AB|150.2|Mal neo abdomin esophag
C0496779|ICD9CM|PT|153.5|Malignant neoplasm of appendix vermiformis
C0496779|ICD9CM|AB|153.5|Malignant neo appendix
C0496814|ICD9CM|PT|184.1|Malignant neoplasm of labia majora
C0496814|ICD9CM|AB|184.1|Mal neo labia majora
C0496815|ICD9CM|PT|184.2|Malignant neoplasm of labia minora
C0496815|ICD9CM|AB|184.2|Mal neo labia minora
C0496826|ICD9CM|PT|188.0|Malignant neoplasm of trigone of urinary bladder
C0496826|ICD9CM|AB|188.0|Mal neo bladder-trigone
C0496827|ICD9CM|PT|188.1|Malignant neoplasm of dome of urinary bladder
C0496827|ICD9CM|AB|188.1|Mal neo bladder-dome
C0496828|ICD9CM|PT|188.2|Malignant neoplasm of lateral wall of urinary bladder
C0496828|ICD9CM|AB|188.2|Mal neo bladder-lateral
C0496836|ICD9CM|HT|190|Malignant neoplasm of eye
C0496836|ICD9CM|PT|190.9|Malignant neoplasm of eye, part unspecified
C0496836|ICD9CM|AB|190.9|Malign neopl eye NOS
C0496854|ICD9CM|PT|230.8|Carcinoma in situ of liver and biliary system
C0496854|ICD9CM|AB|230.8|Ca in situ liver/biliary
C0496858|ICD9CM|PT|210.2|Benign neoplasm of major salivary glands
C0496858|ICD9CM|AB|210.2|Ben neo major salivary
C0496872|ICD9CM|PT|211.7|Benign neoplasm of islets of Langerhans
C0496872|ICD9CM|AB|211.7|Ben neo islets langerhan
C0496876|ICD9CM|HT|215|Other benign neoplasm of connective and other soft tissue
C0496876|ICD9CM|PT|215.9|Other benign neoplasm of connective and other soft tissue, site unspecified
C0496876|ICD9CM|AB|215.9|Ben neo soft tissue NOS
C0496889|ICD9CM|PT|221.0|Benign neoplasm of fallopian tube and uterine ligaments
C0496889|ICD9CM|AB|221.0|Ben neo fallopian tube
C0496891|ICD9CM|HT|222|Benign neoplasm of male genital organs
C0496891|ICD9CM|PT|222.9|Benign neoplasm of male genital organ, site unspecified
C0496891|ICD9CM|AB|222.9|Ben neo male genital NOS
C0496893|ICD9CM|PT|223.9|Benign neoplasm of urinary organ, site unspecified
C0496893|ICD9CM|AB|223.9|Benign neo urinary NOS
C0496897|ICD9CM|HT|224|Benign neoplasm of eye
C0496897|ICD9CM|AB|224.9|Benign neoplasm eye NOS
C0496897|ICD9CM|PT|224.9|Benign neoplasm of eye, part unspecified
C0496899|ICD9CM|PT|225.0|Benign neoplasm of brain
C0496899|ICD9CM|AB|225.0|Benign neoplasm brain
C0496909|ICD9CM|PT|235.3|Neoplasm of uncertain behavior of liver and biliary passages
C0496909|ICD9CM|AB|235.3|Unc behav neo liver
C0496912|ICD9CM|PT|235.6|Neoplasm of uncertain behavior of larynx
C0496912|ICD9CM|AB|235.6|Unc behav neo larynx
C0496919|ICD9CM|PT|236.0|Neoplasm of uncertain behavior of uterus
C0496919|ICD9CM|AB|236.0|Uncert behav neo uterus
C0496920|ICD9CM|PT|236.2|Neoplasm of uncertain behavior of ovary
C0496920|ICD9CM|AB|236.2|Unc behav neo ovary
C0496921|ICD9CM|PT|236.1|Neoplasm of uncertain behavior of placenta
C0496921|ICD9CM|AB|236.1|Unc behav neo placenta
C0496923|ICD9CM|PT|236.5|Neoplasm of uncertain behavior of prostate
C0496923|ICD9CM|AB|236.5|Unc behav neo prostate
C0496924|ICD9CM|PT|236.4|Neoplasm of uncertain behavior of testis
C0496924|ICD9CM|AB|236.4|Unc behav neo testis
C0496930|ICD9CM|PT|236.7|Neoplasm of uncertain behavior of bladder
C0496930|ICD9CM|AB|236.7|Unc behav neo bladder
C0496932|ICD9CM|PT|236.90|Neoplasm of uncertain behavior of urinary organ, unspecified
C0496932|ICD9CM|AB|236.90|Unc behav neo urinar NOS
C0496946|ICD9CM|PT|237.1|Neoplasm of uncertain behavior of pineal gland
C0496946|ICD9CM|AB|237.1|Unc behav neo pineal
C0496955|ICD9CM|PT|238.2|Neoplasm of uncertain behavior of skin
C0496955|ICD9CM|AB|238.2|Unc behav neo skin
C0496956|ICD9CM|PT|238.3|Neoplasm of uncertain behavior of breast
C0496956|ICD9CM|AB|238.3|Unc behav neo breast
C0496964|ICD9CM|PT|961.6|Poisoning by anthelmintics
C0496964|ICD9CM|AB|961.6|Poisoning-anthelmintics
C0496967|ICD9CM|PT|962.3|Poisoning by insulins and antidiabetic agents
C0496967|ICD9CM|AB|962.3|Poison-insulin/antidiab
C0496978|ICD9CM|PT|969.05|Poisoning by tricyclic antidepressants
C0496978|ICD9CM|AB|969.05|Pois tricyclc antidepres
C0497026|ICD9CM|PT|988.1|Toxic effect of mushrooms eaten as food
C0497026|ICD9CM|AB|988.1|Toxic effect mushrooms
C0497073|ICD9CM|PT|E942.7|Antivaricose drugs, including sclerosing agents, causing adverse effects in therapeutic use
C0497073|ICD9CM|AB|E942.7|Adv eff antivaricose
C0497074|ICD9CM|PT|E942.9|Other and unspecified agents primarily affecting the cardiovascular system causing adverse effects in therapeutic use
C0497074|ICD9CM|AB|E942.9|Adv eff cardiovasc NEC
C0497076|ICD9CM|PT|E944.5|Electrolytic, caloric, and water-balance agents causing adverse effects in therapeutic use
C0497076|ICD9CM|AB|E944.5|Adv eff electrolyte agnt
C0497080|ICD9CM|PT|E872.1|Failure of sterile precautions during infusion or transfusion
C0497080|ICD9CM|AB|E872.1|Failure sterile infusion
C0497081|ICD9CM|PT|E872.3|Failure of sterile precautions during injection or vaccination
C0497081|ICD9CM|AB|E872.3|Fail sterile injection
C0497082|ICD9CM|PT|E872.4|Failure of sterile precautions during endoscopic examination
C0497082|ICD9CM|AB|E872.4|Fail sterile endoscopy
C0497083|ICD9CM|PT|E872.6|Failure of sterile precautions during heart catheterization
C0497083|ICD9CM|AB|E872.6|Fail sterile heart cath
C0497134|ICD9CM|PT|780.92|Excessive crying of infant (baby)
C0497134|ICD9CM|AB|780.92|Excess cry infant/baby
C0497217|ICD9CM|HT|379|Other disorders of eye
C0497327|ICD9CM|HT|290|Dementias
C0497327|ICD9CM|HT|294.2|Dementia, unspecified
C0497333|ICD9CM|HT|295-299.99|OTHER PSYCHOSES
C0497406|ICD9CM|AB|278.02|Overweight
C0497406|ICD9CM|PT|278.02|Overweight
C0497538|ICD9CM|HT|211|Benign neoplasm of other parts of digestive system
C0497538|ICD9CM|PT|211.9|Benign neoplasm of other and unspecified site in the digestive system
C0497538|ICD9CM|AB|211.9|Ben neo GI tract NEC/NOS
C0497550|ICD9CM|HT|225|Benign neoplasm of brain and other parts of nervous system
C0497550|ICD9CM|PT|225.9|Benign neoplasm of nervous system, part unspecified
C0497550|ICD9CM|AB|225.9|Benign neo nerv sys NOS
C0497552|ICD9CM|PT|742.9|Unspecified congenital anomaly of brain, spinal cord, and nervous system
C0497552|ICD9CM|AB|742.9|Nervous system anom NOS
C0498276|ICD9CM|PT|76.5|Temporomandibular arthroplasty
C0498276|ICD9CM|AB|76.5|Temporomand arthroplasty
C0519030|ICD9CM|PT|482.0|Pneumonia due to Klebsiella pneumoniae
C0519030|ICD9CM|AB|482.0|K. pneumoniae pneumonia
C0519129|ICD9CM|PT|60.96|Transurethral destruction of prostate tissue by microwave thermotherapy
C0519129|ICD9CM|AB|60.96|Tu destr prostate by mt
C0520473|ICD9CM|HT|290-294.99|ORGANIC PSYCHOTIC CONDITIONS
C0520474|ICD9CM|HT|733.4|Aseptic necrosis of bone
C0520474|ICD9CM|PT|733.40|Aseptic necrosis of bone, site unspecified
C0520474|ICD9CM|AB|733.40|Asept necrosis bone NOS
C0520482|ICD9CM|AB|300.81|Somatization disorder
C0520482|ICD9CM|PT|300.81|Somatization disorder
C0520556|ICD9CM|PT|685.1|Pilonidal cyst without mention of abscess
C0520556|ICD9CM|AB|685.1|Pilonidal cyst w/o absc
C0520569|ICD9CM|HT|553.0|Femoral hernia without mention of obstruction or gangrene
C0520575|ICD9CM|HT|590.1|Acute pyelonephritis
C0520578|ICD9CM|AB|752.52|Retractile testis
C0520578|ICD9CM|PT|752.52|Retractile testis
C0520578|ICD9CM|HT|752.5|Undescended and retractile testicle
C0520679|ICD9CM|AB|327.23|Obstructive sleep apnea
C0520679|ICD9CM|PT|327.23|Obstructive sleep apnea (adult)(pediatric)
C0520728|ICD9CM|AB|369.70|Low vision, one eye
C0520728|ICD9CM|PT|369.70|Moderate or severe impairment, one eye, impairment level not further specified
C0520806|ICD9CM|HT|798|Sudden death, cause unknown
C0520966|ICD9CM|AB|781.3|Lack of coordination
C0520966|ICD9CM|PT|781.3|Lack of coordination
C0521221|ICD9CM|PT|33.20|Thoracoscopic lung biopsy
C0521221|ICD9CM|AB|33.20|Thoracoscopc lung biopsy
C0521223|ICD9CM|PT|32.41|Thoracoscopic lobectomy of lung
C0521223|ICD9CM|AB|32.41|Thorac lobectomy lung
C0521224|ICD9CM|PT|32.50|Thoracoscopic pneumonectomy
C0521224|ICD9CM|AB|32.50|Thoracospc pneumonectomy
C0521232|ICD9CM|PT|36.06|Insertion of non-drug-eluting coronary artery stent(s)
C0521232|ICD9CM|AB|36.06|Ins nondrug elut cor st
C0521254|ICD9CM|PT|42.82|Suture of laceration of esophagus
C0521254|ICD9CM|AB|42.82|Suture esophageal lacer
C0521264|ICD9CM|PT|50.14|Laparoscopic liver biopsy
C0521264|ICD9CM|AB|50.14|Laparoscopic liver bx
C0521590|ICD9CM|PT|524.52|Limited mandibular range of motion
C0521590|ICD9CM|AB|524.52|Limited mandibular ROM
C0521620|ICD9CM|AB|593.5|Hydroureter
C0521620|ICD9CM|PT|593.5|Hydroureter
C0521648|ICD9CM|PT|770.84|Respiratory failure of newborn
C0521648|ICD9CM|AB|770.84|Resp failure of newborn
C0521668|ICD9CM|PT|339.43|Primary thunderclap headache
C0521668|ICD9CM|AB|339.43|Prim thnderclap headache
C0521709|ICD9CM|PT|369.02|Better eye: near-total vision impairment; lesser eye: not further specified
C0521709|ICD9CM|AB|369.02|One eye-near tot/oth-NOS
C0521710|ICD9CM|PT|369.61|One eye: total vision impairment; other eye: not specified
C0521710|ICD9CM|AB|369.61|One eye-total/oth-unknwn
C0521829|ICD9CM|PT|088.9|Arthropod-borne disease, unspecified
C0521829|ICD9CM|AB|088.9|Arthropod-borne dis NOS
C0522214|ICD9CM|PT|794.13|Nonspecific abnormal visually evoked potential
C0522214|ICD9CM|AB|794.13|Abnormal vep
C0522224|ICD9CM|AB|344.9|Paralysis NOS
C0522224|ICD9CM|PT|344.9|Paralysis, unspecified
C0522253|ICD9CM|PT|339.84|Primary exertional headache
C0522253|ICD9CM|AB|339.84|Prim exertion headache
C0522274|ICD9CM|HT|279.0|Deficiency of humoral immunity
C0522274|ICD9CM|PT|279.09|Other deficiency of humoral immunity
C0522274|ICD9CM|AB|279.09|Humoral immunity def NEC
C0522723|ICD9CM|AB|E004.3|Bungee jumping
C0522723|ICD9CM|PT|E004.3|Activities involving bungee jumping
C0524528|ICD9CM|HT|299.9|Unspecified pervasive developmental disorder
C0524528|ICD9CM|HT|299|Pervasive developmental disorders
C0524620|ICD9CM|AB|277.7|Dysmetabolic syndrome x
C0524620|ICD9CM|PT|277.7|Dysmetabolic syndrome X
C0524662|ICD9CM|AB|304.00|Opioid dependence-unspec
C0524662|ICD9CM|HT|304.0|Opioid type dependence
C0524662|ICD9CM|PT|304.00|Opioid type dependence, unspecified
C0524688|ICD9CM|AB|020.5|Pneumonic plague NOS
C0524688|ICD9CM|PT|020.5|Pneumonic plague, unspecified
C0524689|ICD9CM|PT|32.22|Lung volume reduction surgery
C0524689|ICD9CM|AB|32.22|Lung vol reduction surg
C0524850|ICD9CM|HT|01-05.99|OPERATIONS ON THE NERVOUS SYSTEM
C0542408|ICD9CM|HT|72.2|Mid forceps operation
C0543418|ICD9CM|HT|E941|Drugs primarily affecting the autonomic nervous system causing adverse effects in therapeutic use
C0543428|ICD9CM|HT|V02.6|Carrier or suspected carrier of viral hepatitis
C0544793|ICD9CM|PT|562.13|Diverticulitis of colon with hemorrhage
C0544793|ICD9CM|AB|562.13|Dvrtcli colon w hmrhg
C0546812|ICD9CM|HT|599|Other disorders of urethra and urinary tract
C0546817|ICD9CM|HT|276.6|Fluid overload
C0546819|ICD9CM|PT|313.22|Introverted disorder of childhood
C0546819|ICD9CM|AB|313.22|Introverted dis-child
C0546821|ICD9CM|PT|96.06|Insertion of Sengstaken tube
C0546821|ICD9CM|AB|96.06|Insert sengstaken tube
C0546823|ICD9CM|HT|62.9|Other operations on testes
C0546823|ICD9CM|PT|62.99|Other operations on testes
C0546823|ICD9CM|AB|62.99|Testicular operation NEC
C0546826|ICD9CM|PT|110.5|Dermatophytosis of the body
C0546826|ICD9CM|AB|110.5|Dermatophytosis of body
C0546827|ICD9CM|AB|126.8|Ancylostoma NEC
C0546827|ICD9CM|PT|126.8|Other specified ancylostoma
C0546830|ICD9CM|PT|E906.2|Bite of nonvenomous snakes and lizards
C0546830|ICD9CM|AB|E906.2|Nonvenomous snake bite
C0546831|ICD9CM|PT|E957.1|Suicide and self-inflicted injuries by jumping from other man-made structures
C0546831|ICD9CM|AB|E957.1|Injury-jump fm struc NEC
C0546834|ICD9CM|AB|95.23|Visual evoked potential
C0546834|ICD9CM|PT|95.23|Visual evoked potential [VEP]
C0546835|ICD9CM|PT|155.1|Malignant neoplasm of intrahepatic bile ducts
C0546835|ICD9CM|AB|155.1|Mal neo intrahepat ducts
C0546836|ICD9CM|PT|140.9|Malignant neoplasm of lip, unspecified, vermilion border
C0546836|ICD9CM|AB|140.9|Mal neo lip/vermil NOS
C0546837|ICD9CM|HT|150|Malignant neoplasm of esophagus
C0546837|ICD9CM|PT|150.9|Malignant neoplasm of esophagus, unspecified site
C0546837|ICD9CM|AB|150.9|Mal neo esophagus NOS
C0546839|ICD9CM|HT|359.8|Other myopathies
C0546839|ICD9CM|PT|359.89|Other myopathies
C0546839|ICD9CM|AB|359.89|Myopathies NEC
C0546840|ICD9CM|PT|716.59|Unspecified polyarthropathy or polyarthritis, multiple sites
C0546840|ICD9CM|AB|716.59|Polyarthritis NOS-mult
C0546841|ICD9CM|PT|E904.3|Accident due to exposure (to weather conditions), not elsewhere classifiable
C0546841|ICD9CM|AB|E904.3|Exposure NEC
C0546884|ICD9CM|AB|276.52|Hypovolemia
C0546884|ICD9CM|PT|276.52|Hypovolemia
C0546884|ICD9CM|HT|276.5|Volume depletion
C0546884|ICD9CM|AB|276.50|Volume depletion NOS
C0546884|ICD9CM|PT|276.50|Volume depletion, unspecified
C0546949|MTH|PN|NOCODE|Complications of medical care, NEC in ICD9CM_2014
C0546949|ICD9CM|HT|999|Complications of medical care, not elsewhere classified
C0546982|ICD9CM|PT|277.01|Cystic fibrosis with meconium ileus
C0546982|ICD9CM|AB|277.01|Cystic fibrosis w ileus
C0546983|ICD9CM|AB|310.2|Postconcussion syndrome
C0546983|ICD9CM|PT|310.2|Postconcussion syndrome
C0546996|ICD9CM|PT|120.3|Cutaneous schistosomiasis
C0546996|ICD9CM|AB|120.3|Cutaneous schistosoma
C0547030|ICD9CM|HT|368|Visual disturbances
C0547030|ICD9CM|AB|368.9|Visual disturbance NOS
C0547030|ICD9CM|PT|368.9|Unspecified visual disturbance
C0549102|ICD9CM|HT|08.2|Excision or destruction of lesion or tissue of eyelid
C0549103|ICD9CM|PT|08.20|Removal of lesion of eyelid, not otherwise specified
C0549103|ICD9CM|AB|08.20|Remove eyelid lesion NOS
C0549117|ICD9CM|AB|310.0|Frontal lobe syndrome
C0549117|ICD9CM|PT|310.0|Frontal lobe syndrome
C0549126|ICD9CM|PT|V02.60|Viral hepatitis carrier, unspecified
C0549126|ICD9CM|AB|V02.60|Viral hep carrier NOS
C0549147|MTH|PN|NOCODE|Cardiac complications, NEC in ICD9CM_2014
C0549147|ICD9CM|PT|997.1|Cardiac complications, not elsewhere classified
C0549147|ICD9CM|AB|997.1|Surg compl-heart
C0549160|ICD9CM|PT|082.2|North Asian tick fever
C0549160|ICD9CM|AB|082.2|North asian tick fever
C0549211|ICD9CM|PT|426.13|Other second degree atrioventricular block
C0549211|ICD9CM|AB|426.13|Av block-2nd degree NEC
C0549397|ICD9CM|AB|470|Deviated nasal septum
C0549397|ICD9CM|PT|470|Deviated nasal septum
C0549423|ICD9CM|PT|331.4|Obstructive hydrocephalus
C0549423|ICD9CM|AB|331.4|Obstructiv hydrocephalus
C0549470|ICD9CM|AB|365.00|Preglaucoma NOS
C0549470|ICD9CM|PT|365.00|Preglaucoma, unspecified
C0553526|ICD9CM|PT|985.4|Toxic effect of antimony and its compounds
C0553526|ICD9CM|AB|985.4|Toxic effect antimony
C0553570|ICD9CM|AB|454.0|Leg varicosity w ulcer
C0553570|ICD9CM|PT|454.0|Varicose veins of lower extremities with ulcer
C0553604|ICD9CM|HT|359.2|Myotonic disorders
C0553651|MTH|PN|NOCODE|PHYSICAL THERAPY NEC in ICD9CM
C0553651|ICD9CM|PT|93.39|Other physical therapy
C0553651|ICD9CM|AB|93.39|Physical therapy NEC
C0553716|ICD9CM|PT|618.1|Uterine prolapse without mention of vaginal wall prolapse
C0553716|ICD9CM|AB|618.1|Uterine prolapse
C0553730|ICD9CM|HT|712.2|Chondrocalcinosis due to pyrophosphate crystals
C0553730|ICD9CM|HT|712.3|Chondrocalcinosis, cause unspecified
C0553730|ICD9CM|PT|712.20|Chondrocalcinosis, due to pyrophosphate crystals, site unspecified
C0553730|ICD9CM|AB|712.20|Pyrophosph cryst-unspec
C0553794|ICD9CM|AB|03.31|Spinal tap
C0553794|ICD9CM|PT|03.31|Spinal tap
C0553977|ICD9CM|PT|421.0|Acute and subacute bacterial endocarditis
C0553977|ICD9CM|AB|421.0|Ac/subac bact endocard
C0553980|ICD9CM|AB|425.0|Endomyocardial fibrosis
C0553980|ICD9CM|PT|425.0|Endomyocardial fibrosis
C0553983|ICD9CM|HT|443|Other peripheral vascular disease
C0553983|ICD9CM|PT|443.89|Other specified peripheral vascular diseases
C0553983|ICD9CM|AB|443.89|Periph vascular dis NEC
C0554121|ICD9CM|PT|550.13|Inguinal hernia, with obstruction, without mention of gangrene, bilateral, recurrent
C0554121|ICD9CM|AB|550.13|Recur bil ing hern-obstr
C0554123|ICD9CM|PT|550.10|Inguinal hernia, with obstruction, without mention of gangrene, unilateral or unspecified (not specified as recurrent)
C0554123|ICD9CM|AB|550.10|Unilat ing hernia w obst
C0554139|ICD9CM|PT|55.87|Correction of ureteropelvic junction
C0554139|ICD9CM|AB|55.87|Correct ureteropelv junc
C0554472|ICD9CM|HT|704|Diseases of hair and hair follicles
C0554472|ICD9CM|AB|704.9|Hair disease NOS
C0554472|ICD9CM|PT|704.9|Unspecified disease of hair and hair follicles
C0554585|ICD9CM|AB|77.57|Repair of claw toe
C0554585|ICD9CM|PT|77.57|Repair of claw toe
C0554588|ICD9CM|PT|719.05|Effusion of joint, pelvic region and thigh
C0554588|ICD9CM|AB|719.05|Joint effusion-pelvis
C0554634|ICD9CM|PT|090.7|Late congenital syphilis, unspecified
C0554634|ICD9CM|AB|090.7|Late congen syph NOS
C0555219|ICD9CM|PT|751.5|Other anomalies of intestine
C0555219|ICD9CM|AB|751.5|Intestinal anomaly NEC
C0555264|ICD9CM|HT|150-159.99|MALIGNANT NEOPLASM OF DIGESTIVE ORGANS AND PERITONEUM
C0555295|ICD9CM|HT|883|Open wound of finger(s)
C0555330|ICD9CM|HT|812.4|Fracture of lower end of humerus, closed
C0555330|ICD9CM|PT|812.40|Closed fracture of unspecified part of lower end of humerus
C0555330|ICD9CM|AB|812.40|Fx lower humerus NOS-cl
C0555332|ICD9CM|HT|812.5|Fracture of lower end of humerus, open
C0555332|ICD9CM|PT|812.50|Open fracture of unspecified part of lower end of humerus
C0555332|ICD9CM|AB|812.50|Fx lower humer NOS-open
C0555347|ICD9CM|PT|823.82|Closed fracture of unspecified part of fibula with tibia
C0555347|ICD9CM|HT|823.8|Fracture of unspecified part of tibia and fibula, closed
C0555347|ICD9CM|AB|823.82|Fx tibia w fibula NOS-cl
C0556856|ICD9CM|PT|93.56|Application of pressure dressing
C0556856|ICD9CM|AB|93.56|Pressure dressing applic
C0558156|ICD9CM|AB|707.01|Pressure ulcer, elbow
C0558156|ICD9CM|PT|707.01|Pressure ulcer, elbow
C0558158|ICD9CM|AB|707.07|Pressure ulcer, heel
C0558158|ICD9CM|PT|707.07|Pressure ulcer, heel
C0558160|ICD9CM|AB|707.05|Pressure ulcer, buttock
C0558160|ICD9CM|PT|707.05|Pressure ulcer, buttock
C0558338|ICD9CM|PT|66.8|Insufflation of fallopian tube
C0558338|ICD9CM|AB|66.8|Fallopian tube insufflat
C0558421|ICD9CM|HT|915|Superficial injury of finger(s)
C0558960|ICD9CM|PT|E954|Suicide and self-inflicted injury by submersion [drowning]
C0558960|ICD9CM|AB|E954|Injury-submersion
C0558995|ICD9CM|HT|097|Other and unspecified syphilis
C0559043|ICD9CM|HT|805|Fracture of vertebral column without mention of spinal cord injury
C0559051|ICD9CM|HT|E913|Accidental mechanical suffocation
C0559702|ICD9CM|PT|80.21|Arthroscopy, shoulder
C0559702|ICD9CM|AB|80.21|Shoulder arthroscopy
C0562512|ICD9CM|HT|893|Open wound of toe(s)
C0563449|ICD9CM|AB|752.62|Epispadias
C0563449|ICD9CM|PT|752.62|Epispadias
C0563536|ICD9CM|PT|08.91|Electrosurgical epilation of eyelid
C0563536|ICD9CM|AB|08.91|Electrosurg lid epilat
C0564567|ICD9CM|AB|799.23|Impulsiveness
C0564567|ICD9CM|PT|799.23|Impulsiveness
C0565375|ICD9CM|PT|66.63|Bilateral partial salpingectomy, not otherwise specified
C0565375|ICD9CM|AB|66.63|Bilat part salpingec NOS
C0565454|ICD9CM|PT|75.0|Intra-amniotic injection for abortion
C0565454|ICD9CM|AB|75.0|Intra-amnion inj for ab
C0565840|ICD9CM|HT|66.0|Salpingotomy and salpingostomy
C0565864|ICD9CM|PT|93.93|Nonmechanical methods of resuscitation
C0565864|ICD9CM|AB|93.93|Nonmechan resuscitation
C0565898|ICD9CM|AB|E922.1|Shotgun accident
C0565898|ICD9CM|PT|E922.1|Accident caused by shotgun (automatic)
C0566742|ICD9CM|HT|663.1|Cord around neck, with compression, complicating labor and delivery
C0569621|ICD9CM|PT|E940.9|Unspecified central nervous system stimulant causing adverse effects in therapeutic use
C0569621|ICD9CM|HT|E940|Central nervous system stimulants causing adverse effects in therapeutic use
C0569621|ICD9CM|AB|E940.9|Adv eff cns stimulnt NOS
C0575081|ICD9CM|AB|781.2|Abnormality of gait
C0575081|ICD9CM|PT|781.2|Abnormality of gait
C0576748|ICD9CM|PT|04.01|Excision of acoustic neuroma
C0576748|ICD9CM|AB|04.01|Excision acoustc neuroma
C0576995|ICD9CM|AB|784.8|Hemorrhage from throat
C0576995|ICD9CM|PT|784.8|Hemorrhage from throat
C0577712|ICD9CM|AB|707.04|Pressure ulcer, hip
C0577712|ICD9CM|PT|707.04|Pressure ulcer, hip
C0577713|ICD9CM|AB|707.06|Pressure ulcer, ankle
C0577713|ICD9CM|PT|707.06|Pressure ulcer, ankle
C0577719|ICD9CM|AB|707.12|Ulcer of calf
C0577719|ICD9CM|PT|707.12|Ulcer of calf
C0579036|ICD9CM|PT|86.26|Ligation of dermal appendage
C0579036|ICD9CM|AB|86.26|Ligation dermal appendag
C0580546|ICD9CM|HT|790.2|Abnormal glucose
C0581582|ICD9CM|AB|92.11|Cerebral scan
C0581582|ICD9CM|PT|92.11|Cerebral scan
C0581628|ICD9CM|PT|88.74|Diagnostic ultrasound of digestive system
C0581628|ICD9CM|AB|88.74|Dx ultrasound-digestive
C0581654|ICD9CM|PT|88.24|Skeletal x-ray of upper limb, not otherwise specified
C0581654|ICD9CM|AB|88.24|Skel xray-upper limb NOS
C0581655|ICD9CM|PT|88.29|Skeletal x-ray of lower limb, not otherwise specified
C0581655|ICD9CM|AB|88.29|Skel xray-lower limb NOS
C0582114|ICD9CM|PT|V49.86|Do not resuscitate status
C0582114|ICD9CM|AB|V49.86|Do not resusctate status
C0584793|ICD9CM|PT|385.21|Impaired mobility of malleus
C0584793|ICD9CM|AB|385.21|Ankylosis malleus
C0585100|ICD9CM|PT|44.38|Laparoscopic gastroenterostomy
C0585100|ICD9CM|AB|44.38|Lap gastroenterostomy
C0585464|ICD9CM|PT|17.33|Laparoscopic right hemicolectomy
C0585464|ICD9CM|AB|17.33|Lap right hemicolectomy
C0585968|ICD9CM|PT|V12.55|Personal history of pulmonary embolism
C0585968|ICD9CM|AB|V12.55|Hx pulmonary embolism
C0587245|ICD9CM|HT|536.4|Gastrostomy complications
C0587245|ICD9CM|PT|536.40|Gastrostomy complication, unspecified
C0587245|ICD9CM|AB|536.40|Gastrostomy comp NOS
C0587909|ICD9CM|PT|33.43|Closure of laceration of lung
C0587909|ICD9CM|AB|33.43|Lung laceration closure
C0587958|ICD9CM|PT|14.41|Scleral buckling with implant
C0587958|ICD9CM|AB|14.41|Scleral buckle w implant
C0595943|MTH|PN|NOCODE|Urinary complications, NEC in ICD9CM_2014
C0595943|ICD9CM|PT|997.5|Urinary complications, not elsewhere classified
C0595943|ICD9CM|AB|997.5|Surg compl-urinary tract
C0595979|ICD9CM|PT|009.1|Colitis, enteritis, and gastroenteritis of presumed infectious origin
C0595979|ICD9CM|AB|009.1|Enteritis of infect orig
C0595983|ICD9CM|PT|379.57|Deficiencies of saccadic eye movements
C0595983|ICD9CM|AB|379.57|Saccadic eye movmnt def
C0598894|ICD9CM|HT|206|Monocytic leukemia
C0598894|ICD9CM|HT|206.9|Unspecified monocytic leukemia
C0599986|ICD9CM|AB|V26.33|Genetic counseling
C0599986|ICD9CM|PT|V26.33|Genetic counseling
C0600000|ICD9CM|HT|26|Operations on salivary glands and ducts
C0600027|ICD9CM|PT|V79.9|Screening for unspecified mental disorder and developmental handicap
C0600027|ICD9CM|AB|V79.9|Screen-mental dis NOS
C0600040|ICD9CM|PT|595.1|Chronic interstitial cystitis
C0600040|ICD9CM|AB|595.1|Chr interstit cystitis
C0600042|ICD9CM|PT|635.81|Legally induced abortion, with unspecified complication, incomplete
C0600042|ICD9CM|AB|635.81|Leg ab w compl NOS-inc
C0600043|ICD9CM|PT|635.91|Legally induced abortion, without mention of complication, incomplete
C0600043|ICD9CM|AB|635.91|Legal abort uncompl-inc
C0600057|ICD9CM|HT|40|Operations on lymphatic system
C0600126|ICD9CM|HT|433.1|Occlusion and stenosis of carotid artery
C0600298|ICD9CM|AB|523.5|Periodontosis
C0600298|ICD9CM|PT|523.5|Periodontosis
C0600327|ICD9CM|AB|040.82|Toxic shock syndrome
C0600327|ICD9CM|PT|040.82|Toxic shock syndrome
C0600336|ICD9CM|PT|694.1|Subcorneal pustular dermatosis
C0600336|ICD9CM|AB|694.1|Subcorneal pust dermatos
C0600427|ICD9CM|HT|304.2|Cocaine dependence
C0600427|ICD9CM|PT|304.20|Cocaine dependence, unspecified
C0600427|ICD9CM|AB|304.20|Cocaine depend-unspec
C0600452|ICD9CM|PT|573.5|Hepatopulmonary syndrome
C0600452|ICD9CM|AB|573.5|Hepatopulmonary syndrome
C0677061|ICD9CM|AB|724.1|Pain in thoracic spine
C0677061|ICD9CM|PT|724.1|Pain in thoracic spine
C0677491|ICD9CM|PT|V42.0|Kidney replaced by transplant
C0677491|ICD9CM|AB|V42.0|Kidney transplant status
C0677519|ICD9CM|AB|E928.2|Exposure to vibration
C0677519|ICD9CM|PT|E928.2|Vibration
C0677545|ICD9CM|PT|290.10|Presenile dementia, uncomplicated
C0677545|ICD9CM|AB|290.10|Presenile dementia
C0677548|ICD9CM|AB|V21.1|Puberty
C0677548|ICD9CM|PT|V21.1|Puberty
C0677577|MTH|PN|NOCODE|Dwarfism, NEC in ICD9CM_2014
C0677577|ICD9CM|PT|259.4|Dwarfism, not elsewhere classified
C0677577|ICD9CM|AB|259.4|Dwarfism NEC
C0677586|ICD9CM|HT|426.5|Bundle branch block, other and unspecified
C0677607|ICD9CM|PT|245.2|Chronic lymphocytic thyroiditis
C0677607|ICD9CM|AB|245.2|Chr lymphocyt thyroidit
C0677614|ICD9CM|AB|V66.9|Convalescence NOS
C0677614|ICD9CM|PT|V66.9|Unspecified convalescence
C0677631|ICD9CM|AB|V42.2|Heart valve transplant
C0677631|ICD9CM|PT|V42.2|Heart valve replaced by transplant
C0677639|ICD9CM|AB|V62.4|Social maladjustment
C0677639|ICD9CM|PT|V62.4|Social maladjustment
C0677640|ICD9CM|PT|115.90|Histoplasmosis, unspecified, without mention of manifestation
C0677640|ICD9CM|AB|115.90|Histoplasmosis NOS
C0678189|ICD9CM|PT|272.0|Pure hypercholesterolemia
C0678189|ICD9CM|AB|272.0|Pure hypercholesterolem
C0678202|ICD9CM|HT|555|Regional enteritis
C0678202|ICD9CM|AB|555.9|Regional enteritis NOS
C0678202|ICD9CM|PT|555.9|Regional enteritis of unspecified site
C0683416|ICD9CM|PT|300.6|Depersonalization disorder
C0683416|ICD9CM|AB|300.6|Depersonalization disord
C0684250|ICD9CM|PT|V42.83|Pancreas replaced by transplant
C0684250|ICD9CM|AB|V42.83|Trnspl status-pancreas
C0684255|ICD9CM|PT|V62.82|Bereavement, uncomplicated
C0684255|ICD9CM|AB|V62.82|Bereavement, uncomplicat
C0684333|ICD9CM|PT|141.3|Malignant neoplasm of ventral surface of tongue
C0684333|ICD9CM|AB|141.3|Mal neo ventral tongue
C0685874|ICD9CM|AB|744.05|Anomalies of inner ear
C0685874|ICD9CM|PT|744.05|Anomalies of inner ear
C0685898|ICD9CM|HT|995.6|Anaphylactic reaction due to food
C0685925|ICD9CM|PT|524.63|Temporomandibular joint disorders, articular disc disorder (reducing or non-reducing)
C0685925|ICD9CM|AB|524.63|Articular disc disorder
C0686277|ICD9CM|AB|233.31|Carcinoma in situ vagina
C0686277|ICD9CM|PT|233.31|Carcinoma in situ, vagina
C0686546|ICD9CM|PT|200.27|Burkitt's tumor or lymphoma, spleen
C0686546|ICD9CM|AB|200.27|Burkitt's tumor spleen
C0686560|ICD9CM|PT|201.00|Hodgkin's paragranuloma, unspecified site, extranodal and solid organ sites
C0686560|ICD9CM|AB|201.00|Hdgk prg unsp xtrndl org
C0686574|ICD9CM|PT|202.61|Malignant mast cell tumors, lymph nodes of head, face, and neck
C0686574|ICD9CM|AB|202.61|Mal mastocytosis head
C0686584|ICD9CM|PT|208.91|Unspecified leukemia, in remission
C0686584|ICD9CM|AB|208.91|Leukemia NOS w remission
C0686586|ICD9CM|PT|208.01|Acute leukemia of unspecified cell type, in remission
C0686586|ICD9CM|AB|208.01|Act leuk uns cl w rmson
C0686589|ICD9CM|PT|208.11|Chronic leukemia of unspecified cell type, in remission
C0686589|ICD9CM|AB|208.11|Chr leuk uns cl w rmson
C0686591|ICD9CM|PT|208.21|Subacute leukemia of unspecified cell type, in remission
C0686591|ICD9CM|AB|208.21|Sbac leuk uns cl w rmson
C0686593|ICD9CM|PT|205.91|Unspecified myeloid leukemia, in remission
C0686593|ICD9CM|AB|205.91|Uns myl leuk w rmsion
C0686595|ICD9CM|PT|206.91|Unspecified monocytic leukemia, in remission
C0686595|ICD9CM|AB|206.91|Uns mono leuk w rmsion
C0686597|ICD9CM|PT|204.91|Unspecified lymphoid leukemia, in remission
C0686597|ICD9CM|AB|204.91|Uns lym leuk w rmsion
C0686619|ICD9CM|HT|196|Secondary and unspecified malignant neoplasm of lymph nodes
C0686619|ICD9CM|PT|196.9|Secondary and unspecified malignant neoplasm of lymph nodes, site unspecified
C0686619|ICD9CM|AB|196.9|Mal neo lymph node NOS
C0686645|ICD9CM|PT|196.1|Secondary and unspecified malignant neoplasm of intrathoracic lymph nodes
C0686645|ICD9CM|AB|196.1|Mal neo lymph-intrathor
C0686655|ICD9CM|PT|196.2|Secondary and unspecified malignant neoplasm of intra-abdominal lymph nodes
C0686655|ICD9CM|AB|196.2|Mal neo lymph intra-abd
C0686689|ICD9CM|PT|196.6|Secondary and unspecified malignant neoplasm of intrapelvic lymph nodes
C0686689|ICD9CM|AB|196.6|Mal neo lymph-intrapelv
C0686705|ICD9CM|HT|934|Foreign body in trachea, bronchus, and lung
C0686721|ICD9CM|PT|995.55|Shaken baby syndrome
C0686721|ICD9CM|AB|995.55|Shaken infant syndrome
C0687122|ICD9CM|PT|93.53|Application of other cast
C0687122|ICD9CM|AB|93.53|Other cast application
C0687129|ICD9CM|AB|V60.0|Lack of housing
C0687129|ICD9CM|PT|V60.0|Lack of housing
C0687718|ICD9CM|PT|571.9|Unspecified chronic liver disease without mention of alcohol
C0687718|ICD9CM|AB|571.9|Chronic liver dis NOS
C0687719|MTH|PN|NOCODE|Autoimmune disease NEC in ICD9CM
C0687719|ICD9CM|AB|279.49|Autoimmune disease NEC
C0687719|ICD9CM|HT|279.4|Autoimmune disease, not elsewhere classified
C0687719|ICD9CM|PT|279.49|Autoimmune disease, not elsewhere classified
C0687762|ICD9CM|HT|263|Other and unspecified protein-calorie malnutrition
C0694548|ICD9CM|AB|493.82|Cough variant asthma
C0694548|ICD9CM|PT|493.82|Cough variant asthma
C0694551|ICD9CM|PT|789.03|Abdominal pain, right lower quadrant
C0694551|ICD9CM|AB|789.03|Abdmnal pain rt lwr quad
C0695214|ICD9CM|PT|655.70|Decreased fetal movements, affecting management of mother, unspecified as to episode of care
C0695214|ICD9CM|AB|655.70|Decrease fetl movmt unsp
C0695215|ICD9CM|PT|655.71|Decreased fetal movements, affecting management of mother, delivered, with or without mention of antepartum condition
C0695215|ICD9CM|AB|655.71|Decrease fetal movmt del
C0695216|ICD9CM|PT|655.73|Decreased fetal movements, affecting management of mother, antepartum condition or complication
C0695216|ICD9CM|AB|655.73|Dec fetal movmt antepart
C0695217|ICD9CM|PT|851.09|Cortex (cerebral) contusion without mention of open intracranial wound, with concussion, unspecified
C0695217|ICD9CM|AB|851.09|Cortex contus-concus NOS
C0695221|ICD9CM|PT|851.49|Cerebellar or brain stem contusion without mention of open intracranial wound, with concussion, unspecified
C0695221|ICD9CM|AB|851.49|Cerebell contus-concuss
C0695222|ICD9CM|PT|851.59|Cerebellar or brain stem contusion with open intracranial wound, with concussion, unspecified
C0695222|ICD9CM|AB|851.59|Opn cerebel cont-concuss
C0695223|ICD9CM|PT|851.69|Cerebellar or brain stem laceration without mention of open intracranial wound, with concussion, unspecified
C0695223|ICD9CM|AB|851.69|Cerebel lacer-concussion
C0695224|ICD9CM|PT|851.79|Cerebellar or brain stem laceration with open intracranial wound, with concussion, unspecified
C0695224|ICD9CM|AB|851.79|Opn cerebell lac-concuss
C0695225|ICD9CM|PT|851.89|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with concussion, unspecified
C0695225|ICD9CM|AB|851.89|Brain lacer NEC-concuss
C0695226|ICD9CM|PT|851.99|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with concussion, unspecified
C0695226|ICD9CM|AB|851.99|Open brain lacer-concuss
C0695231|ICD9CM|PT|V23.7|Supervision of high-risk pregnancy with insufficient prenatal care
C0695231|ICD9CM|AB|V23.7|Insufficnt prenatal care
C0695232|ICD9CM|PT|438.53|Late effects of cerebrovascular disease, other paralytic syndrome, bilateral
C0695232|ICD9CM|AB|438.53|Lt ef oth parals-bilat
C0695234|ICD9CM|PT|482.49|Other Staphylococcus pneumonia
C0695234|ICD9CM|AB|482.49|Staph pneumonia NEC
C0695236|ICD9CM|AB|519.01|Tracheostomy infection
C0695236|ICD9CM|PT|519.01|Infection of tracheostomy
C0695237|ICD9CM|PT|519.02|Mechanical complication of tracheostomy
C0695237|ICD9CM|AB|519.02|Tracheostomy - mech comp
C0695238|ICD9CM|PT|519.09|Other tracheostomy complications
C0695238|ICD9CM|AB|519.09|Tracheostomy comp NEC
C0695239|ICD9CM|AB|536.41|Gastrostomy infection
C0695239|ICD9CM|PT|536.41|Infection of gastrostomy
C0695240|ICD9CM|PT|536.42|Mechanical complication of gastrostomy
C0695240|ICD9CM|AB|536.42|Gastrostomy comp - mech
C0695241|ICD9CM|PT|536.49|Other gastrostomy complications
C0695241|ICD9CM|AB|536.49|Gastrostomy comp NEC
C0695242|ICD9CM|AB|564.81|Neurogenic bowel
C0695242|ICD9CM|PT|564.81|Neurogenic bowel
C0695243|ICD9CM|PT|569.62|Mechanical complication of colostomy and enterostomy
C0695243|ICD9CM|AB|569.62|Colosty/enter comp-mech
C0695244|ICD9CM|PT|V23.82|Supervision of high-risk pregnancy with elderly multigravida
C0695244|ICD9CM|AB|V23.82|Suprv elderly multigrav
C0695245|ICD9CM|HT|659.7|Abnormality in fetal heart rate or rhythm
C0695246|ICD9CM|PT|659.70|Abnormality in fetal heart rate or rhythm, unspecified as to episode of care or not applicable
C0695246|ICD9CM|AB|659.70|Abn ftl hrt rate/rhy-uns
C0695247|ICD9CM|PT|659.71|Abnormality in fetal heart rate or rhythm, delivered, with or without mention of antepartum condition
C0695247|ICD9CM|AB|659.71|Abn ftl hrt rate/rhy-del
C0695248|ICD9CM|PT|659.73|Abnormality in fetal heart rate or rhythm, antepartum condition or complication
C0695248|ICD9CM|AB|659.73|Abn ftl hrt rate/rhy-ant
C0695249|ICD9CM|PT|763.81|Abnormality in fetal heart rate or rhythm before the onset of labor
C0695249|ICD9CM|AB|763.81|Ab ftl hrt rt/rh b/f lab
C0695250|ICD9CM|PT|763.82|Abnormality in fetal heart rate or rhythm during labor
C0695250|ICD9CM|AB|763.82|Ab ftl hrt rt/rh dur lab
C0695251|ICD9CM|PT|763.83|Abnormality in fetal heart rate or rhythm, unspecified as to time of onset
C0695251|ICD9CM|AB|763.83|Ab ftl hrt rt/rhy NOS
C0695252|ICD9CM|PT|780.79|Other malaise and fatigue
C0695252|ICD9CM|AB|780.79|Malaise and fatigue NEC
C0695253|ICD9CM|PT|965.69|Poisoning by other antirheumatics
C0695253|ICD9CM|AB|965.69|Poison-antirheumatic NEC
C0695254|ICD9CM|PT|996.55|Mechanical complication due to artificial skin graft and decellularized allodermis
C0695254|ICD9CM|AB|996.55|Comp-artificial skin grf
C0695255|ICD9CM|PT|996.56|Mechanical complication due to peritoneal dialysis catheter
C0695255|ICD9CM|AB|996.56|Comp-periton dialys cath
C0695256|ICD9CM|PT|996.68|Infection and inflammatory reaction due to peritoneal dialysis catheter
C0695256|ICD9CM|AB|996.68|React-periton dialy cath
C0695257|ICD9CM|PT|V02.52|Carrier or suspected carrier of other streptococcus
C0695257|ICD9CM|AB|V02.52|Streptococus carrier NEC
C0695259|ICD9CM|PT|V18.69|Family history of other kidney diseases
C0695259|ICD9CM|AB|V18.69|Fam hx-kidney dis NEC
C0695260|ICD9CM|PT|V23.83|Supervision of high-risk pregnancy with young primigravida
C0695260|ICD9CM|AB|V23.83|Suprv young primigravida
C0695261|ICD9CM|PT|V23.84|Supervision of high-risk pregnancy with young multigravida
C0695261|ICD9CM|AB|V23.84|Suprv young multigravida
C0695263|ICD9CM|HT|V26.5|Sterilization status
C0695264|ICD9CM|AB|V26.51|Tubal ligation status
C0695264|ICD9CM|PT|V26.51|Tubal ligation status
C0695265|ICD9CM|AB|V26.52|Vasectomy status
C0695265|ICD9CM|PT|V26.52|Vasectomy status
C0695266|ICD9CM|PT|V29.3|Observation for suspected genetic or metabolic condition
C0695266|ICD9CM|AB|V29.3|NB obs genetc/metabl cnd
C0695272|ICD9CM|PT|V82.4|Maternal postnatal screening for chromosomal anomalies
C0695272|ICD9CM|AB|V82.4|Mat pstntl scr-chrm anom
C0695273|ICD9CM|PT|V43.83|Artificial skin replacement
C0695273|ICD9CM|AB|V43.83|Artific skin repl status
C0695274|ICD9CM|PT|965.61|Poisoning by propionic acid derivatives
C0695274|ICD9CM|AB|965.61|Pois-propionic acid derv
C0699739|ICD9CM|PT|356.2|Hereditary sensory neuropathy
C0699739|ICD9CM|AB|356.2|Hered sensory neuropathy
C0699815|ICD9CM|PT|783.3|Feeding difficulties and mismanagement
C0699815|ICD9CM|AB|783.3|Feeding problem
C0699895|ICD9CM|AB|V26.1|Artificial insemination
C0699895|ICD9CM|PT|V26.1|Artificial insemination
C0699899|ICD9CM|PT|723.7|Ossification of posterior longitudinal ligament in cervical region
C0699899|ICD9CM|AB|723.7|Ossification cerv lig
C0699916|ICD9CM|PT|V76.44|Screening for malignant neoplasms of prostate
C0699916|ICD9CM|AB|V76.44|Scrn malig neop-prostate
C0699976|ICD9CM|AB|91.95|Toxicology NOS
C0699976|ICD9CM|PT|91.95|Microscopic examination of specimen from unspecified site, toxicology
C0700102|ICD9CM|PT|V16.51|Family history of malignant neoplasm of kidney
C0700102|ICD9CM|AB|V16.51|Family hx-kidney malig
C0700112|ICD9CM|PT|V10.48|Personal history of malignant neoplasm of epididymis
C0700112|ICD9CM|AB|V10.48|Hx-epididymis malignancy
C0700143|ICD9CM|PT|201.17|Hodgkin's granuloma, spleen
C0700143|ICD9CM|AB|201.17|Hodgkins granulom spleen
C0700172|ICD9CM|AB|V04.6|Vaccin for mumps
C0700172|ICD9CM|PT|V04.6|Need for prophylactic vaccination and inoculation against mumps alone
C0700173|ICD9CM|AB|V04.2|Vaccin for measles
C0700173|ICD9CM|PT|V04.2|Need for prophylactic vaccination and inoculation against measles alone
C0700174|ICD9CM|AB|V04.3|Vaccin for rubella
C0700174|ICD9CM|PT|V04.3|Need for prophylactic vaccination and inoculation against rubella alone
C0700211|ICD9CM|HT|070.3|Viral hepatitis B without mention of hepatic coma
C0700232|ICD9CM|PT|V13.69|Personal history of other (corrected) congenital malformations
C0700232|ICD9CM|AB|V13.69|Hx-congenital malfor NEC
C0700292|ICD9CM|AB|799.02|Hypoxemia
C0700292|ICD9CM|PT|799.02|Hypoxemia
C0700297|ICD9CM|PT|V02.51|Carrier or suspected carrier of group B streptococcus
C0700297|ICD9CM|AB|V02.51|Group b streptoc carrier
C0700322|ICD9CM|AB|V61.5|Multiparity
C0700322|ICD9CM|PT|V61.5|Multiparity
C0700345|ICD9CM|AB|112.1|Candidal vulvovaginitis
C0700345|ICD9CM|PT|112.1|Candidiasis of vulva and vagina
C0700433|ICD9CM|PT|V73.99|Special screening examination for unspecified viral disease
C0700433|ICD9CM|HT|V73.9|Screening examination for unspecified viral disease
C0700433|ICD9CM|AB|V73.99|Scrn unspcf viral dis
C0700498|ICD9CM|HT|V61.2|Parent-child problems
C0700501|ICD9CM|AB|379.51|Congenital nystagmus
C0700501|ICD9CM|PT|379.51|Congenital nystagmus
C0700502|ICD9CM|HT|244|Acquired hypothyroidism
C0700503|ICD9CM|PT|053.0|Herpes zoster with meningitis
C0700503|ICD9CM|AB|053.0|Herpes zoster meningitis
C0700508|ICD9CM|HT|361.3|Retinal defects without detachment
C0700510|ICD9CM|PT|552.3|Diaphragmatic hernia with obstruction
C0700510|ICD9CM|AB|552.3|Diaphragm hernia w obstr
C0700516|ICD9CM|HT|V13.0|Personal history of disorders of urinary system
C0700522|ICD9CM|AB|E928.1|Exposure to noise
C0700522|ICD9CM|PT|E928.1|Exposure to noise
C0700573|ICD9CM|HT|V22|Normal pregnancy
C0700587|ICD9CM|AB|759.0|Anomalies of spleen
C0700587|ICD9CM|PT|759.0|Anomalies of spleen
C0700588|ICD9CM|PT|537.0|Acquired hypertrophic pyloric stenosis
C0700588|ICD9CM|AB|537.0|Acq pyloric stenosis
C0700613|ICD9CM|HT|300.0|Anxiety states
C0700613|ICD9CM|AB|300.00|Anxiety state NOS
C0700613|ICD9CM|PT|300.00|Anxiety state, unspecified
C0700615|ICD9CM|HT|659.6|Elderly multigravida
C0700625|MTH|PN|NOCODE|Allergy, unspecified, NEC in ICD9CM
C0700625|ICD9CM|AB|995.3|Allergy, unspecified
C0700625|ICD9CM|PT|995.3|Allergy, unspecified, not elsewhere classified
C0700639|ICD9CM|PT|750.5|Congenital hypertrophic pyloric stenosis
C0700639|ICD9CM|AB|750.5|Cong pyloric stenosis
C0700643|ICD9CM|PT|767.3|Other injuries to skeleton due to birth trauma
C0700643|ICD9CM|AB|767.3|Bone injury NEC at birth
C0700644|ICD9CM|PT|114.1|Primary extrapulmonary coccidioidomycosis
C0700644|ICD9CM|AB|114.1|Prim cutan coccidioid
C0700645|ICD9CM|AB|V50.3|Ear piercing
C0700645|ICD9CM|PT|V50.3|Ear piercing
C0701144|ICD9CM|PT|774.1|Perinatal jaundice from other excessive hemolysis
C0701144|ICD9CM|AB|774.1|Perinat jaund:hemolysis
C0701146|ICD9CM|PT|743.44|Specified congenital anomalies of anterior chamber, chamber angle, and related structures
C0701146|ICD9CM|AB|743.44|Anom anter chamber-eye
C0701156|ICD9CM|PT|34.92|Injection into thoracic cavity
C0701156|ICD9CM|AB|34.92|Inject into thorax cavit
C0701157|ICD9CM|HT|287.3|Primary thrombocytopenia
C0701162|ICD9CM|PT|253.4|Other anterior pituitary disorders
C0701162|ICD9CM|AB|253.4|Anter pituitary dis NEC
C0701163|ICD9CM|AB|255.2|Adrenogenital disorders
C0701163|ICD9CM|PT|255.2|Adrenogenital disorders
C0701168|ICD9CM|PT|424.2|Tricuspid valve disorders, specified as nonrheumatic
C0701168|ICD9CM|AB|424.2|Nonrheum tricusp val dis
C0701169|ICD9CM|PT|84.14|Amputation of ankle through malleoli of tibia and fibula
C0701169|ICD9CM|AB|84.14|Amputat through malleoli
C0701795|ICD9CM|PT|349.0|Reaction to spinal or lumbar puncture
C0701795|ICD9CM|AB|349.0|Lumbar puncture reaction
C0701804|ICD9CM|PT|54.22|Biopsy of abdominal wall or umbilicus
C0701804|ICD9CM|AB|54.22|Abdominal wall biopsy
C0701814|ICD9CM|PT|715.18|Osteoarthrosis, localized, primary, other specified sites
C0701814|ICD9CM|AB|715.18|Loc prim osteoarthr NEC
C0701822|ICD9CM|PT|246.0|Disorders of thyrocalcitonin secretion
C0701822|ICD9CM|AB|246.0|Dis thyrocalciton secret
C0701825|ICD9CM|HT|383.0|Acute mastoiditis
C0701828|ICD9CM|PT|34.3|Excision or destruction of lesion or tissue of mediastinum
C0701828|ICD9CM|AB|34.3|Destruct mediastin les
C0701842|ICD9CM|PT|84.02|Amputation and disarticulation of thumb
C0701842|ICD9CM|AB|84.02|Thumb amputation
C0701843|ICD9CM|PT|77.54|Excision or correction of bunionette
C0701843|ICD9CM|AB|77.54|Exc correct bunionette
C0701844|ICD9CM|PT|96.36|Irrigation of gastrostomy or enterostomy
C0701844|ICD9CM|AB|96.36|GI ostomy irrigation
C0702090|ICD9CM|PT|E871.0|Foreign object left in body during surgical operation
C0702090|ICD9CM|AB|E871.0|Post-surgical forgn body
C0702139|ICD9CM|PT|744.01|Absence of external ear
C0702139|ICD9CM|AB|744.01|Cong absence ext ear
C0702141|ICD9CM|AB|333.3|Tics of organic origin
C0702141|ICD9CM|PT|333.3|Tics of organic origin
C0702143|ICD9CM|AB|378.81|Palsy of conjugate gaze
C0702143|ICD9CM|PT|378.81|Palsy of conjugate gaze
C0702151|ICD9CM|HT|50.6|Repair of liver
C0702152|ICD9CM|AB|51.72|Choledochoplasty
C0702152|ICD9CM|PT|51.72|Choledochoplasty
C0702159|ICD9CM|HT|284.0|Constitutional aplastic anemia
C0702197|ICD9CM|PT|213.2|Benign neoplasm of vertebral column, excluding sacrum and coccyx
C0702197|ICD9CM|AB|213.2|Benign neo vertebrae
C0702266|ICD9CM|PT|288.65|Basophilia
C0702266|ICD9CM|AB|288.65|Basophilia
C0728716|ICD9CM|PT|81.40|Repair of hip, not elsewhere classified
C0728716|ICD9CM|AB|81.40|Repair of hip, NEC
C0728813|ICD9CM|HT|669.6|Breech extraction, without mention of indication
C0728829|ICD9CM|AB|754.71|Talipes cavus
C0728829|ICD9CM|PT|754.71|Talipes cavus
C0728859|ICD9CM|AB|V04.5|Vaccin for rabies
C0728859|ICD9CM|PT|V04.5|Need for prophylactic vaccination and inoculation against rabies
C0728864|ICD9CM|PT|160.0|Malignant neoplasm of nasal cavities
C0728864|ICD9CM|AB|160.0|Mal neo nasal cavities
C0728871|ICD9CM|PT|98.28|Removal of foreign body from foot without incision
C0728871|ICD9CM|AB|98.28|Removal FB from foot
C0728903|ICD9CM|PT|202.88|Other malignant lymphomas, lymph nodes of multiple sites
C0728903|ICD9CM|AB|202.88|Lymphomas NEC mult
C0728908|ICD9CM|PT|V42.84|Organ or tissue replaced by transplant, intestines
C0728908|ICD9CM|AB|V42.84|Trnspl status-intestines
C0728910|ICD9CM|HT|074|Specific diseases due to Coxsackie virus
C0728936|ICD9CM|PT|459.9|Unspecified circulatory system disorder
C0728936|ICD9CM|HT|390-459.99|DISEASES OF THE CIRCULATORY SYSTEM
C0728936|ICD9CM|AB|459.9|Circulatory disease NOS
C0728950|ICD9CM|AB|787.03|Vomiting alone
C0728950|ICD9CM|PT|787.03|Vomiting alone
C0728984|ICD9CM|AB|V41.0|Problems with sight
C0728984|ICD9CM|PT|V41.0|Problems with sight
C0729205|ICD9CM|PT|634.91|Spontaneous abortion, without mention of complication, incomplete
C0729205|ICD9CM|AB|634.91|Spon abort uncompl-inc
C0729233|ICD9CM|PT|441.01|Dissection of aorta, thoracic
C0729233|ICD9CM|AB|441.01|Dsct of thoracic aorta
C0729250|MTH|PN|NOCODE|Respiratory complications, NEC in ICD9CM_2014
C0729250|ICD9CM|HT|997.3|Respiratory complications, not elsewhere classified
C0729258|ICD9CM|AB|44.31|High gastric bypass
C0729258|ICD9CM|PT|44.31|High gastric bypass
C0729262|ICD9CM|PT|564.01|Slow transit constipation
C0729262|ICD9CM|AB|564.01|Slow transt constipation
C0730032|ICD9CM|PT|510.9|Empyema without mention of fistula
C0730032|ICD9CM|AB|510.9|Empyema w/o fistula
C0730276|ICD9CM|PT|362.04|Mild nonproliferative diabetic retinopathy
C0730276|ICD9CM|AB|362.04|Mild nonprolf db retnoph
C0730277|ICD9CM|PT|362.05|Moderate nonproliferative diabetic retinopathy
C0730277|ICD9CM|AB|362.05|Mod nonprolf db retinoph
C0730278|ICD9CM|PT|362.06|Severe nonproliferative diabetic retinopathy
C0730278|ICD9CM|AB|362.06|Sev nonprolf db retinoph
C0730285|ICD9CM|AB|362.07|Diabetic macular edema
C0730285|ICD9CM|PT|362.07|Diabetic macular edema
C0730328|ICD9CM|PT|362.41|Central serous retinopathy
C0730328|ICD9CM|AB|362.41|Cent serous retinopathy
C0730421|ICD9CM|PT|V65.42|Counseling on substance use and abuse
C0730421|ICD9CM|AB|V65.42|Counslng sbstn use abuse
C0730521|ICD9CM|PT|765.21|Less than 24 completed weeks of gestation
C0730521|ICD9CM|AB|765.21|<24 comp wks gestation
C0730522|ICD9CM|PT|765.22|24 completed weeks of gestation
C0730522|ICD9CM|AB|765.22|24 comp weeks gestation
C0730554|ICD9CM|PT|V15.41|History of physical abuse
C0730554|ICD9CM|AB|V15.41|Hx of physical abuse
C0730556|ICD9CM|PT|V15.42|History of emotional abuse
C0730556|ICD9CM|AB|V15.42|Hx of emotional abuse
C0733455|ICD9CM|PT|378.87|Other dissociated deviation of eye movements
C0733455|ICD9CM|AB|378.87|Skew deviation, eye
C0733940|ICD9CM|PT|140.4|Malignant neoplasm of lower lip, inner aspect
C0733940|ICD9CM|AB|140.4|Mal neo lower lip, inner
C0740080|ICD9CM|HT|V03.8|Need for other specified vaccinations against single bacterial diseases
C0740088|ICD9CM|PT|V12.50|Personal history of unspecified circulatory disease
C0740088|ICD9CM|AB|V12.50|Hx-circulatory dis NOS
C0740089|ICD9CM|PT|V12.70|Personal history of unspecified digestive disease
C0740089|ICD9CM|AB|V12.70|Prsnl hst unspc dgstv ds
C0740177|ICD9CM|PT|V23.81|Supervision of high-risk pregnancy with elderly primigravida
C0740177|ICD9CM|AB|V23.81|Suprv elderly primigrav
C0740179|ICD9CM|PT|V42.81|Bone marrow replaced by transplant
C0740179|ICD9CM|AB|V42.81|Trnspl status-bne marrow
C0740181|ICD9CM|AB|V50.0|Hair transplant
C0740181|ICD9CM|PT|V50.0|Elective hair transplant for purposes other than remedying health states
C0740203|ICD9CM|HT|V55|Attention to artificial openings
C0740203|ICD9CM|PT|V55.9|Attention to unspecified artificial opening
C0740203|ICD9CM|AB|V55.9|Attn to artif open NOS
C0740209|ICD9CM|AB|V65.40|Counseling NOS
C0740209|ICD9CM|PT|V65.40|Counseling NOS
C0740225|ICD9CM|AB|V82.6|Multiphasic screening
C0740225|ICD9CM|PT|V82.6|Multiphasic screening
C0740253|ICD9CM|AB|510.0|Empyema with fistula
C0740253|ICD9CM|PT|510.0|Empyema with fistula
C0740287|ICD9CM|PT|42.92|Dilation of esophagus
C0740287|ICD9CM|AB|42.92|Esophageal dilation
C0740331|ICD9CM|PT|279.05|Immunodeficiency with increased IgM
C0740331|ICD9CM|AB|279.05|Immunodefic w hyper-igm
C0741085|ICD9CM|AB|707.13|Ulcer of ankle
C0741085|ICD9CM|PT|707.13|Ulcer of ankle
C0741160|ICD9CM|PT|441.5|Aortic aneurysm of unspecified site, ruptured
C0741160|ICD9CM|AB|441.5|Rupt aortic aneurysm NOS
C0741305|ICD9CM|AB|380.03|Chondritis of pinna
C0741305|ICD9CM|PT|380.03|Chondritis of pinna
C0741439|ICD9CM|PT|288.66|Bandemia
C0741439|ICD9CM|AB|288.66|Bandemia
C0741646|ICD9CM|PT|675.13|Abscess of breast associated with childbirth, antepartum condition or complication
C0741646|ICD9CM|AB|675.13|Breast abscess-antepart
C0741804|ICD9CM|PT|519.11|Acute bronchospasm
C0741804|ICD9CM|AB|519.11|Acute bronchospasm
C0742343|ICD9CM|AB|517.3|Acute chest syndrome
C0742343|ICD9CM|PT|517.3|Acute chest syndrome
C0744374|ICD9CM|HT|629.2|Female genital mutilation status
C0744374|ICD9CM|AB|629.20|Genital mutilation NOS
C0744374|ICD9CM|PT|629.20|Female genital mutilation status, unspecified
C0744667|ICD9CM|PT|389.15|Sensorineural hearing loss, unilateral
C0744667|ICD9CM|AB|389.15|Sensorneur hear loss uni
C0745890|ICD9CM|PT|337.22|Reflex sympathetic dystrophy of the lower limb
C0745890|ICD9CM|AB|337.22|Rflx sym dystrph lwr lmb
C0746674|ICD9CM|PT|728.87|Muscle weakness (generalized)
C0746674|ICD9CM|AB|728.87|Muscle weakness-general
C0747273|ICD9CM|PT|142.0|Malignant neoplasm of parotid gland
C0747273|ICD9CM|AB|142.0|Malig neo parotid
C0747817|ICD9CM|AB|647.13|Gonorrhea-antepartum
C0747817|ICD9CM|PT|647.13|Gonorrhea of mother, complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C0747820|ICD9CM|AB|647.43|Malaria-antepartum
C0747820|ICD9CM|PT|647.43|Malaria in the mother, antepartum condition or complication
C0747833|ICD9CM|AB|647.03|Syphilis-antepartum
C0747833|ICD9CM|PT|647.03|Syphilis of mother, complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C0747834|ICD9CM|PT|648.13|Thyroid dysfunction of mother, antepartum condition or complication
C0747834|ICD9CM|AB|648.13|Thyroid dysfunc-antepart
C0748012|ICD9CM|HT|600.1|Nodular prostate
C0748659|ICD9CM|PT|660.41|Shoulder (girdle) dystocia, delivered, with or without mention of antepartum condition
C0748659|ICD9CM|AB|660.41|Shoulder dystocia-deliv
C0748830|ICD9CM|HT|801|Fracture of base of skull
C0749165|ICD9CM|HT|464.5|Supraglottitis, unspecified
C0749173|ICD9CM|AB|840.6|Sprain supraspinatus
C0749173|ICD9CM|PT|840.6|Supraspinatus (muscle) (tendon) sprain
C0749794|ICD9CM|PT|755.50|Unspecified anomaly of upper limb
C0749794|ICD9CM|AB|755.50|Upper limb anomaly NOS
C0750394|ICD9CM|HT|288.5|Decreased white blood cell count
C0750426|ICD9CM|HT|288.6|Elevated white blood cell count
C0750862|ICD9CM|AB|89.31|Dental examination
C0750862|ICD9CM|PT|89.31|Dental examination
C0750887|ICD9CM|PT|194.0|Malignant neoplasm of adrenal gland
C0750887|ICD9CM|AB|194.0|Malign neopl adrenal
C0750903|ICD9CM|AB|368.01|Strabismic amblyopia
C0750903|ICD9CM|PT|368.01|Strabismic amblyopia
C0750952|ICD9CM|PT|156.9|Malignant neoplasm of biliary tract, part unspecified site
C0750952|ICD9CM|AB|156.9|Malig neo biliary NOS
C0751057|ICD9CM|PT|780.32|Complex febrile convulsions
C0751057|ICD9CM|AB|780.32|Complx febrile convulsns
C0751098|ICD9CM|HT|062|Mosquito-borne viral encephalitis
C0751098|ICD9CM|PT|062.9|Mosquito-borne viral encephalitis, unspecified
C0751098|ICD9CM|AB|062.9|Mosquit-borne enceph NOS
C0751185|ICD9CM|PT|339.83|Primary cough headache
C0751185|ICD9CM|AB|339.83|Primary cough headache
C0751191|ICD9CM|PT|339.85|Primary stabbing headache
C0751191|ICD9CM|AB|339.85|Prim stabbing headache
C0751226|ICD9CM|AB|327.13|Recurrent hypersomnia
C0751226|ICD9CM|PT|327.13|Recurrent hypersomnia
C0751295|ICD9CM|AB|780.93|Memory loss
C0751295|ICD9CM|PT|780.93|Memory loss
C0751343|ICD9CM|AB|323.63|Postinfectious myelitis
C0751343|ICD9CM|PT|323.63|Postinfectious myelitis
C0751362|ICD9CM|HT|347|Cataplexy and narcolepsy
C0751362|ICD9CM|PT|347.01|Narcolepsy, with cataplexy
C0751362|ICD9CM|AB|347.01|Narcolepsy w cataplexy
C0751552|ICD9CM|PT|164.0|Malignant neoplasm of thymus
C0751552|ICD9CM|AB|164.0|Malignant neopl thymus
C0751560|ICD9CM|PT|146.0|Malignant neoplasm of tonsil
C0751560|ICD9CM|AB|146.0|Malignant neopl tonsil
C0751583|ICD9CM|PT|066.41|West Nile Fever with encephalitis
C0751583|ICD9CM|AB|066.41|West Nile Fever w/enceph
C0751674|ICD9CM|PT|516.4|Lymphangioleiomyomatosis
C0751674|ICD9CM|AB|516.4|Lymphangioleiomyomatosis
C0751758|ICD9CM|PT|327.32|Circadian rhythm sleep disorder, advanced sleep phase type
C0751758|ICD9CM|AB|327.32|Circadian rhy-advc sleep
C0751762|ICD9CM|PT|327.21|Primary central sleep apnea
C0751762|ICD9CM|AB|327.21|Prim central sleep apnea
C0751772|ICD9CM|PT|327.42|REM sleep behavior disorder
C0751772|ICD9CM|AB|327.42|REM sleep behavior dis
C0751774|ICD9CM|PT|327.51|Periodic limb movement disorder
C0751774|ICD9CM|AB|327.51|Periodic limb movement
C0751908|ICD9CM|AB|386.12|Vestibular neuronitis
C0751908|ICD9CM|PT|386.12|Vestibular neuronitis
C0751908|ICD9CM|AB|078.81|Epidemic vertigo
C0751908|ICD9CM|PT|078.81|Epidemic vertigo
C0751937|ICD9CM|AB|352.0|Olfactory nerve disorder
C0751937|ICD9CM|PT|352.0|Disorders of olfactory (1st) nerve
C0752150|ICD9CM|PT|339.81|Hypnic headache
C0752150|ICD9CM|AB|339.81|Hypnic headache
C0752294|ICD9CM|AB|307.46|Sleep arousal disorder
C0752294|ICD9CM|PT|307.46|Sleep arousal disorder
C0752295|ICD9CM|AB|327.41|Confusional arousals
C0752295|ICD9CM|PT|327.41|Confusional arousals
C0752304|ICD9CM|HT|768.7|Hypoxic-ischemic encephalopathy (HIE)
C0752304|ICD9CM|AB|768.70|Hypoxc-ischem enceph NOS
C0752304|ICD9CM|PT|768.70|Hypoxic-ischemic encephalopathy, unspecified
C0752347|ICD9CM|PT|331.82|Dementia with lewy bodies
C0752347|ICD9CM|AB|331.82|Dementia w Lewy bodies
C0795685|ICD9CM|PT|349.2|Disorders of meninges, not elsewhere classified
C0795685|ICD9CM|AB|349.2|Disorder of meninges NEC
C0795686|ICD9CM|PT|321.3|Meningitis due to trypanosomiasis
C0795686|ICD9CM|AB|321.3|Trypanosomiasis meningit
C0795690|ICD9CM|PT|756.72|Omphalocele
C0795690|ICD9CM|AB|756.72|Omphalocele
C0795698|ICD9CM|PT|053.29|Herpes zoster with other ophthalmic complications
C0795698|ICD9CM|AB|053.29|Herpes zoster of eye NEC
C0795699|MTH|PN|NOCODE|Other diseases of pharynx, NEC in ICD9CM
C0795699|ICD9CM|HT|478.2|Other diseases of pharynx, not elsewhere classified
C0795699|ICD9CM|PT|478.29|Other diseases of pharynx, not elsewhere classified
C0795699|ICD9CM|AB|478.29|Disease of pharynx NEC
C0795702|ICD9CM|PT|383.00|Acute mastoiditis without complications
C0795702|ICD9CM|AB|383.00|Ac mastoiditis w/o compl
C0795772|ICD9CM|PT|36.31|Open chest transmyocardial revascularization
C0795772|ICD9CM|AB|36.31|Open chest trans revasc
C0795773|ICD9CM|PT|36.32|Other transmyocardial revascularization
C0795773|ICD9CM|AB|36.32|Oth transmyo revascular
C0795774|ICD9CM|AB|37.35|Partial ventriculectomy
C0795774|ICD9CM|PT|37.35|Partial ventriculectomy
C0795775|ICD9CM|PT|37.67|Implantation of cardiomyostimulation system
C0795775|ICD9CM|AB|37.67|Imp cardiomyostimul sys
C0795778|ICD9CM|PT|86.67|Dermal regenerative graft
C0795778|ICD9CM|AB|86.67|Dermal regener graft
C0795779|ICD9CM|PT|92.31|Single source photon radiosurgery
C0795779|ICD9CM|AB|92.31|Sing source radiosurgery
C0795780|ICD9CM|PT|92.32|Multi-source photon radiosurgery
C0795780|ICD9CM|AB|92.32|Multisource radiosurgery
C0795781|ICD9CM|AB|92.33|Particulate radiosurgery
C0795781|ICD9CM|PT|92.33|Particulate radiosurgery
C0795782|ICD9CM|PT|92.39|Stereotactic radiosurgery, not elsewhere classified
C0795782|ICD9CM|AB|92.39|Stereo radiosurgery NEC
C0795783|ICD9CM|PT|96.29|Reduction of intussusception of alimentary tract
C0795783|ICD9CM|AB|96.29|Reduct intuss ali tract
C0795784|ICD9CM|PT|99.10|Injection or infusion of thrombolytic agent
C0795784|ICD9CM|AB|99.10|Inject/inf thrombo agent
C0795785|ICD9CM|PT|99.20|Injection or infusion of platelet inhibitor
C0795785|ICD9CM|AB|99.20|Inj/inf platelet inhibit
C0795786|ICD9CM|PT|V61.22|Counseling for perpetrator of spousal and partner abuse
C0795786|ICD9CM|PT|V61.12|Counseling for perpetrator of spousal and partner abuse
C0795786|ICD9CM|AB|V61.12|Cnsl perp partner abuse
C0795786|ICD9CM|AB|V61.22|Cnsl perp parent chld ab
C0812420|MTH|PN|NOCODE|Shock due to anesthesia, NEC in ICD9CM_2014
C0812420|ICD9CM|AB|995.4|Shock due to anesthesia
C0812420|ICD9CM|PT|995.4|Shock due to anesthesia, not elsewhere classified
C0812427|ICD9CM|AB|84.12|Amputation through foot
C0812427|ICD9CM|PT|84.12|Amputation through foot
C0812429|ICD9CM|PT|303.00|Acute alcoholic intoxication in alcoholism, unspecified
C0812429|ICD9CM|AB|303.00|Ac alcohol intox-unspec
C0812450|ICD9CM|AB|69.7|Insertion of iud
C0812450|ICD9CM|PT|69.7|Insertion of intrauterine contraceptive device
C0813173|ICD9CM|PT|295.40|Schizophreniform disorder, unspecified
C0813173|ICD9CM|AB|295.40|Schizophreniform dis NOS
C0815336|ICD9CM|PT|646.13|Edema or excessive weight gain in pregnancy, without mention of hypertension, antepartum condition or complication
C0815336|ICD9CM|AB|646.13|Edema in preg-antepartum
C0836917|ICD9CM|PT|767.0|Subdural and cerebral hemorrhage
C0836917|ICD9CM|AB|767.0|Cerebral hem at birth
C0837133|ICD9CM|PT|414.00|Coronary atherosclerosis of unspecified type of vessel, native or graft
C0837133|ICD9CM|AB|414.00|Cor ath unsp vsl ntv/gft
C0837134|ICD9CM|PT|414.01|Coronary atherosclerosis of native coronary artery
C0837134|ICD9CM|AB|414.01|Crnry athrscl natve vssl
C0837135|ICD9CM|PT|414.02|Coronary atherosclerosis of autologous vein bypass graft
C0837135|ICD9CM|AB|414.02|Crn ath atlg vn bps grft
C0837136|ICD9CM|PT|414.03|Coronary atherosclerosis of nonautologous biological bypass graft
C0837136|ICD9CM|AB|414.03|Crn ath nonatlg blg grft
C0837158|ICD9CM|PT|306.50|Psychogenic genitourinary malfunction, unspecified
C0837158|ICD9CM|AB|306.50|Psychogenic gu dis NOS
C0837418|ICD9CM|PT|711.39|Postdysenteric arthropathy, multiple sites
C0837418|ICD9CM|AB|711.39|Dysenter arthrit-mult
C0837419|ICD9CM|PT|711.31|Postdysenteric arthropathy, shoulder region
C0837419|ICD9CM|AB|711.31|Dysenter arthrit-shlder
C0837420|ICD9CM|PT|711.32|Postdysenteric arthropathy, upper arm
C0837420|ICD9CM|AB|711.32|Dysenter arthrit-up/arm
C0837421|ICD9CM|PT|711.33|Postdysenteric arthropathy, forearm
C0837421|ICD9CM|AB|711.33|Dysenter arthrit-forearm
C0837422|ICD9CM|PT|711.34|Postdysenteric arthropathy, hand
C0837422|ICD9CM|AB|711.34|Dysenter arthrit-hand
C0837423|ICD9CM|PT|711.35|Postdysenteric arthropathy, pelvic region and thigh
C0837423|ICD9CM|AB|711.35|Dysenter arthrit-pelvis
C0837424|ICD9CM|PT|711.36|Postdysenteric arthropathy, lower leg
C0837424|ICD9CM|AB|711.36|Dysenter arthrit-l/leg
C0837425|ICD9CM|PT|711.37|Postdysenteric arthropathy, ankle and foot
C0837425|ICD9CM|AB|711.37|Dysenter arthrit-ankle
C0837691|ICD9CM|PT|714.30|Polyarticular juvenile rheumatoid arthritis, chronic or unspecified
C0837691|ICD9CM|AB|714.30|Juv rheum arthritis NOS
C0837881|ICD9CM|PT|712.89|Other specified crystal arthropathies, multiple sites
C0837881|ICD9CM|AB|712.89|Cryst arthrop NEC-mult
C0837882|ICD9CM|PT|712.81|Other specified crystal arthropathies, shoulder region
C0837882|ICD9CM|AB|712.81|Cryst arthrop NEC-shlder
C0837883|ICD9CM|PT|712.82|Other specified crystal arthropathies, upper arm
C0837883|ICD9CM|AB|712.82|Cryst arthrop NEC-up/arm
C0837884|ICD9CM|PT|712.83|Other specified crystal arthropathies, forearm
C0837884|ICD9CM|AB|712.83|Crys arthrop NEC-forearm
C0837885|ICD9CM|PT|712.84|Other specified crystal arthropathies, hand
C0837885|ICD9CM|AB|712.84|Cryst arthrop NEC-hand
C0837886|ICD9CM|PT|712.85|Other specified crystal arthropathies, pelvic region and thigh
C0837886|ICD9CM|AB|712.85|Cryst arthrop NEC-pelvis
C0837887|ICD9CM|PT|712.86|Other specified crystal arthropathies, lower leg
C0837887|ICD9CM|AB|712.86|Cryst arthrop NEC-l/leg
C0837888|ICD9CM|PT|712.87|Other specified crystal arthropathies, ankle and foot
C0837888|ICD9CM|AB|712.87|Cryst arthrop NEC-ankle
C0837909|ICD9CM|PT|719.29|Villonodular synovitis, multiple sites
C0837909|ICD9CM|AB|719.29|Villonod synovit-mult jt
C0838222|ICD9CM|PT|719.41|Pain in joint, shoulder region
C0838222|ICD9CM|AB|719.41|Joint pain-shlder
C0838223|ICD9CM|PT|719.42|Pain in joint, upper arm
C0838223|ICD9CM|AB|719.42|Joint pain-up/arm
C0838224|ICD9CM|PT|719.43|Pain in joint, forearm
C0838224|ICD9CM|AB|719.43|Joint pain-forearm
C0838226|ICD9CM|PT|719.45|Pain in joint, pelvic region and thigh
C0838226|ICD9CM|AB|719.45|Joint pain-pelvis
C0838227|ICD9CM|PT|719.46|Pain in joint, lower leg
C0838227|ICD9CM|AB|719.46|Joint pain-l/leg
C0840764|ICD9CM|PT|911.8|Other and unspecified superficial injury of trunk, without mention of infection
C0840764|ICD9CM|AB|911.8|Superfic inj trunk NEC
C0840791|ICD9CM|PT|942.02|Burn of unspecified degree of chest wall, excluding breast and nipple
C0840791|ICD9CM|AB|942.02|Burn NOS chest wall
C0840795|ICD9CM|PT|942.10|Erythema [first degree] of trunk, unspecified site
C0840795|ICD9CM|AB|942.10|1st deg burn trunk NOS
C0840797|ICD9CM|PT|942.13|Erythema [first degree] of abdominal wall
C0840797|ICD9CM|AB|942.13|1st deg burn abdomn wall
C0840798|ICD9CM|PT|942.14|Erythema [first degree] of back [any part]
C0840798|ICD9CM|AB|942.14|1st deg burn back
C0840801|ICD9CM|PT|942.20|Blisters, epidermal loss [second degree] of trunk, unspecified site
C0840801|ICD9CM|AB|942.20|2nd deg burn trunk NOS
C0840802|ICD9CM|PT|942.21|Blisters, epidermal loss [second degree] of breast
C0840802|ICD9CM|AB|942.21|2nd deg burn breast
C0840804|ICD9CM|PT|942.23|Blisters, epidermal loss [second degree] of abdominal wall
C0840804|ICD9CM|AB|942.23|2nd deg burn abdomn wall
C0840805|ICD9CM|PT|942.24|Blisters, epidermal loss [second degree] of back [any part]
C0840805|ICD9CM|AB|942.24|2nd deg burn back
C0840808|ICD9CM|PT|942.30|Full-thickness skin loss [third degree, not otherwise specified] of trunk, unspecified site
C0840808|ICD9CM|AB|942.30|3rd deg burn trunk NOS
C0840810|ICD9CM|PT|942.34|Full-thickness skin loss [third degree,not otherwise specified] of back [any part]
C0840810|ICD9CM|AB|942.34|3rd deg burn back
C0840880|ICD9CM|PT|996.75|Other complications due to nervous system device, implant, and graft
C0840880|ICD9CM|AB|996.75|Comp-nerv sys dev/graft
C0840927|ICD9CM|PT|781.8|Neurologic neglect syndrome
C0840927|ICD9CM|AB|781.8|Neurologic neglect syndr
C0840982|ICD9CM|PT|E030|Unspecified activity
C0840982|ICD9CM|AB|E030|Activity NOS
C0840990|ICD9CM|AB|V02.62|Hepatitis C carrier
C0840990|ICD9CM|PT|V02.62|Hepatitis C carrier
C0841057|ICD9CM|HT|56.9|Other operations on ureter
C0841057|ICD9CM|PT|56.99|Other operations on ureter
C0841057|ICD9CM|AB|56.99|Ureteral operation NEC
C0841108|ICD9CM|HT|61.9|Other operations on scrotum and tunica vaginalis
C0841108|ICD9CM|PT|61.99|Other operations on scrotum and tunica vaginalis
C0841108|ICD9CM|AB|61.99|Scrotum & tunica op NEC
C0841133|ICD9CM|HT|64.9|Other operations on male genital organs
C0841133|ICD9CM|PT|64.99|Other operations on male genital organs
C0841133|ICD9CM|AB|64.99|Male genital op NEC
C0841595|ICD9CM|HT|99.5|Other vaccination and inoculation
C0841595|ICD9CM|PT|99.59|Other vaccination and inoculation
C0841595|ICD9CM|AB|99.59|Vaccination/innocula NEC
C0841706|ICD9CM|PT|14.79|Other operations on vitreous
C0841706|ICD9CM|AB|14.79|Vitreous operation NEC
C0841903|ICD9CM|PT|31.99|Other operations on trachea
C0841903|ICD9CM|AB|31.99|Other tracheal operation
C0841930|ICD9CM|HT|03.9|Other operations on spinal cord and spinal canal structures
C0841930|ICD9CM|PT|03.99|Other operations on spinal cord and spinal canal structures
C0841930|ICD9CM|AB|03.99|Spine canal struc op NEC
C0842094|ICD9CM|PT|41.98|Other operations on bone marrow
C0842094|ICD9CM|AB|41.98|Bone marrow ops NEC
C0842101|ICD9CM|PT|40.9|Other operations on lymphatic structures
C0842101|ICD9CM|AB|40.9|Lymph structure op NEC
C0842217|ICD9CM|HT|52.9|Other operations on pancreas
C0842217|ICD9CM|PT|52.99|Other operations on pancreas
C0842217|ICD9CM|AB|52.99|Pancreatic operation NEC
C0842378|ICD9CM|PT|99.73|Therapeutic erythrocytapheresis
C0842378|ICD9CM|AB|99.73|Therapeu erythropheresis
C0842626|ICD9CM|PT|07.11|Closed [percutaneous] [needle] biopsy of adrenal gland
C0842626|ICD9CM|AB|07.11|Closed adrenal gland bx
C0842627|ICD9CM|PT|51.12|Percutaneous biopsy of gallbladder or bile ducts
C0842627|ICD9CM|AB|51.12|Percu bx gb/bile duct
C0842628|ICD9CM|PT|54.24|Closed [percutaneous] [needle] biopsy of intra-abdominal mass
C0842628|ICD9CM|AB|54.24|Closed intra-abd mass bx
C0842630|ICD9CM|PT|60.13|Closed [percutaneous] biopsy of seminal vesicles
C0842630|ICD9CM|AB|60.13|Clos seminal vesicles bx
C0842631|ICD9CM|PT|26.11|Closed [needle] biopsy of salivary gland or duct
C0842631|ICD9CM|AB|26.11|Clos bx saliv gland/duct
C0842720|ICD9CM|HT|40.4|Radical excision of cervical lymph nodes
C0842950|ICD9CM|HT|17.1|Laparoscopic unilateral repair of inguinal hernia
C0842951|ICD9CM|HT|17.2|Laparoscopic bilateral repair of inguinal hernia
C0843081|ICD9CM|AB|48.75|Abdominal proctopexy
C0843081|ICD9CM|PT|48.75|Abdominal proctopexy
C0843593|ICD9CM|PT|68.51|Laparoscopically assisted vaginal hysterectomy (LAVH)
C0843593|ICD9CM|AB|68.51|Lap ast vag hysterectomy
C0843622|ICD9CM|AB|55.23|Closed renal biopsy
C0843622|ICD9CM|PT|55.23|Closed [percutaneous] [needle] biopsy of kidney
C0843999|ICD9CM|PT|37.95|Implantation of automatic cardioverter/defibrillator lead(s) only
C0843999|ICD9CM|AB|37.95|Implt cardiodefib leads
C0844429|ICD9CM|PT|31.95|Tracheoesophageal fistulization
C0844429|ICD9CM|AB|31.95|Tracheoesoph fistulizat
C0844519|ICD9CM|PT|11.0|Magnetic removal of embedded foreign body from cornea
C0844519|ICD9CM|AB|11.0|Magnet removal cornea FB
C0844541|ICD9CM|PT|13.3|Extracapsular extraction of lens by simple aspiration (and irrigation) technique
C0844541|ICD9CM|AB|13.3|Simpl aspir lens extract
C0844573|ICD9CM|PT|12.92|Injection into anterior chamber
C0844573|ICD9CM|AB|12.92|Anterior chamber inject
C0844969|ICD9CM|PT|08.36|Repair of blepharoptosis by other techniques
C0844969|ICD9CM|AB|08.36|Blepharoptos repair NEC
C0844977|ICD9CM|PT|08.42|Repair of entropion or ectropion by suture technique
C0844977|ICD9CM|AB|08.42|Suture entropion repair
C0844978|ICD9CM|PT|08.43|Repair of entropion or ectropion with wedge resection
C0844978|ICD9CM|AB|08.43|Wedg resec entropion rep
C0845085|ICD9CM|AB|81.28|Interphalangeal fusion
C0845085|ICD9CM|PT|81.28|Interphalangeal fusion
C0845973|ICD9CM|AB|95.14|X-ray study of eye
C0845973|ICD9CM|PT|95.14|X-ray study of eye
C0846208|ICD9CM|HT|26.9|Other operations on salivary gland or duct
C0846208|ICD9CM|PT|26.99|Other operations on salivary gland or duct
C0846208|ICD9CM|AB|26.99|Salivary operation NEC
C0846215|ICD9CM|PT|27.79|Other operations on uvula
C0846215|ICD9CM|AB|27.79|Other uvula operations
C0846218|ICD9CM|HT|28.9|Other operations on tonsils and adenoids
C0846218|ICD9CM|PT|28.99|Other operations on tonsils and adenoids
C0846218|ICD9CM|AB|28.99|Tonsil/adenoid ops NEC
C0846290|ICD9CM|HT|51.9|Other operations on biliary tract
C0846290|ICD9CM|PT|51.99|Other operations on biliary tract
C0846290|ICD9CM|AB|51.99|Biliary tract op NEC
C0846305|ICD9CM|PT|49.95|Control of (postoperative) hemorrhage of anus
C0846305|ICD9CM|AB|49.95|Control anal hemorrhage
C0846318|ICD9CM|PT|60.79|Other operations on seminal vesicles
C0846318|ICD9CM|AB|60.79|Seminal vesicle op NEC
C0846319|ICD9CM|PT|61.41|Suture of laceration of scrotum and tunica vaginalis
C0846319|ICD9CM|AB|61.41|Suture scrotal lacerat
C0846321|ICD9CM|PT|61.19|Other diagnostic procedures on scrotum and tunica vaginalis
C0846321|ICD9CM|AB|61.19|Scrot/tunica dx proc NEC
C0846357|ICD9CM|PT|73.8|Operations on fetus to facilitate delivery
C0846357|ICD9CM|AB|73.8|Fetal ops-facilitate del
C0846363|ICD9CM|PT|75.91|Evacuation of obstetrical incisional hematoma of perineum
C0846363|ICD9CM|AB|75.91|Evac ob inc hemat perin
C0846381|ICD9CM|HT|82.8|Other plastic operations on hand
C0846381|ICD9CM|PT|82.89|Other plastic operations on hand
C0846381|ICD9CM|AB|82.89|Hand plastic op NEC
C0846400|ICD9CM|PT|83.43|Excision of muscle or fascia for graft
C0846400|ICD9CM|AB|83.43|Musc/fasc excis for grft
C0846489|ICD9CM|AB|87.78|Ileal conduitogram
C0846489|ICD9CM|PT|87.78|Ileal conduitogram
C0846510|ICD9CM|PT|96.43|Digestive tract instillation, except gastric gavage
C0846510|ICD9CM|AB|96.43|GI tract instillat NEC
C0846521|ICD9CM|PT|96.45|Irrigation of nephrostomy and pyelostomy
C0846521|ICD9CM|AB|96.45|Nephrost/pyelost irrigat
C0846859|ICD9CM|PT|23.43|Insertion of removable bridge
C0846859|ICD9CM|AB|23.43|Insert removable bridge
C0847244|ICD9CM|AB|18.11|Otoscopy
C0847244|ICD9CM|PT|18.11|Otoscopy
C0848548|ICD9CM|HT|403.9|Hypertensive renal disease, unspecified
C0850128|ICD9CM|PT|V43.64|Hip joint replacement
C0850128|ICD9CM|AB|V43.64|Joint replaced hip
C0851140|ICD9CM|PT|233.1|Carcinoma in situ of cervix uteri
C0851140|ICD9CM|AB|233.1|Ca in situ cervix uteri
C0851225|ICD9CM|HT|228|Hemangioma and lymphangioma, any site
C0851252|ICD9CM|HT|72.5|Breech extraction
C0851258|ICD9CM|AB|726.65|Prepatellar bursitis
C0851258|ICD9CM|PT|726.65|Prepatellar bursitis
C0851311|ICD9CM|PT|V65.5|Person with feared complaint in whom no diagnosis was made
C0851311|ICD9CM|AB|V65.5|Persn w feared complaint
C0851314|ICD9CM|PT|E932.8|Antithyroid agents causing adverse effects in therapeutic use
C0851314|ICD9CM|AB|E932.8|Adv eff antithyroid agnt
C0851315|ICD9CM|PT|091.81|Acute syphilitic meningitis (secondary)
C0851315|ICD9CM|AB|091.81|Acute syphil meningitis
C0851323|ICD9CM|PT|E935.3|Salicylates causing adverse effects in therapeutic use
C0851323|ICD9CM|AB|E935.3|Adv eff salicylates
C0851324|ICD9CM|PT|E936.2|Succinimides causing adverse effects in therapeutic use
C0851324|ICD9CM|AB|E936.2|Adv eff succinimides
C0851325|ICD9CM|PT|E937.2|Paraldehyde causing adverse effects in therapeutic use
C0851325|ICD9CM|AB|E937.2|Adv eff paraldehyde
C0851326|ICD9CM|PT|E945.5|Expectorants causing adverse effects in therapeutic use
C0851326|ICD9CM|AB|E945.5|Adv eff expectorants
C0851327|ICD9CM|HT|E948|Bacterial vaccines causing adverse effects in therapeutic use
C0851328|ICD9CM|PT|E948.0|Bcg vaccine causing adverse effects in therapeutic use
C0851328|ICD9CM|AB|E948.0|Adv eff bcg vaccine
C0851329|ICD9CM|PT|E948.3|Plague vaccine causing adverse effects in therapeutic use
C0851329|ICD9CM|AB|E948.3|Adv eff plague vaccine
C0851330|ICD9CM|PT|E930.2|Chloramphenicol group causing adverse effects in therapeutic use
C0851330|ICD9CM|AB|E930.2|Adv eff chloramphenicol
C0851341|ICD9CM|AB|134.9|Infestation NOS
C0851341|ICD9CM|PT|134.9|Infestation, unspecified
C0854172|ICD9CM|PT|772.2|Subarachnoid hemorrhage of fetus or newborn
C0854172|ICD9CM|AB|772.2|NB subarachnoid hemorr
C0854248|ICD9CM|PT|482.83|Pneumonia due to other gram-negative bacteria
C0854248|ICD9CM|AB|482.83|Pneumo oth grm-neg bact
C0854530|ICD9CM|PT|058.81|Human herpesvirus 6 infection
C0854530|ICD9CM|AB|058.81|Human herpesvirus 6 infc
C0854802|ICD9CM|PT|204.12|Chronic lymphoid leukemia, in relapse
C0854802|ICD9CM|AB|204.12|Chr lymp leuk in relapse
C0856722|ICD9CM|PT|416.2|Chronic pulmonary embolism
C0856722|ICD9CM|AB|416.2|Chr pulmonary embolism
C0856761|ICD9CM|AB|453.0|Budd-chiari syndrome
C0856761|ICD9CM|PT|453.0|Budd-chiari syndrome
C0856825|ICD9CM|PT|279.51|Acute graft-versus-host disease
C0856825|ICD9CM|AB|279.51|Ac graft-versus-host dis
C0857751|ICD9CM|PT|695.11|Erythema multiforme minor
C0857751|ICD9CM|AB|695.11|Erythma multiforme minor
C0858895|ICD9CM|AB|112.85|Candidal enteritis
C0858895|ICD9CM|PT|112.85|Candidal enteritis
C0859058|ICD9CM|HT|253|Disorders of the pituitary gland and its hypothalamic control
C0859058|ICD9CM|PT|253.9|Unspecified disorder of the pituitary gland and its hypothalamic control
C0859058|ICD9CM|AB|253.9|Pituitary disorder NOS
C0859118|ICD9CM|PT|524.79|Other specified alveolar anomaly
C0859118|ICD9CM|AB|524.79|Oth spcf alveolar anmaly
C0859172|ICD9CM|HT|647|Infectious and parasitic conditions in the mother classifiable elsewhere, but complicating pregnancy, childbirth, or the puerperium
C0859268|ICD9CM|PT|864.15|Injury to liver with open wound into cavity, laceration, unspecified
C0859268|ICD9CM|AB|864.15|Liver lacerat unspcf opn
C0859273|ICD9CM|AB|952.9|Spinal cord injury NOS
C0859273|ICD9CM|PT|952.9|Unspecified site of spinal cord injury without evidence of spinal bone injury
C0859375|ICD9CM|PT|952.11|T1-T6 level with complete lesion of spinal cord
C0859375|ICD9CM|AB|952.11|Complete les cord/t1-t6
C0859376|ICD9CM|PT|952.12|T1-T6 level with anterior cord syndrome
C0859376|ICD9CM|AB|952.12|Anterior cord synd/t1-t6
C0859377|ICD9CM|PT|952.13|T1-T6 level with central cord syndrome
C0859377|ICD9CM|AB|952.13|Central cord synd/t1-t6
C0859378|ICD9CM|PT|952.14|T1-T6 level with other specified spinal cord injury
C0859378|ICD9CM|AB|952.14|T1-t6 spin cord inj NEC
C0859379|ICD9CM|PT|952.16|T7-T12 level with complete lesion of spinal cord
C0859379|ICD9CM|AB|952.16|Complete les cord/t7-t12
C0859380|ICD9CM|PT|952.17|T7-T12 level with anterior cord syndrome
C0859380|ICD9CM|AB|952.17|Anterior cord syn/t7-t12
C0859381|ICD9CM|PT|952.18|T7-T12 level with central cord syndrome
C0859381|ICD9CM|AB|952.18|Central cord syn/t7-t12
C0859643|ICD9CM|HT|290.2|Senile dementia with delusional or depressive features
C0859673|ICD9CM|PT|356.9|Unspecified hereditary and idiopathic peripheral neuropathy
C0859673|ICD9CM|AB|356.9|Idio periph neurpthy NOS
C0859693|ICD9CM|HT|805.0|Closed fracture of cervical vertebra without mention of spinal cord injury
C0859694|ICD9CM|HT|805.1|Open fracture of cervical vertebra without mention of spinal cord injury
C0859697|ICD9CM|PT|805.4|Closed fracture of lumbar vertebra without mention of spinal cord injury
C0859697|ICD9CM|AB|805.4|Fx lumbar vertebra-close
C0859698|ICD9CM|PT|805.5|Open fracture of lumbar vertebra without mention of spinal cord injury
C0859698|ICD9CM|AB|805.5|Fx lumbar vertebra-open
C0859703|ICD9CM|HT|806.0|Closed fracture of cervical vertebra with spinal cord injury
C0859704|ICD9CM|HT|806.1|Open fracture of cervical vertebra with spinal cord injury
C0859705|ICD9CM|HT|806.2|Closed fracture of dorsal vertebra with spinal cord injury
C0859706|ICD9CM|HT|806.3|Open fracture of dorsal vertebra with spinal cord injury
C0859760|ICD9CM|HT|974|Poisoning by water, mineral, and uric acid metabolism drugs
C0859814|ICD9CM|HT|516|Other alveolar and parietoalveolar pneumonopathy
C0859820|ICD9CM|HT|654.4|Other abnormalities in shape or position of gravid uterus and of neighboring structures
C0859825|ICD9CM|HT|760.7|Noxious influences affecting fetus or newborn via placenta or breast milk
C0859827|ICD9CM|PT|908.1|Late effect of internal injury to intra-abdominal organs
C0859827|ICD9CM|AB|908.1|Late eff int inj abdomen
C0859831|ICD9CM|PT|078.89|Other specified diseases due to viruses
C0859831|ICD9CM|AB|078.89|Oth spec dis viruses
C0859832|ICD9CM|PT|344.32|Monoplegia of lower limb affecting nondominant side
C0859832|ICD9CM|AB|344.32|Mnplg lwr lmb nondmnt sd
C0859851|ICD9CM|HT|943.5|Deep necrosis of underlying tissues due to burn [deep third degree] of upper limb, except wrist and hand, with loss of a body part
C0859855|ICD9CM|PT|995.61|Anaphylactic reaction due to peanuts
C0859855|ICD9CM|AB|995.61|Anphylct react peanuts
C0859856|ICD9CM|PT|995.62|Anaphylactic reaction due to crustaceans
C0859856|ICD9CM|AB|995.62|Anphylct react crstacns
C0859857|ICD9CM|PT|995.63|Anaphylactic reaction due to fruits and vegetables
C0859857|ICD9CM|AB|995.63|Anphylct react frts veg
C0859858|ICD9CM|PT|995.65|Anaphylactic reaction due to fish
C0859858|ICD9CM|AB|995.65|Anphylct reaction fish
C0859859|ICD9CM|PT|995.66|Anaphylactic reaction due to food additives
C0859859|ICD9CM|AB|995.66|Anphylct react food addv
C0859860|ICD9CM|PT|995.67|Anaphylactic reaction due to milk products
C0859860|ICD9CM|AB|995.67|Anphylct react milk prod
C0859861|ICD9CM|PT|995.68|Anaphylactic reaction due to eggs
C0859861|ICD9CM|AB|995.68|Anphylct reaction eggs
C0863239|ICD9CM|PT|02.39|Ventricular shunt to extracranial site NEC
C0863239|ICD9CM|AB|02.39|Vent shunt extracran NEC
C0864706|ICD9CM|PT|051.02|Vaccinia not from vaccination
C0864706|ICD9CM|AB|051.02|Vaccinia n/f vaccination
C0865240|ICD9CM|PT|284.81|Red cell aplasia (acquired)(adult)(with thymoma)
C0865240|ICD9CM|AB|284.81|Red cell aplasia
C0865505|ICD9CM|HT|V90|Retained foreign body
C0865505|ICD9CM|HT|V90-V90.99|RETAINED FOREIGN BODY
C0866710|ICD9CM|PT|735.1|Hallux varus (acquired)
C0866710|ICD9CM|AB|735.1|Hallux varus
C0867389|ICD9CM|PT|279.52|Chronic graft-versus-host disease
C0867389|ICD9CM|AB|279.52|Chronc graft-vs-host dis
C0868739|MTH|PN|NOCODE|Disorders of impulse control, NEC in ICD9CM_2014
C0868739|ICD9CM|HT|312.3|Disorders of impulse control, not elsewhere classified
C0868743|MTH|PN|NOCODE|Derangement of meniscus, NEC in ICD9CM_2014
C0868743|ICD9CM|AB|717.5|Derangement meniscus NEC
C0868743|ICD9CM|PT|717.5|Derangement of meniscus, not elsewhere classified
C0868752|MTH|PN|NOCODE|Muscular wasting and disuse atrophy, not elsewhere classified in ICD9CM
C0868752|ICD9CM|PT|728.2|Muscular wasting and disuse atrophy, not elsewhere classified
C0868752|ICD9CM|AB|728.2|Musc disuse atrophy NEC
C0868755|MTH|PN|NOCODE|Other complications of labor and delivery, not elsewhere classified in ICD9CM
C0868755|ICD9CM|HT|669|Other complications of labor and delivery, not elsewhere classified
C0868762|MTH|PN|NOCODE|Crushing injury of multiple sites, NEC in ICD9CM_2014
C0868762|ICD9CM|PT|929.0|Crushing injury of multiple sites, not elsewhere classified
C0868762|ICD9CM|AB|929.0|Crush inj mult site NEC
C0868767|MTH|PN|NOCODE|Posttraumatic wound infection NEC in ICD9CM_2014
C0868767|ICD9CM|PT|958.3|Posttraumatic wound infection not elsewhere classified
C0868767|ICD9CM|AB|958.3|Posttraum wnd infec NEC
C0868769|MTH|PN|NOCODE|Complications affecting specified body systems, NEC in ICD9CM_2014
C0868769|ICD9CM|HT|997|Complications affecting specified body systems, not elsewhere classified
C0868775|MTH|PN|NOCODE|Poisoning by aromatic analgesics, NEC in ICD9CM_2014
C0868775|ICD9CM|PT|965.4|Poisoning by aromatic analgesics, not elsewhere classified
C0868775|ICD9CM|AB|965.4|Pois-arom analgesics NEC
C0868777|ICD9CM|PT|307.42|Persistent disorder of initiating or maintaining sleep
C0868777|ICD9CM|AB|307.42|Persistent insomnia
C0868779|ICD9CM|PT|31.43|Closed [endoscopic] biopsy of larynx
C0868779|ICD9CM|AB|31.43|Closed biopsy larynx
C0868780|MTH|PN|NOCODE|Poisoning by mixed sedatives, NEC in ICD9CM_2014
C0868780|ICD9CM|AB|967.6|Poison-mix sedative NEC
C0868780|ICD9CM|PT|967.6|Poisoning by mixed sedatives, not elsewhere classified
C0868783|MTH|PN|NOCODE|Meningitis due to viruses NEC in ICD9CM_2014
C0868783|ICD9CM|PT|321.2|Meningitis due to viruses not elsewhere classified
C0868783|ICD9CM|AB|321.2|Mening in oth viral dis
C0868842|MTH|PN|NOCODE|Thoracic root lesions, NEC in ICD9CM_2014
C0868842|ICD9CM|PT|353.3|Thoracic root lesions, not elsewhere classified
C0868842|ICD9CM|AB|353.3|Thoracic root lesion NEC
C0868848|MTH|PN|NOCODE|Hereditary disturbances in tooth structure, NEC in ICD9CM_2014
C0868848|ICD9CM|PT|520.5|Hereditary disturbances in tooth structure, not elsewhere classified
C0868848|ICD9CM|AB|520.5|Heredit tooth struct NEC
C0868850|ICD9CM|AB|596.2|Vesical fistula NEC
C0868850|ICD9CM|PT|596.2|Vesical fistula, not elsewhere classified
C0868853|MTH|PN|NOCODE|Disorders of uterus, NEC in ICD9CM_2014
C0868853|ICD9CM|HT|621|Disorders of uterus, not elsewhere classified
C0868855|MTH|PN|NOCODE|Other and unspecified complications of the puerperium, NEC in ICD9CM
C0868855|ICD9CM|HT|674|Other and unspecified complications of the puerperium, not elsewhere classified
C0868862|ICD9CM|PT|720.2|Sacroiliitis, not elsewhere classified
C0868862|ICD9CM|AB|720.2|Sacroiliitis NEC
C0868867|ICD9CM|HT|E860|Accidental poisoning by alcohol, not elsewhere classified
C0868868|ICD9CM|PT|755.67|Anomalies of foot, not elsewhere classified
C0868868|ICD9CM|AB|755.67|Anomalies of foot NEC
C0868870|MTH|PN|NOCODE|Other lichen, NEC in ICD9CM
C0868870|ICD9CM|AB|697.8|Lichen NEC
C0868870|ICD9CM|PT|697.8|Other lichen, not elsewhere classified
C0868890|MTH|PN|NOCODE|Electrolyte and fluid disorders NEC in ICD9CM_2014
C0868890|ICD9CM|PT|276.9|Electrolyte and fluid disorders not elsewhere classified
C0868890|ICD9CM|AB|276.9|Electrolyt/fluid dis NEC
C0868892|MTH|PN|NOCODE|Depressive disorder, NEC in ICD9CM_2014
C0868892|ICD9CM|AB|311|Depressive disorder NEC
C0868892|ICD9CM|PT|311|Depressive disorder, not elsewhere classified
C0869062|ICD9CM|PT|719.80|Other specified disorders of joint, site unspecified
C0869062|ICD9CM|PT|716.80|Other specified arthropathy, site unspecified
C0869062|ICD9CM|AB|716.80|Arthropathy NEC-unspec
C0869062|ICD9CM|AB|719.80|Joint dis NEC-unspec
C0869063|ICD9CM|HT|718.8|Other joint derangement, not elsewhere classified
C0869063|ICD9CM|PT|718.80|Other joint derangement, not elsewhere classified, site unspecified
C0869063|ICD9CM|AB|718.80|Jt derangmnt NEC-unsp jt
C0869095|ICD9CM|PT|744.9|Unspecified congenital anomalies of face and neck
C0869095|ICD9CM|AB|744.9|Cong face/neck anom NOS
C0869098|ICD9CM|PT|995.7|Other adverse food reactions, not elsewhere classified
C0869098|ICD9CM|AB|995.7|Adverse food react NEC
C0869208|MTH|PN|NOCODE|Cervical root lesions, NEC in ICD9CM_2014
C0869208|ICD9CM|AB|353.2|Cervical root lesion NEC
C0869208|ICD9CM|PT|353.2|Cervical root lesions, not elsewhere classified
C0869240|ICD9CM|PT|941.05|Burn of unspecified degree of nose (septum)
C0869240|ICD9CM|AB|941.05|Burn NOS nose
C0869256|ICD9CM|PT|788.33|Mixed incontinence (male) (female)
C0869256|ICD9CM|AB|788.33|Mixed incontinence
C0869265|MTH|PN|NOCODE|Other complications of pregnancy, NEC in ICD9CM
C0869265|ICD9CM|HT|646|Other complications of pregnancy, not elsewhere classified
C0869267|ICD9CM|HT|E864|Accidental poisoning by corrosives and caustics, not elsewhere classified
C0869269|MTH|PN|NOCODE|Nonallopathic lesions, NEC in ICD9CM_2014
C0869269|ICD9CM|HT|739|Nonallopathic lesions, not elsewhere classified
C0869272|ICD9CM|HT|996-999.99|COMPLICATIONS OF SURGICAL AND MEDICAL CARE, NOT ELSEWHERE CLASSIFIED
C0869273|MTH|PN|NOCODE|Disturbance of conduct, NEC in ICD9CM_2014
C0869273|ICD9CM|HT|312|Disturbance of conduct, not elsewhere classified
C0869275|MTH|PN|NOCODE|Other diseases of mediastinum, NEC in ICD9CM
C0869275|ICD9CM|AB|519.3|Mediastinum disease NEC
C0869275|ICD9CM|PT|519.3|Other diseases of mediastinum, not elsewhere classified
C0869277|ICD9CM|PT|42.84|Repair of esophageal fistula, not elsewhere classified
C0869277|ICD9CM|AB|42.84|Esoph fistula repair NEC
C0869278|MTH|PN|NOCODE|Malignant neoplasm of spleen, NEC in ICD9CM_2014
C0869278|ICD9CM|PT|159.1|Malignant neoplasm of spleen, not elsewhere classified
C0869278|ICD9CM|AB|159.1|Malignant neo spleen NEC
C0869280|MTH|PN|NOCODE|Hematocele, female, NEC in ICD9CM_2014
C0869280|ICD9CM|AB|629.0|Hematocele, female NEC
C0869280|ICD9CM|PT|629.0|Hematocele, female, not elsewhere classified
C0869286|MTH|PN|NOCODE|Other complications of procedures, NEC in ICD9CM
C0869286|ICD9CM|HT|998|Other complications of procedures, NEC
C0869289|ICD9CM|PT|V62.81|Interpersonal problems, not elsewhere classified
C0869289|ICD9CM|AB|V62.81|Interpersonal probl NEC
C0869291|MTH|PN|NOCODE|Radiological examination, NEC in ICD9CM_2014
C0869291|ICD9CM|PT|V72.5|Radiological examination, not elsewhere classified
C0869291|ICD9CM|AB|V72.5|Radiological exam NEC
C0869292|MTH|PN|NOCODE|Other diseases of trachea and bronchus, NEC in ICD9CM
C0869292|ICD9CM|HT|519.1|Other diseases of trachea and bronchus, not elsewhere classified
C0869296|ICD9CM|PT|718.81|Other joint derangement, not elsewhere classified, shoulder region
C0869296|ICD9CM|AB|718.81|Jt derangment NEC-shlder
C0869298|ICD9CM|PT|718.82|Other joint derangement, not elsewhere classified, upper arm
C0869298|ICD9CM|AB|718.82|Jt derangment NEC-up/arm
C0869300|ICD9CM|PT|718.83|Other joint derangement, not elsewhere classified, forearm
C0869300|ICD9CM|AB|718.83|Jt derangmnt NEC-forearm
C0869419|ICD9CM|PT|746.84|Obstructive anomalies of heart, not elsewhere classified
C0869419|ICD9CM|AB|746.84|Obstruct heart anom NEC
C0869423|MTH|PN|NOCODE|Mineral deficiency, NEC in ICD9CM_2014
C0869423|ICD9CM|AB|269.3|Mineral deficiency NEC
C0869423|ICD9CM|PT|269.3|Mineral deficiency, not elsewhere classified
C0869426|ICD9CM|PT|718.84|Other joint derangement, not elsewhere classified, hand
C0869426|ICD9CM|AB|718.84|Jt derangement NEC-hand
C0869428|ICD9CM|PT|718.85|Other joint derangement, not elsewhere classified, pelvic region and thigh
C0869428|ICD9CM|AB|718.85|Jt derangment NEC-pelvis
C0869430|ICD9CM|PT|718.86|Other joint derangement, not elsewhere classified, lower leg
C0869430|ICD9CM|AB|718.86|Jt derangement NEC-l/leg
C0869432|ICD9CM|PT|718.87|Other joint derangement, not elsewhere classified, ankle and foot
C0869432|ICD9CM|AB|718.87|Jt derangement NEC-ankle
C0869434|ICD9CM|PT|718.88|Other joint derangement, not elsewhere classified, other specified sites
C0869434|ICD9CM|AB|718.88|Jt derangment NEC-oth jt
C0869436|ICD9CM|PT|718.89|Other joint derangement, not elsewhere classified, multiple sites
C0869436|ICD9CM|AB|718.89|Jt derangement NEC-mult
C0869438|MTH|PN|NOCODE|Other affections of shoulder region, NEC in ICD9CM
C0869438|ICD9CM|PT|726.2|Other affections of shoulder region, not elsewhere classified
C0869438|ICD9CM|AB|726.2|Shoulder region dis NEC
C0869440|MTH|PN|NOCODE|Poisoning by antidotes and chelating agents, NEC in ICD9CM_2014
C0869440|ICD9CM|PT|977.2|Poisoning by antidotes and chelating agents, not elsewhere classified
C0869440|ICD9CM|AB|977.2|Poisoning-antidotes NEC
C0869442|MTH|PN|NOCODE|Unspecified complication of procedure, NEC in ICD9CM_2014
C0869442|ICD9CM|PT|998.9|Unspecified complication of procedure, not elsewhere classified
C0869442|ICD9CM|AB|998.9|Surgical complicat NOS
C0869445|ICD9CM|PT|E852.5|Accidental poisoning by mixed sedatives, not elsewhere classified
C0869445|ICD9CM|AB|E852.5|Acc poison-mix sedtv NEC
C0869447|MTH|PN|NOCODE|Lumbosacral root lesions, NEC in ICD9CM_2014
C0869447|ICD9CM|PT|353.4|Lumbosacral root lesions, not elsewhere classified
C0869447|ICD9CM|AB|353.4|Lumbsacral root les NEC
C0869450|ICD9CM|HT|719.5|Stiffness of joint, not elsewhere classified
C0869452|MTH|PN|NOCODE|Other diseases of respiratory system, NEC in ICD9CM
C0869452|ICD9CM|PT|519.8|Other diseases of respiratory system, not elsewhere classified
C0869452|ICD9CM|AB|519.8|Resp system disease NEC
C0869474|ICD9CM|AB|315.1|Mathematics disorder
C0869474|ICD9CM|PT|315.1|Mathematics disorder
C0869476|MTH|PN|NOCODE|Revision of operative wound of anterior segment, NEC in ICD9CM_2014
C0869476|ICD9CM|PT|12.83|Revision of operative wound of anterior segment, not elsewhere classified
C0869476|ICD9CM|AB|12.83|Revis ant seg op wnd NEC
C0869477|MTH|PN|NOCODE|Removal of packing from trunk, NEC in ICD9CM_2014
C0869477|ICD9CM|PT|97.85|Removal of packing from trunk, not elsewhere classified
C0869477|ICD9CM|AB|97.85|Remov trunk packing NEC
C0869481|ICD9CM|HT|V65.4|Other counseling, not elsewhere classified
C0869483|MTH|PN|NOCODE|Other known or suspected fetal abnormality, NEC, affecting management of mother in ICD9CM
C0869483|ICD9CM|HT|655.8|Other known or suspected fetal abnormality, not elsewhere classified, affecting management of mother
C0869496|ICD9CM|PT|259.3|Ectopic hormone secretion, not elsewhere classified
C0869496|ICD9CM|AB|259.3|Ectopic hormone secr NEC
C0869499|MTH|PN|NOCODE|Delay in sexual development and puberty, NEC in ICD9CM_2014
C0869499|ICD9CM|AB|259.0|Delay sexual develop NEC
C0869499|ICD9CM|PT|259.0|Delay in sexual development and puberty, not elsewhere classified
C0869502|ICD9CM|PT|E933.4|Enzymes, not elsewhere classified, causing adverse effects in therapeutic use
C0869502|ICD9CM|AB|E933.4|Adv eff enzymes NEC
C0869504|ICD9CM|PT|E933.5|Vitamins, not elsewhere classified, causing adverse effects in therapeutic use
C0869504|ICD9CM|AB|E933.5|Adv eff vitamins NEC
C0869507|MTH|PN|NOCODE|Poisoning by enzymes, NEC in ICD9CM_2014
C0869507|ICD9CM|AB|963.4|Poisoning-enzymes NEC
C0869507|ICD9CM|PT|963.4|Poisoning by enzymes, not elsewhere classified
C0869511|MTH|PN|NOCODE|Poisoning by vitamins, NEC in ICD9CM_2014
C0869511|ICD9CM|AB|963.5|Poisoning-vitamins NEC
C0869511|ICD9CM|PT|963.5|Poisoning by vitamins, not elsewhere classified
C0869513|ICD9CM|PT|E850.4|Accidental poisoning by aromatic analgesics, not elsewhere classified
C0869513|ICD9CM|AB|E850.4|Acc poison-arom analgesc
C0869515|MTH|PN|NOCODE|Precocious sexual development and puberty, NEC in ICD9CM_2014
C0869515|ICD9CM|AB|259.1|Sexual precocity NEC
C0869515|ICD9CM|PT|259.1|Precocious sexual development and puberty, not elsewhere classified
C0869528|ICD9CM|HT|711.6|Arthropathy associated with mycoses
C0869528|ICD9CM|PT|711.60|Arthropathy associated with mycoses, site unspecified
C0869528|ICD9CM|AB|711.60|Mycotic arthritis-unspec
C0869904|ICD9CM|HT|72-75.99|OBSTETRICAL PROCEDURES
C0870073|ICD9CM|HT|28|Operations on tonsils and adenoids
C0876943|ICD9CM|PT|98.20|Removal of foreign body, not otherwise specified
C0876943|ICD9CM|AB|98.20|Removal of FB NOS
C0877176|ICD9CM|AB|038.12|MRSA septicemia
C0877176|ICD9CM|PT|038.12|Methicillin resistant Staphylococcus aureus septicemia
C0877208|ICD9CM|HT|674.5|Peripartum cardiomyopathy
C0877308|ICD9CM|AB|779.82|Neonatal tachycardia
C0877308|ICD9CM|PT|779.82|Neonatal tachycardia
C0877720|ICD9CM|PT|739.0|Nonallopathic lesions, head region
C0877720|ICD9CM|AB|739.0|Somat dys head region
C0877722|ICD9CM|PT|739.1|Nonallopathic lesions, cervical region
C0877722|ICD9CM|AB|739.1|Somat dysfunc cervic reg
C0877724|ICD9CM|PT|739.2|Nonallopathic lesions, thoracic region
C0877724|ICD9CM|AB|739.2|Somat dysfunc thorac reg
C0877726|ICD9CM|PT|739.3|Nonallopathic lesions, lumbar region
C0877726|ICD9CM|AB|739.3|Somat dysfunc lumbar reg
C0877728|ICD9CM|PT|739.4|Nonallopathic lesions, sacral region
C0877728|ICD9CM|AB|739.4|Somat dysfunc sacral reg
C0877730|ICD9CM|PT|739.5|Nonallopathic lesions, pelvic region
C0877730|ICD9CM|AB|739.5|Somat dysfunc pelvic reg
C0877732|ICD9CM|PT|739.6|Nonallopathic lesions, lower extremities
C0877732|ICD9CM|AB|739.6|Somat dysfunc lower extr
C0877734|ICD9CM|PT|739.7|Nonallopathic lesions, upper extremities
C0877734|ICD9CM|AB|739.7|Somat dysfunc upper extr
C0877736|ICD9CM|PT|739.8|Nonallopathic lesions, rib cage
C0877736|ICD9CM|AB|739.8|Somat dysfunc rib cage
C0877738|MTH|PN|NOCODE|Peripheral vascular complications, NEC in ICD9CM_2014
C0877738|ICD9CM|PT|997.2|Peripheral vascular complications, not elsewhere classified
C0877738|ICD9CM|AB|997.2|Surg comp-peri vasc syst
C0877771|MTH|PN|NOCODE|Angioneurotic edema, NEC in ICD9CM_2014
C0877771|ICD9CM|AB|995.1|Angioneurotic edema
C0877771|ICD9CM|PT|995.1|Angioneurotic edema, not elsewhere classified
C0877792|ICD9CM|HT|327.3|Circadian rhythm sleep disorder
C0877841|ICD9CM|HT|V15.0|Personal history of allergy, other than to medicinal agents, presenting hazards to health
C0877842|ICD9CM|HT|V26.2|Procreation management investigation and testing
C0877843|ICD9CM|PT|V76.49|Special screening for malignant neoplasms of other sites
C0877843|ICD9CM|HT|V76.4|Screening for malignant neoplasms of other sites
C0877843|ICD9CM|AB|V76.49|Screen mal neop oth site
C0877844|ICD9CM|HT|V76.8|Screening for other malignant neoplasms
C0877845|ICD9CM|PT|V77.99|Screening for other and unspecified endocrine, nutritional, metabolic, and immunity disorders
C0877845|ICD9CM|HT|V77.9|Screening for other and unspecified endocrine, nutritional, metabolic and immunity disorders
C0877845|ICD9CM|AB|V77.99|Screen-endoc/nut/met NEC
C0878514|ICD9CM|PT|35.84|Total correction of transposition of great vessels, not elsewhere classified
C0878514|ICD9CM|AB|35.84|Tot cor transpos grt ves
C0878518|ICD9CM|PT|E909.4|Tidalwave caused by earthquake
C0878518|ICD9CM|AB|E909.4|Acc d/t tidalwave NOS
C0878544|ICD9CM|HT|425|Cardiomyopathy
C0878688|ICD9CM|PT|082.49|Other ehrlichiosis
C0878688|ICD9CM|AB|082.49|Ehrlichiosis NEC
C0878691|ICD9CM|PT|294.10|Dementia in conditions classified elsewhere without behavioral disturbance
C0878691|ICD9CM|AB|294.10|Dementia w/o behav dist
C0878692|ICD9CM|PT|294.11|Dementia in conditions classified elsewhere with behavioral disturbance
C0878692|ICD9CM|AB|294.11|Dementia w behavior dist
C0878693|ICD9CM|AB|372.81|Conjunctivochalasis
C0878693|ICD9CM|PT|372.81|Conjunctivochalasis
C0878694|ICD9CM|PT|477.1|Allergic rhinitis due to food
C0878694|ICD9CM|AB|477.1|Allergic rhinitis-food
C0878695|ICD9CM|PT|494.0|Bronchiectasis without acute exacerbation
C0878695|ICD9CM|AB|494.0|Bronchiectas w/o ac exac
C0878696|ICD9CM|PT|494.1|Bronchiectasis with acute exacerbation
C0878696|ICD9CM|AB|494.1|Bronchiectasis w ac exac
C0878697|ICD9CM|HT|600.2|Benign localized hyperplasia of prostate
C0878700|ICD9CM|PT|707.10|Ulcer of lower limb, unspecified
C0878700|ICD9CM|AB|707.10|Ulcer of lower limb NOS
C0878701|ICD9CM|AB|707.11|Ulcer of thigh
C0878701|ICD9CM|PT|707.11|Ulcer of thigh
C0878702|ICD9CM|PT|707.14|Ulcer of heel and midfoot
C0878702|ICD9CM|AB|707.14|Ulcer of heel & midfoot
C0878703|ICD9CM|PT|707.15|Ulcer of other part of foot
C0878703|ICD9CM|AB|707.15|Ulcer other part of foot
C0878704|ICD9CM|PT|707.19|Ulcer of other part of lower limb
C0878704|ICD9CM|AB|707.19|Ulcer oth part low limb
C0878705|ICD9CM|AB|727.83|Plica syndrome
C0878705|ICD9CM|PT|727.83|Plica syndrome
C0878706|ICD9CM|PT|783.40|Lack of normal physiological development, unspecified
C0878706|ICD9CM|AB|783.40|Lack norm physio dev NOS
C0878707|ICD9CM|PT|790.01|Precipitous drop in hematocrit
C0878707|ICD9CM|AB|790.01|Drop, hematocrit, precip
C0878708|ICD9CM|PT|790.09|Other abnormality of red blood cells
C0878708|ICD9CM|AB|790.09|Abnormal RBC NEC
C0878709|ICD9CM|PT|792.5|Cloudy (hemodialysis) (peritoneal) dialysis effluent
C0878709|ICD9CM|AB|792.5|Cloudy dialysis effluent
C0878710|ICD9CM|PT|V15.02|Allergy to milk products
C0878710|ICD9CM|AB|V15.02|Hx-milk prod allergy
C0878711|ICD9CM|PT|V15.05|Allergy to other foods
C0878711|ICD9CM|AB|V15.05|Hx-other food allergy
C0878713|ICD9CM|PT|V15.08|Allergy to radiographic dye
C0878713|ICD9CM|AB|V15.08|Hx-radiogrphc dye allrgy
C0878714|ICD9CM|PT|V15.09|Other allergy, other than to medicinal agents
C0878714|ICD9CM|AB|V15.09|Hx-allergy NEC
C0878715|ICD9CM|HT|V21.3|Low birth weight status
C0878716|ICD9CM|PT|V21.30|Low birth weight status, unspecified
C0878716|ICD9CM|AB|V21.30|Low birthwt status NOS
C0878717|ICD9CM|PT|V21.31|Low birth weight status, less than 500 grams
C0878717|ICD9CM|AB|V21.31|Low birthwt status <500g
C0878718|ICD9CM|PT|V21.32|Low birth weight status, 500-999 grams
C0878718|ICD9CM|AB|V21.32|Low birthwt 500-999g
C0878719|ICD9CM|PT|V21.33|Low birth weight status, 1000-1499 grams
C0878719|ICD9CM|AB|V21.33|Low birthwt 1000-1499g
C0878720|ICD9CM|PT|V21.34|Low birth weight status, 1500-1999 grams
C0878720|ICD9CM|AB|V21.34|Low birthwt 1500-1999g
C0878721|ICD9CM|PT|V21.35|Low birth weight status, 2000-2500 grams
C0878721|ICD9CM|AB|V21.35|Low birthwt 2000-2500g
C0878722|ICD9CM|PT|V26.22|Aftercare following sterilization reversal
C0878722|ICD9CM|AB|V26.22|Sterilzation rev aftcare
C0878723|ICD9CM|PT|V26.29|Other investigation and testing
C0878723|ICD9CM|AB|V26.29|Investigate & test NEC
C0878725|ICD9CM|PT|V45.74|Acquired absence of organ, other parts of urinary tract
C0878725|ICD9CM|AB|V45.74|Acq absence urinary trct
C0878726|ICD9CM|PT|V45.75|Acquired absence of organ, stomach
C0878726|ICD9CM|AB|V45.75|Acq absence of stomach
C0878727|ICD9CM|PT|V45.76|Acquired absence of organ, lung
C0878727|ICD9CM|AB|V45.76|Acq absence of lung
C0878729|ICD9CM|HT|V49.8|Other specified conditions influencing health status
C0878729|ICD9CM|PT|V49.89|Other specified conditions influencing health status
C0878729|ICD9CM|AB|V49.89|Conditn influ health NEC
C0878730|ICD9CM|HT|V56.3|Encounter for adequacy testing for dialysis
C0878731|ICD9CM|PT|V56.31|Encounter for adequacy testing for hemodialysis
C0878731|ICD9CM|AB|V56.31|Hemodialysis testing
C0878732|ICD9CM|PT|V56.32|Encounter for adequacy testing for peritoneal dialysis
C0878732|ICD9CM|AB|V56.32|Peritoneal dialysis test
C0878734|ICD9CM|PT|V67.00|Follow-up examination, following surgery, unspecified
C0878734|ICD9CM|AB|V67.00|Follow-up surgery NOS
C0878735|ICD9CM|PT|V67.01|Following surgery, follow-up vaginal pap smear
C0878735|ICD9CM|AB|V67.01|Follow-up vag pap smear
C0878736|ICD9CM|PT|V67.09|Follow-up examination, following other surgery
C0878736|ICD9CM|AB|V67.09|Follow-up surgery NEC
C0878737|ICD9CM|PT|V71.81|Observation and evaluation for suspected abuse and neglect
C0878737|ICD9CM|AB|V71.81|Observe-abuse & neglect
C0878739|ICD9CM|PT|V76.47|Special screening for malignant neoplasms of vagina
C0878739|ICD9CM|AB|V76.47|Screen malig neop-vagina
C0878740|ICD9CM|HT|V76.5|Screening for malignant neoplasms of intestine
C0878741|ICD9CM|PT|V76.50|Special screening for malignant neoplasms for intestine, unspecified
C0878741|ICD9CM|AB|V76.50|Scrn malig neo-intes NOS
C0878742|ICD9CM|PT|V76.51|Special screening for malignant neoplasms of colon
C0878742|ICD9CM|AB|V76.51|Screen malig neop-colon
C0878746|ICD9CM|AB|E885.1|Fall from roller skates
C0878746|ICD9CM|PT|E885.1|Fall from roller skates
C0878747|ICD9CM|AB|E885.2|Fall from skateboard
C0878747|ICD9CM|PT|E885.2|Fall from skateboard
C0878748|ICD9CM|AB|E885.3|Fall from skis
C0878748|ICD9CM|PT|E885.3|Fall from skis
C0878749|ICD9CM|AB|E885.4|Fall from snowboard
C0878749|ICD9CM|PT|E885.4|Fall from snowboard
C0878750|ICD9CM|PT|E885.9|Fall from other slipping, tripping, or stumbling
C0878750|ICD9CM|AB|E885.9|Fall from slipping NEC
C0878751|ICD9CM|HT|645|Late pregnancy
C0878752|ICD9CM|HT|783.2|Abnormal loss of weight and underweight
C0878753|ICD9CM|HT|783.4|Lack of expected normal physiological development in childhood
C0878754|ICD9CM|HT|V26.3|Genetic counseling and testing on procreative management
C0878755|ICD9CM|HT|V49|Other conditions influencing health status
C0878756|ICD9CM|HT|E967|Perpetrator of child and adult abuse
C0878757|ICD9CM|PT|E967.0|Perpetrator of child and adult abuse, by father, stepfather, or boyfriend
C0878757|ICD9CM|AB|E967.0|Abuse by fther/stpfth/bf
C0878758|ICD9CM|PT|E967.2|Perpetrator of child and adult abuse, by mother, stepmother, or girlfriend
C0878758|ICD9CM|AB|E967.2|Abuse by mther/stpmth/gf
C0878773|ICD9CM|AB|596.51|Hypertonicity of bladder
C0878773|ICD9CM|PT|596.51|Hypertonicity of bladder
C0886366|MTH|PN|NOCODE|Encounter due to other acquired absence of organ NEC in ICD9CM
C0886366|ICD9CM|AB|V45.79|Acq absence of organ NEC
C0886366|ICD9CM|PT|V45.79|Other acquired absence of organ
C0886496|ICD9CM|AB|V26.21|Fertility testing
C0886496|ICD9CM|PT|V26.21|Fertility testing
C0917799|ICD9CM|AB|780.54|Hypersomnia NOS
C0917799|ICD9CM|PT|780.54|Hypersomnia, unspecified
C0917801|ICD9CM|AB|780.52|Insomnia NOS
C0917801|ICD9CM|PT|780.52|Insomnia, unspecified
C0917805|ICD9CM|HT|435|Transient cerebral ischemia
C0917805|ICD9CM|PT|435.9|Unspecified transient cerebral ischemia
C0917805|ICD9CM|AB|435.9|Trans cereb ischemia NOS
C0917918|ICD9CM|PT|V15.01|Allergy to peanuts
C0917918|ICD9CM|AB|V15.01|Hx-peanut allergy
C0917919|ICD9CM|PT|V15.03|Allergy to eggs
C0917919|ICD9CM|AB|V15.03|Hx-eggs allergy
C0917920|ICD9CM|PT|V15.04|Allergy to seafood
C0917920|ICD9CM|AB|V15.04|Hx-seafood allergy
C0917921|ICD9CM|PT|V15.07|Allergy to latex
C0917921|ICD9CM|AB|V15.07|Hx-latex allergy
C0917922|ICD9CM|AB|V45.78|Acquired absence of eye
C0917922|ICD9CM|PT|V45.78|Acquired absence of organ, eye
C0917967|ICD9CM|HT|379.4|Anomalies of pupillary function
C0917967|ICD9CM|PT|379.40|Abnormal pupillary function, unspecified
C0917967|ICD9CM|AB|379.40|Abn pupil function NOS
C0917981|ICD9CM|PT|335.21|Progressive muscular atrophy
C0917981|ICD9CM|AB|335.21|Prog muscular atrophy
C0919563|ICD9CM|PT|443.23|Dissection of renal artery
C0919563|ICD9CM|AB|443.23|Dissection renal artery
C0920028|ICD9CM|AB|208.92|Leukemia NOS in relapse
C0920028|ICD9CM|PT|208.92|Unspecified leukemia, in relapse
C0920049|ICD9CM|HT|567.3|Retroperitoneal infections
C0920296|ICD9CM|HT|315.0|Developmental reading disorder
C0920296|ICD9CM|AB|315.02|Developmental dyslexia
C0920296|ICD9CM|PT|315.02|Developmental dyslexia
C0920296|ICD9CM|AB|315.00|Reading disorder NOS
C0920296|ICD9CM|PT|315.00|Developmental reading disorder, unspecified
C0936215|ICD9CM|PT|266.1|Vitamin B6 deficiency
C0936215|ICD9CM|AB|266.1|Vitamin b6 deficiency
C0936250|ICD9CM|AB|054.0|Eczema herpeticum
C0936250|ICD9CM|PT|054.0|Eczema herpeticum
C0948343|ICD9CM|PT|518.7|Transfusion related acute lung injury (TRALI)
C0948343|ICD9CM|AB|518.7|Transfsn rel ac lung inj
C0948364|ICD9CM|PT|996.45|Peri-prosthetic osteolysis
C0948364|ICD9CM|AB|996.45|Periprosthetc osteolysis
C0949022|ICD9CM|PT|154.1|Malignant neoplasm of rectum
C0949022|ICD9CM|AB|154.1|Malignant neopl rectum
C0949122|ICD9CM|PT|464.00|Acute laryngitis without mention of obstruction
C0949122|ICD9CM|AB|464.00|Ac laryngitis w/o obst
C0949123|ICD9CM|PT|464.01|Acute laryngitis with obstruction
C0949123|ICD9CM|AB|464.01|Ac laryngitis w obstruct
C0949126|ICD9CM|PT|464.51|Supraglottitis unspecified, with obstruction
C0949126|ICD9CM|AB|464.51|Supraglottis w obstr NOS
C0949130|ICD9CM|PT|525.11|Loss of teeth due to trauma
C0949130|ICD9CM|AB|525.11|Loss of teeth d/t trauma
C0949131|ICD9CM|PT|525.12|Loss of teeth due to periodontal disease
C0949131|ICD9CM|AB|525.12|Loss teeth d/t peri dis
C0949132|ICD9CM|PT|525.13|Loss of teeth due to caries
C0949132|ICD9CM|AB|525.13|Loss of teeth d/t caries
C0949133|ICD9CM|PT|525.19|Other loss of teeth
C0949133|ICD9CM|AB|525.19|Loss of teeth NEC
C0949134|ICD9CM|PT|564.02|Outlet dysfunction constipation
C0949134|ICD9CM|AB|564.02|Outlet dysfnc constption
C0949135|ICD9CM|PT|564.09|Other constipation
C0949135|ICD9CM|AB|564.09|Constipation NEC
C0949136|ICD9CM|AB|602.3|Dysplasia of prostate
C0949136|ICD9CM|PT|602.3|Dysplasia of prostate
C0949138|ICD9CM|PT|733.93|Stress fracture of tibia or fibula
C0949138|ICD9CM|AB|733.93|Stress fx tibia/fibula
C0949139|ICD9CM|PT|733.94|Stress fracture of the metatarsals
C0949139|ICD9CM|AB|733.94|Stress fx metatarsals
C0949140|ICD9CM|PT|733.95|Stress fracture of other bone
C0949140|ICD9CM|AB|733.95|Stress fracture bone NEC
C0949141|ICD9CM|PT|772.10|Intraventricular hemorrhage unspecified grade
C0949141|ICD9CM|AB|772.10|NB intraven hem NOS
C0949142|ICD9CM|PT|772.11|Intraventricular hemorrhage, grade I
C0949142|ICD9CM|AB|772.11|NB intraven hem,grade i
C0949143|ICD9CM|PT|772.12|Intraventricular hemorrhage, grade II
C0949143|ICD9CM|AB|772.12|NB intraven hem,grade ii
C0949144|ICD9CM|PT|772.13|Intraventricular hemorrhage, grade III
C0949144|ICD9CM|AB|772.13|NB intravn hem,grade iii
C0949145|ICD9CM|PT|772.14|Intraventricular hemorrhage, grade IV
C0949145|ICD9CM|AB|772.14|NB intraven hem,grade iv
C0949146|ICD9CM|PT|793.80|Abnormal mammogram, unspecified
C0949146|ICD9CM|AB|793.80|Ab mammogram NOS
C0949148|ICD9CM|PT|793.89|Other (abnormal) findings on radiological examination of breast
C0949148|ICD9CM|AB|793.89|Abn finding-breast NEC
C0949149|ICD9CM|PT|840.7|Superior glenoid labrum lesion
C0949149|ICD9CM|AB|840.7|Sup glenoid labrm lesion
C0949150|ICD9CM|PT|997.71|Vascular complications of mesenteric artery
C0949150|ICD9CM|AB|997.71|Vasc comp mesenteric art
C0949151|ICD9CM|PT|997.72|Vascular complications of renal artery
C0949151|ICD9CM|AB|997.72|Vasc comp renal artery
C0949152|ICD9CM|HT|997.7|Vascular complications of other vessels
C0949152|ICD9CM|PT|997.79|Vascular complications of other vessels
C0949152|ICD9CM|AB|997.79|Vascular comp vessel NEC
C0949153|ICD9CM|PT|V10.53|Personal history of malignant neoplasm of renal pelvis
C0949153|ICD9CM|AB|V10.53|Hx malig renal pelvis
C0949155|ICD9CM|AB|V49.82|Dental sealant status
C0949155|ICD9CM|PT|V49.82|Dental sealant status
C0949156|ICD9CM|HT|V83|Genetic carrier status
C0949159|ICD9CM|PT|E888.0|Fall resulting in striking against sharp object
C0949159|ICD9CM|AB|E888.0|Fall striking sharp obj
C0949160|ICD9CM|PT|E888.1|Fall resulting in striking against other object
C0949160|ICD9CM|AB|E888.1|Fall striking object NEC
C0949161|ICD9CM|PT|E917.3|Striking against or struck accidentally by furniture without subsequent fall
C0949161|ICD9CM|AB|E917.3|Furnit w/o sub fall
C0949162|ICD9CM|PT|E917.4|Striking against or struck accidentally by other stationary object without subsequent fall
C0949162|ICD9CM|AB|E917.4|Stat ob w/o sub fall NEC
C0949163|ICD9CM|PT|E917.5|Striking against or struck accidentally by object in sports with subsequent fall
C0949163|ICD9CM|AB|E917.5|Sports acc w sub fall
C0949164|ICD9CM|PT|E917.6|Striking against or struck accidentally caused by a crowd, by collective fear or panic with subsequent fall
C0949164|ICD9CM|AB|E917.6|Crowd accidnt w sub fall
C0949165|ICD9CM|PT|E917.7|Striking against or struck accidentally by furniture with subsequent fall
C0949165|ICD9CM|AB|E917.7|Furniture acc w sub fall
C0949166|ICD9CM|PT|E917.8|Striking against or struck accidentally by other stationary object with subsequent fall
C0949166|ICD9CM|AB|E917.8|Stat obj w sub fall NEC
C0949167|ICD9CM|PT|411.81|Acute coronary occlusion without myocardial infarction
C0949167|ICD9CM|AB|411.81|Acute cor occlsn w/o MI
C0949168|ICD9CM|PT|V70.7|Examination of participant in clinical trial
C0949168|ICD9CM|AB|V70.7|Exam-clincal trial
C0949169|ICD9CM|PT|E917.0|Striking against or struck accidentally by objects or persons in sports
C0949169|ICD9CM|AB|E917.0|Sports acc w/o sub fall
C0949170|ICD9CM|PT|E917.1|Striking against or struck accidentally by a crowd, by collective fear or panic
C0949170|ICD9CM|AB|E917.1|Crowd w/o sub fall
C0949171|ICD9CM|PT|E917.2|Striking against or struck accidentally in running water
C0949171|ICD9CM|AB|E917.2|Run water w/o sub fall
C0949172|ICD9CM|PT|E917.9|Other accident caused by striking against or being struck accidentally by objects or persons
C0949172|ICD9CM|AB|E917.9|Obj w-w/o sub fall NEC
C0949744|ICD9CM|HT|93.6|Osteopathic manipulative treatment
C0994344|ICD9CM|AB|714.81|Rheumatoid lung
C0994344|ICD9CM|PT|714.81|Rheumatoid lung
C0994526|ICD9CM|PT|39.71|Endovascular implantation of other graft in abdominal aorta
C0994526|ICD9CM|AB|39.71|Endo imp oth grf abd aor
C0994528|ICD9CM|PT|41.04|Autologous hematopoietic stem cell transplant without purging
C0994528|ICD9CM|AB|41.04|Auto hem stem ct w/o pur
C0994529|ICD9CM|PT|41.05|Allogeneic hematopoietic stem cell transpant without purging
C0994529|ICD9CM|AB|41.05|Allo hem stem ct w/o pur
C0994530|ICD9CM|PT|41.07|Autologous hematopoietic stem cell transplant with purging
C0994530|ICD9CM|AB|41.07|Auto hem stem ct w purg
C0994531|ICD9CM|PT|60.97|Other transurethral destruction of prostate tissue by other thermotherapy
C0994531|ICD9CM|AB|60.97|Oth tu destr pros - rt
C0994532|ICD9CM|HT|86.5|Suture or other closure of skin and subcutaneous tissue
C0994533|ICD9CM|PT|86.59|Closure of skin and subcutaneous tissue of other sites
C0994533|ICD9CM|AB|86.59|Skin closure NEC
C0994534|ICD9CM|HT|99.7|Therapeutic apheresis or other injection, administration, or infusion of other therapeutic or prophylactic substance
C0994535|ICD9CM|PT|99.75|Administration of neuroprotective agent
C0994535|ICD9CM|AB|99.75|Adm neuroprotective agnt
C0994536|ICD9CM|PT|37.28|Intracardiac echocardiography
C0994536|ICD9CM|AB|37.28|Intracardiac echocardio
C0994537|ICD9CM|PT|44.32|Percutaneous [endoscopic] gastrojejunostomy
C0994537|ICD9CM|AB|44.32|Percu gastrojejunostomy
C0994538|ICD9CM|PT|67.51|Transabdominal cerclage of cervix
C0994538|ICD9CM|AB|67.51|Transab cerclage cervix
C0994539|ICD9CM|PT|67.59|Other repair of internal cervical os
C0994539|ICD9CM|AB|67.59|Oth rep int cervical os
C0994540|ICD9CM|AB|75.34|Other fetal monitoring
C0994540|ICD9CM|PT|75.34|Other fetal monitoring
C0994541|ICD9CM|AB|75.38|Fetal pulse oximetry
C0994541|ICD9CM|PT|75.38|Fetal pulse oximetry
C0994542|ICD9CM|PT|81.31|Refusion of atlas-axis spine
C0994542|ICD9CM|AB|81.31|Refusion of atlas-axis
C0994543|ICD9CM|PT|81.32|Refusion of other cervical spine, anterior column, anterior technique
C0994543|ICD9CM|AB|81.32|Refus oth cervcl ant/ant
C0994544|ICD9CM|PT|81.33|Refusion of other cervical spine, posterior column, posterior technique
C0994544|ICD9CM|AB|81.33|Refus oth cerv post/post
C0994545|ICD9CM|PT|81.34|Refusion of dorsal and dorsolumbar spine, anterior column, anterior technique
C0994545|ICD9CM|AB|81.34|Refus drs/drslmb ant/ant
C0994546|ICD9CM|PT|81.35|Refusion of dorsal and dorsolumbar spine, posterior column, posterior technique
C0994546|ICD9CM|AB|81.35|Refus drs/drslmb pst/pst
C0994547|ICD9CM|PT|81.38|Refusion of lumbar and lumbosacral spine, anterior column, posterior technique
C0994547|ICD9CM|AB|81.38|Refus lmb/lmbsc ant/post
C0994549|ICD9CM|PT|81.37|Refusion of lumbar and lumbosacral spine, posterior column, posterior technique
C0994549|ICD9CM|AB|81.37|Refus lmb/lmbsac pst/pst
C0994550|ICD9CM|PT|81.39|Refusion of spine, not elsewhere classified
C0994550|ICD9CM|AB|81.39|Refusion of spine NEC
C0994551|ICD9CM|PT|97.44|Nonoperative removal of heart assist system
C0994551|ICD9CM|AB|97.44|Nonop remov hrt asst sys
C0995154|ICD9CM|HT|338|Pain, not elsewhere classified
C1096116|ICD9CM|AB|286.52|Acquired hemophilia
C1096116|ICD9CM|PT|286.52|Acquired hemophilia
C1096624|ICD9CM|PT|789.05|Abdominal pain, periumbilic
C1096624|ICD9CM|AB|789.05|Abdmnal pain periumbilic
C1112318|ICD9CM|AB|779.84|Meconium staining
C1112318|ICD9CM|PT|779.84|Meconium staining
C1112452|ICD9CM|AB|055.1|Postmeasles pneumonia
C1112452|ICD9CM|PT|055.1|Postmeasles pneumonia
C1112488|ICD9CM|AB|779.81|Neonatal bradycardia
C1112488|ICD9CM|PT|779.81|Neonatal bradycardia
C1112529|ICD9CM|PT|944.14|Erythema [first degree] of two or more digits of hand including thumb
C1112529|ICD9CM|AB|944.14|1 deg burn fingr w thumb
C1112530|ICD9CM|PT|528.6|Leukoplakia of oral mucosa, including tongue
C1112530|ICD9CM|AB|528.6|Leukoplakia oral mucosa
C1112532|ICD9CM|PT|172.7|Malignant melanoma of skin of lower limb, including hip
C1112532|ICD9CM|AB|172.7|Malig melanoma leg
C1112533|ICD9CM|PT|172.6|Malignant melanoma of skin of upper limb, including shoulder
C1112533|ICD9CM|AB|172.6|Malig melanoma arm
C1112685|ICD9CM|PT|045.21|Acute nonparalytic poliomyelitis, poliovirus type I
C1112685|ICD9CM|AB|045.21|Nonparalyt polio-type 1
C1112686|ICD9CM|PT|045.22|Acute nonparalytic poliomyelitis, poliovirus type II
C1112686|ICD9CM|AB|045.22|Nonparalyt polio-type 2
C1112687|ICD9CM|PT|045.23|Acute nonparalytic poliomyelitis, poliovirus type III
C1112687|ICD9CM|AB|045.23|Nonparalyt polio-type 3
C1112690|ICD9CM|PT|366.01|Anterior subcapsular polar cataract
C1112690|ICD9CM|AB|366.01|Ant subcaps pol cataract
C1112691|ICD9CM|AB|440.32|Ath ext nonautlg bps gft
C1112691|ICD9CM|PT|440.32|Atherosclerosis of nonautologous biological bypass graft of the extremities
C1112693|ICD9CM|PT|345.01|Generalized nonconvulsive epilepsy, with intractable epilepsy
C1112693|ICD9CM|AB|345.01|Gen nonconv ep w intr ep
C1112700|ICD9CM|HT|099.4|Other nongonococcal urethritis [NGU]
C1112702|ICD9CM|AB|675.24|Mastitis-postpartum
C1112702|ICD9CM|PT|675.24|Nonpurulent mastitis associated with childbirth, postpartum condition or complication
C1112705|ICD9CM|AB|366.04|Nuclear cataract
C1112705|ICD9CM|PT|366.04|Nuclear cataract
C1112753|ICD9CM|HT|152|Malignant neoplasm of small intestine, including duodenum
C1112781|ICD9CM|PT|366.02|Posterior subcapsular polar cataract
C1112781|ICD9CM|AB|366.02|Post subcaps pol catarct
C1112782|ICD9CM|PT|172.5|Malignant melanoma of skin of trunk, except scrotum
C1112782|ICD9CM|AB|172.5|Malig melanoma trunk
C1112795|ICD9CM|PT|675.23|Nonpurulent mastitis associated with childbirth, antepartum condition or complication
C1112795|ICD9CM|AB|675.23|Mastitis-antepartum
C1135187|ICD9CM|PT|277.03|Cystic fibrosis with gastrointestinal manifestations
C1135187|ICD9CM|AB|277.03|Cystic fibrosis w GI man
C1135188|ICD9CM|PT|359.81|Critical illness myopathy
C1135188|ICD9CM|AB|359.81|Critical illness myopthy
C1135189|ICD9CM|AB|365.83|Aqueous misdirection
C1135189|ICD9CM|PT|365.83|Aqueous misdirection
C1135190|ICD9CM|PT|414.06|Coronary atherosclerosis of native coronary artery of transplanted heart
C1135190|ICD9CM|AB|414.06|Cor ath natv art tp hrt
C1135191|ICD9CM|HT|428.2|Systolic heart failure
C1135191|ICD9CM|PT|428.20|Systolic heart failure, unspecified
C1135191|ICD9CM|AB|428.20|Systolic hrt failure NOS
C1135194|ICD9CM|PT|428.22|Chronic systolic heart failure
C1135194|ICD9CM|AB|428.22|Chr systolic hrt failure
C1135196|ICD9CM|HT|428.3|Diastolic heart failure
C1135196|ICD9CM|PT|428.30|Diastolic heart failure, unspecified
C1135196|ICD9CM|AB|428.30|Diastolc hrt failure NOS
C1135206|ICD9CM|PT|438.6|Late effects of cerebrovascular disease, alterations of sensations
C1135206|ICD9CM|AB|438.6|Alteration of sensations
C1135207|ICD9CM|AB|438.84|Ataxia
C1135207|ICD9CM|PT|438.84|Other late effects of cerebrovascular disease, ataxia
C1135208|ICD9CM|AB|438.85|Vertigo
C1135208|ICD9CM|PT|438.85|Other late effects of cerebrovascular disease, vertigo
C1135209|ICD9CM|HT|443.2|Other arterial dissection
C1135210|ICD9CM|PT|443.29|Dissection of other artery
C1135210|ICD9CM|AB|443.29|Dissection artery NEC
C1135211|ICD9CM|HT|445.0|Atheroembolism Of extremities
C1135212|ICD9CM|PT|445.01|Atheroembolism of upper extremity
C1135212|ICD9CM|AB|445.01|Atheroembolism,upper ext
C1135213|ICD9CM|PT|445.02|Atheroembolism of lower extremity
C1135213|ICD9CM|AB|445.02|Atheroembolism,lower ext
C1135216|ICD9CM|PT|445.89|Atheroembolism of other site
C1135216|ICD9CM|HT|445.8|Atheroembolism of other sites
C1135216|ICD9CM|AB|445.89|Atheroembolism, site NEC
C1135217|ICD9CM|PT|454.8|Varicose veins of lower extremities with other complications
C1135217|ICD9CM|AB|454.8|Varic vein leg,comp NEC
C1135218|ICD9CM|PT|459.10|Postphlebetic syndrome without complications
C1135218|ICD9CM|AB|459.10|Postphlbtc synd w/o comp
C1135219|ICD9CM|PT|459.11|Postphlebetic syndrome with ulcer
C1135219|ICD9CM|AB|459.11|Postphlebtc synd w ulcer
C1135220|ICD9CM|PT|459.12|Postphlebetic syndrome with inflammation
C1135220|ICD9CM|AB|459.12|Postphlebtc syn w inflam
C1135221|ICD9CM|PT|459.13|Postphlebetic syndrome with ulcer and inflammation
C1135221|ICD9CM|AB|459.13|Postphl syn w ulc&inflam
C1135222|ICD9CM|PT|459.19|Postphlebetic syndrome with other complication
C1135222|ICD9CM|AB|459.19|Postphleb synd comp NEC
C1135223|ICD9CM|HT|459.3|Chronic venous hypertension (idiopathic)
C1135224|ICD9CM|PT|459.30|Chronic venous hypertension without complications
C1135224|ICD9CM|AB|459.30|Chr venous hypr w/o comp
C1135225|ICD9CM|PT|459.31|Chronic venous hypertension with ulcer
C1135225|ICD9CM|AB|459.31|Chr venous hyper w ulcer
C1135226|ICD9CM|PT|459.32|Chronic venous hypertension with inflammation
C1135226|ICD9CM|AB|459.32|Chr venous hypr w inflam
C1135227|ICD9CM|PT|459.33|Chronic venous hypertension with ulcer and inflammation
C1135227|ICD9CM|AB|459.33|Chr ven hyp w ulc&inflam
C1135228|ICD9CM|PT|459.39|Chronic venous hypertension with other complication
C1135228|ICD9CM|AB|459.39|Chr venous hyp comp NEC
C1135229|ICD9CM|PT|537.84|Dieulafoy lesion (hemorrhagic) of stomach and duodenum
C1135229|ICD9CM|AB|537.84|Dieulafoy les,stom&duod
C1135231|ICD9CM|PT|633.00|Abdominal pregnancy without intrauterine pregnancy
C1135231|ICD9CM|AB|633.00|Abd preg w/o intrau preg
C1135232|ICD9CM|PT|633.01|Abdominal pregnancy with intrauterine pregnancy
C1135232|ICD9CM|AB|633.01|Abd preg w intraut preg
C1135233|ICD9CM|PT|633.10|Tubal pregnancy without intrauterine pregnancy
C1135233|ICD9CM|AB|633.10|Tubal preg w/o intra prg
C1135234|ICD9CM|PT|633.11|Tubal pregnancy with intrauterine pregnancy
C1135234|ICD9CM|AB|633.11|Tubal preg w intra preg
C1135235|ICD9CM|PT|633.20|Ovarian pregnancy without intrauterine pregnancy
C1135235|ICD9CM|AB|633.20|Ovarn preg w/o intra prg
C1135236|ICD9CM|PT|633.21|Ovarian pregnancy with intrauterine pregnancy
C1135236|ICD9CM|AB|633.21|Ovarian preg w intra prg
C1135237|ICD9CM|PT|633.80|Other ectopic pregnancy without intrauterine pregnancy
C1135237|ICD9CM|AB|633.80|Ect preg NEC w/o int prg
C1135238|ICD9CM|PT|633.81|Other ectopic pregnancy with intrauterine pregnancy
C1135238|ICD9CM|AB|633.81|Ectpc prg NEC w int preg
C1135239|ICD9CM|PT|633.90|Unspecified ectopic pregnancy without intrauterine pregnancy
C1135239|ICD9CM|AB|633.90|Ect preg NOS w/o int prg
C1135240|ICD9CM|PT|633.91|Unspecified ectopic pregnancy with intrauterine pregnancy
C1135240|ICD9CM|AB|633.91|Ectp preg NOS w int preg
C1135241|ICD9CM|PT|765.20|Unspecified weeks of gestation
C1135241|ICD9CM|HT|765.2|Weeks of gestation
C1135241|ICD9CM|AB|765.20|Weeks of gestation NOS
C1135242|ICD9CM|PT|765.23|25-26 completed weeks of gestation
C1135242|ICD9CM|AB|765.23|25-26 comp wks gestation
C1135243|ICD9CM|PT|765.24|27-28 completed weeks of gestation
C1135243|ICD9CM|AB|765.24|27-28 comp wks gestation
C1135244|ICD9CM|PT|765.25|29-30 completed weeks of gestation
C1135244|ICD9CM|AB|765.25|29-30 comp wks gestation
C1135245|ICD9CM|PT|765.26|31-32 completed weeks of gestation
C1135245|ICD9CM|AB|765.26|31-32 comp wks gestation
C1135246|ICD9CM|PT|765.27|33-34 completed weeks of gestation
C1135246|ICD9CM|AB|765.27|33-34 comp wks gestation
C1135247|ICD9CM|PT|765.28|35-36 completed weeks of gestation
C1135247|ICD9CM|AB|765.28|35-36 comp wks gestation
C1135248|ICD9CM|PT|765.29|37 or more completed weeks of gestation
C1135248|ICD9CM|AB|765.29|37+ comp wks gestation
C1135250|ICD9CM|PT|770.89|Other respiratory problems after birth
C1135250|ICD9CM|AB|770.89|Resp prob after brth NEC
C1135251|ICD9CM|PT|771.81|Septicemia [sepsis] of newborn
C1135251|ICD9CM|AB|771.81|NB septicemia [sepsis]
C1135253|ICD9CM|AB|771.83|Bacteremia of newborn
C1135253|ICD9CM|PT|771.83|Bacteremia of newborn
C1135254|ICD9CM|PT|780.91|Fussy infant (baby)
C1135254|ICD9CM|AB|780.91|Fussy infant/baby
C1135260|ICD9CM|PT|795.31|Nonspecific positive findings for anthrax
C1135260|ICD9CM|AB|795.31|Nonsp postv find-anthrax
C1135261|ICD9CM|PT|795.39|Other nonspecific positive culture findings
C1135261|ICD9CM|AB|795.39|Nonsp positive cult NEC
C1135269|ICD9CM|AB|998.31|Disrup internal op wound
C1135269|ICD9CM|PT|998.31|Disruption of internal operation (surgical) wound
C1135270|ICD9CM|AB|998.32|Disrup-external op wound
C1135270|ICD9CM|PT|998.32|Disruption of external operation (surgical) wound
C1135271|ICD9CM|PT|V01.81|Contact with or exposure to anthrax
C1135271|ICD9CM|AB|V01.81|Contact/exposure-anthrax
C1135273|ICD9CM|PT|V13.21|Personal history of pre-term labor
C1135273|ICD9CM|AB|V13.21|History-pre-term labor
C1135275|ICD9CM|PT|V23.41|Pregnancy with history of pre-term labor
C1135275|ICD9CM|AB|V23.41|Preg w hx pre-term labor
C1135277|ICD9CM|HT|V54.1|Aftercare for healing traumatic fracture
C1135278|ICD9CM|PT|V54.10|Aftercare for healing traumatic fracture of arm, unspecified
C1135278|ICD9CM|AB|V54.10|Aftrcre traum fx arm NOS
C1135279|ICD9CM|PT|V54.11|Aftercare for healing traumatic fracture of upper arm
C1135279|ICD9CM|AB|V54.11|Aftrcare traum fx up arm
C1135280|ICD9CM|PT|V54.12|Aftercare for healing traumatic fracture of lower arm
C1135280|ICD9CM|AB|V54.12|Aftrcre traum fx low arm
C1135281|ICD9CM|PT|V54.13|Aftercare for healing traumatic fracture of hip
C1135281|ICD9CM|AB|V54.13|Aftrcre traumatic fx hip
C1135282|ICD9CM|PT|V54.14|Aftercare for healing traumatic fracture of leg, unspecified
C1135282|ICD9CM|AB|V54.14|Aftrcre traum fx leg NOS
C1135283|ICD9CM|PT|V54.15|Aftercare for healing traumatic fracture of upper leg
C1135283|ICD9CM|AB|V54.15|Aftrcare traum fx up leg
C1135284|ICD9CM|PT|V54.16|Aftercare for healing traumatic fracture of lower leg
C1135284|ICD9CM|AB|V54.16|Aftrcre traum fx low leg
C1135285|ICD9CM|PT|V54.17|Aftercare for healing traumatic fracture of vertebrae
C1135285|ICD9CM|AB|V54.17|Aftrcre traum fx vertebr
C1135286|ICD9CM|PT|V54.19|Aftercare for healing traumatic fracture of other bone
C1135286|ICD9CM|AB|V54.19|Aftrce traum fx bone NEC
C1135287|ICD9CM|HT|V54.2|Aftercare for healing pathologic fracture
C1135288|ICD9CM|PT|V54.20|Aftercare for healing pathologic fracture of arm, unspecified
C1135288|ICD9CM|AB|V54.20|Aftrcare path fx arm NOS
C1135289|ICD9CM|PT|V54.21|Aftercare for healing pathologic fracture of upper arm
C1135289|ICD9CM|AB|V54.21|Aftercare path fx up arm
C1135290|ICD9CM|PT|V54.22|Aftercare for healing pathologic fracture of lower arm
C1135290|ICD9CM|AB|V54.22|Aftrcare path fx low arm
C1135291|ICD9CM|PT|V54.23|Aftercare for healing pathologic fracture of hip
C1135291|ICD9CM|AB|V54.23|Aftercare path fx hip
C1135292|ICD9CM|PT|V54.24|Aftercare for healing pathologic fracture of leg, unspecified
C1135292|ICD9CM|AB|V54.24|Aftrcare path fx leg NOS
C1135293|ICD9CM|PT|V54.25|Aftercare for healing pathologic fracture of upper leg
C1135293|ICD9CM|AB|V54.25|Aftrcare path fx up leg
C1135294|ICD9CM|PT|V54.26|Aftercare for healing pathologic fracture of lower leg
C1135294|ICD9CM|AB|V54.26|Aftrcare path fx low leg
C1135295|ICD9CM|PT|V54.27|Aftercare for healing pathologic fracture of vertebrae
C1135295|ICD9CM|AB|V54.27|Aftrcare path fx vertebr
C1135296|ICD9CM|PT|V54.29|Aftercare for healing pathologic fracture of other bone
C1135296|ICD9CM|AB|V54.29|Aftrcre path fx bone NEC
C1135297|ICD9CM|PT|V54.81|Aftercare following joint replacement
C1135297|ICD9CM|AB|V54.81|Aftercare joint replace
C1135298|ICD9CM|PT|V58.42|Aftercare following surgery for neoplasm
C1135298|ICD9CM|AB|V58.42|Aftercare neoplasm surg
C1135299|ICD9CM|PT|V58.43|Aftercare following surgery for injury and trauma
C1135299|ICD9CM|AB|V58.43|Aftrcare inj/trauma surg
C1135300|ICD9CM|HT|V58.7|Aftercare following surgery to specified body systems, not elsewhere classified
C1135301|ICD9CM|PT|V58.71|Aftercare following surgery of the sense organs, NEC
C1135301|ICD9CM|AB|V58.71|Aft surg sense org NEC
C1135302|ICD9CM|PT|V58.72|Aftercare following surgery of the nervous system, NEC
C1135302|ICD9CM|AB|V58.72|Aftcre surg nerv sys NEC
C1135303|ICD9CM|PT|V58.73|Aftercare following surgery of the circulatory system, NEC
C1135303|ICD9CM|AB|V58.73|Aft surg circ syst NEC
C1135304|ICD9CM|PT|V58.74|Aftercare following surgery of the respiratory system, NEC
C1135304|ICD9CM|AB|V58.74|Aftrcre surg respsys NEC
C1135305|ICD9CM|PT|V58.75|Aftercare following surgery of the teeth, oral cavity and digestive system, NEC
C1135305|ICD9CM|AB|V58.75|Aft oral cav/dig sys NEC
C1135306|ICD9CM|PT|V58.76|Aftercare following surgery of the genitourinary system, NEC
C1135306|ICD9CM|AB|V58.76|Aftrcre surg GU syst NEC
C1135307|ICD9CM|PT|V58.77|Aftercare following surgery of the skin and subcutaneous tissue, NEC
C1135307|ICD9CM|AB|V58.77|Aft surg skin/subcu NEC
C1135308|ICD9CM|PT|V58.78|Aftercare following surgery of the musculoskeletal system, NEC
C1135308|ICD9CM|AB|V58.78|Aftrcre surg MS syst NEC
C1135309|ICD9CM|PT|V71.82|Observation and evaluation for suspected exposure to anthrax
C1135309|ICD9CM|AB|V71.82|Obs/eval sus exp anthrax
C1135310|ICD9CM|PT|V71.83|Observation and evaluation for suspected exposure to other biological agent
C1135310|ICD9CM|AB|V71.83|Obs/eval exp biol NEC
C1135312|ICD9CM|HT|V83.8|Other genetic carrier status
C1135312|ICD9CM|PT|V83.89|Other genetic carrier status
C1135312|ICD9CM|AB|V83.89|Genetic carrier stat NEC
C1135313|ICD9CM|PT|E885.0|Fall from (nonmotorized) scooter
C1135313|ICD9CM|AB|E885.0|Fall-nonmotor scooter
C1135314|ICD9CM|PT|E922.5|Accident caused by paintball gun
C1135314|ICD9CM|AB|E922.5|Accident-paintball gun
C1135315|ICD9CM|PT|E955.7|Suicide and self-inflicted injury by paintball gun
C1135315|ICD9CM|AB|E955.7|Self inj-paintball gun
C1135316|ICD9CM|PT|E979.0|Terrorism involving explosion of marine weapons
C1135316|ICD9CM|AB|E979.0|Terrorism,marine weapons
C1135317|ICD9CM|PT|E979.1|Terrorism involving destruction of aircraft
C1135317|ICD9CM|AB|E979.1|Terrorism,dest aircraft
C1135318|ICD9CM|PT|E979.2|Terrorism involving other explosions and fragments
C1135318|ICD9CM|AB|E979.2|Terrorism,explosions
C1135319|ICD9CM|PT|E979.3|Terrorism involving fires
C1135319|ICD9CM|AB|E979.3|Terrorism, fires
C1135320|ICD9CM|PT|E979.4|Terrorism involving firearms
C1135320|ICD9CM|AB|E979.4|Terrorism, firearms
C1135321|ICD9CM|PT|E979.5|Terrorism involving nuclear weapons
C1135321|ICD9CM|AB|E979.5|Terrorism, nuc weapons
C1135322|ICD9CM|PT|E979.6|Terrorism involving biological weapons
C1135322|ICD9CM|AB|E979.6|Terrorism, biologicals
C1135323|ICD9CM|PT|E979.7|Terrorism involving chemical weapons
C1135323|ICD9CM|AB|E979.7|Terrorism, chemicals
C1135324|ICD9CM|PT|E979.8|Terrorism involving other means
C1135324|ICD9CM|AB|E979.8|Terrorism, NEC/NOS
C1135325|ICD9CM|PT|E979.9|Terrorism secondary effects
C1135325|ICD9CM|AB|E979.9|Terrorism, secondary
C1135326|ICD9CM|PT|E985.7|Injury by paintball gun, undetermined whether accidental or purposely inflicted
C1135326|ICD9CM|AB|E985.7|Injury paintball gun NOS
C1135327|ICD9CM|PT|E999.1|Late effect of injury due to terrorism
C1135327|ICD9CM|AB|E999.1|Late effect, terrorism
C1135328|ICD9CM|PT|402.00|Malignant hypertensive heart disease without heart failure
C1135328|ICD9CM|AB|402.00|Mal hyp ht dis w/o hf
C1135329|ICD9CM|PT|402.01|Malignant hypertensive heart disease with heart failure
C1135329|ICD9CM|AB|402.01|Mal hypert hrt dis w hf
C1135330|ICD9CM|PT|402.10|Benign hypertensive heart disease without heart failure
C1135330|ICD9CM|AB|402.10|Benign hyp ht dis w/o hf
C1135331|ICD9CM|PT|402.11|Benign hypertensive heart disease with heart failure
C1135331|ICD9CM|AB|402.11|Benign hyp ht dis w hf
C1135332|ICD9CM|PT|402.90|Unspecified hypertensive heart disease without heart failure
C1135332|ICD9CM|AB|402.90|Hyp hrt dis NOS w/o hf
C1135333|ICD9CM|PT|402.91|Unspecified hypertensive heart disease with heart failure
C1135333|ICD9CM|AB|402.91|Hyp ht dis NOS w ht fail
C1135334|ICD9CM|HT|414.1|Aneurysm and dissection of heart
C1135335|ICD9CM|PT|454.9|Asymptomatic varicose veins
C1135335|ICD9CM|AB|454.9|Asympt varicose veins
C1135336|ICD9CM|PT|627.2|Symptomatic menopausal or female climacteric states
C1135336|ICD9CM|AB|627.2|Sympt fem climact state
C1135337|ICD9CM|PT|627.4|Symptomatic states associated with artificial menopause
C1135337|ICD9CM|AB|627.4|Sympt state w artif meno
C1135338|ICD9CM|PT|V49.81|Asymptomatic postmenopausal status (age-related) (natural)
C1135338|ICD9CM|AB|V49.81|Asympt postmeno status
C1135340|ICD9CM|HT|E999|Late effect of injury due to war operations and terrorism
C1135435|ICD9CM|HT|00|Procedures and interventions, Not Elsewhere Classified
C1135435|ICD9CM|HT|00-00.99|PROCEDURES AND INTERVENTIONS, NOT ELSEWHERE CLASSIFIED
C1135436|ICD9CM|PT|00.01|Therapeutic ultrasound of vessels of head and neck
C1135436|ICD9CM|AB|00.01|Ther ult head & neck ves
C1135437|ICD9CM|PT|00.02|Therapeutic ultrasound of heart
C1135437|ICD9CM|AB|00.02|Ther ultrasound of heart
C1135438|ICD9CM|PT|00.03|Therapeutic ultrasound of peripheral vascular vessels
C1135438|ICD9CM|AB|00.03|Ther ult peripheral ves
C1135439|ICD9CM|PT|00.09|Other therapeutic ultrasound
C1135439|ICD9CM|AB|00.09|Other therapeutic ultsnd
C1135440|ICD9CM|HT|00.1|Pharmaceuticals
C1135441|ICD9CM|PT|00.10|Implantation of chemotherapeutic agent
C1135441|ICD9CM|AB|00.10|Implant chemothera agent
C1135442|ICD9CM|PT|00.11|Infusion of drotrecogin alfa (activated)
C1135442|ICD9CM|AB|00.11|Infus drotrecogin alfa
C1135443|ICD9CM|PT|00.12|Administration of inhaled nitric oxide
C1135443|ICD9CM|AB|00.12|Adm inhal nitric oxide
C1135444|ICD9CM|PT|00.13|Injection or infusion of nesiritide
C1135444|ICD9CM|AB|00.13|Inject/infus nesiritide
C1135445|ICD9CM|PT|00.14|Injection or infusion of oxazolidinone class of antibiotics
C1135445|ICD9CM|AB|00.14|Injection oxazolidinone
C1135446|ICD9CM|PT|00.50|Implantation of cardiac resynchronization pacemaker without mention of defibrillation, total system [CRT-P]
C1135446|ICD9CM|AB|00.50|Impl CRT pacemaker sys
C1135447|ICD9CM|PT|00.51|Implantation of cardiac resynchronization defibrillator, total system [CRT-D]
C1135447|ICD9CM|AB|00.51|Impl CRT defibrillat sys
C1135448|ICD9CM|PT|00.52|Implantation or replacement of transvenous lead [electrode] into left ventricular coronary venous system
C1135448|ICD9CM|AB|00.52|Imp/rep lead lf ven sys
C1135449|ICD9CM|PT|00.53|Implantation or replacement of cardiac resynchronization pacemaker pulse generator only [CRT-P]
C1135449|ICD9CM|AB|00.53|Imp/rep CRT pacemakr gen
C1135450|ICD9CM|PT|00.54|Implantation or replacement of cardiac resynchronization defibrillator pulse generator only [CRT-D]
C1135450|ICD9CM|AB|00.54|Imp/rep CRT defib genat
C1135452|ICD9CM|PT|36.07|Insertion of drug-eluting coronary artery stent(s)
C1135452|ICD9CM|AB|36.07|Ins drug-elut coronry st
C1135454|ICD9CM|PT|49.75|Implantation or revision of artificial anal sphincter
C1135454|ICD9CM|AB|49.75|Impl or rev art anal sph
C1135455|ICD9CM|PT|49.76|Removal of artificial anal sphincter
C1135455|ICD9CM|AB|49.76|Remov art anal sphincter
C1135456|ICD9CM|HT|81.6|Other procedures on spine
C1135458|ICD9CM|HT|84.5|Implantation of other musculoskeletal devices and substances
C1135459|ICD9CM|PT|84.51|Insertion of interbody spinal fusion device
C1135459|ICD9CM|AB|84.51|Ins spinal fusion device
C1135460|ICD9CM|PT|84.52|Insertion of recombinant bone morphogenetic protein
C1135460|ICD9CM|AB|84.52|Insert recombinant BMP
C1135461|ICD9CM|PT|88.96|Other intraoperative magnetic resonance imaging
C1135461|ICD9CM|AB|88.96|Oth intraop mag res imag
C1135462|ICD9CM|PT|89.60|Continuous intra-arterial blood gas monitoring
C1135462|ICD9CM|AB|89.60|Cnt intraart bld gas mon
C1135463|ICD9CM|PT|99.77|Application or administration of an adhesion barrier substance
C1135463|ICD9CM|AB|99.77|App adhesion barrier sub
C1135976|ICD9CM|PT|41.06|Cord blood stem cell transplant
C1135976|ICD9CM|AB|41.06|Cord bld stem cell trans
C1137112|SRC|RHT|V-ICD9CM|ICD-9-CM
C1137112|SRC|RAB|V-ICD9CM|ICD9CM
C1137112|SRC|RPT|V-ICD9CM|International Classification of Diseases, Ninth Revision, Clinical Modification
C1137112|SRC|SSN|V-ICD9CM|International Classification of Diseases, Ninth Revision, Clinical Modification
C1140680|ICD9CM|PT|183.0|Malignant neoplasm of ovary
C1140680|ICD9CM|AB|183.0|Malign neopl ovary
C1142292|ICD9CM|AB|653.43|Fetopel disprop-antepart
C1142292|ICD9CM|PT|653.43|Fetopelvic disproportion, antepartum condition or complication
C1142293|ICD9CM|PT|653.40|Fetopelvic disproportion, unspecified as to episode of care or not applicable
C1142293|ICD9CM|AB|653.40|Fetopelv disprop-unspec
C1142536|ICD9CM|PT|482.42|Methicillin resistant pneumonia due to Staphylococcus aureus
C1142536|ICD9CM|AB|482.42|Meth res pneu d/t Staph
C1145628|ICD9CM|HT|337|Disorders of the autonomic nervous system
C1145628|ICD9CM|AB|337.9|Autonomic nerve dis NEC
C1145628|ICD9CM|PT|337.9|Unspecified disorder of autonomic nervous system
C1145757|ICD9CM|HT|718.7|Developmental dislocation of joint
C1146542|ICD9CM|HT|823.4|Torus fracture
C1168590|ICD9CM|HT|525.1|Loss of teeth due to trauma, extraction, or periodontal disease
C1175175|ICD9CM|PT|079.82|SARS-associated coronavirus
C1175175|ICD9CM|AB|079.82|SARS assoc coronavirus
C1176339|ICD9CM|PT|493.02|Extrinsic asthma with (acute) exacerbation
C1176339|ICD9CM|AB|493.02|Ext asthma w(acute) exac
C1176340|ICD9CM|PT|493.12|Intrinsic asthma with (acute) exacerbation
C1176340|ICD9CM|AB|493.12|Int asthma w (ac) exac
C1176341|ICD9CM|PT|493.22|Chronic obstructive asthma with (acute) exacerbation
C1176341|ICD9CM|AB|493.22|Ch obst asth w (ac) exac
C1176342|ICD9CM|PT|493.92|Asthma, unspecified type, with (acute) exacerbation
C1176342|ICD9CM|AB|493.92|Asthma NOS w (ac) exac
C1176343|ICD9CM|PT|645.10|Post term pregnancy, unspecified as to episode of care or not applicable
C1176343|ICD9CM|AB|645.10|Post term preg-unsp
C1176344|ICD9CM|PT|645.11|Post term pregnancy, delivered, with or without mention of antepartum condition
C1176344|ICD9CM|AB|645.11|Post term preg-del
C1176345|ICD9CM|PT|645.13|Post term pregnancy, antepartum condition or complication
C1176345|ICD9CM|AB|645.13|Post term preg-antepar
C1176346|ICD9CM|PT|645.20|Prolonged pregnancy, unspecified as to episode of care or not applicable
C1176346|ICD9CM|AB|645.20|Prolonged preg-unsp
C1176347|ICD9CM|PT|645.21|Prolonged pregnancy, delivered, with or without mention of antepartum condition
C1176347|ICD9CM|AB|645.21|Prolonged preg-del
C1176348|ICD9CM|PT|645.23|Prolonged pregnancy, antepartum condition or complication
C1176348|ICD9CM|AB|645.23|Prolonged preg-antepar
C1176349|ICD9CM|PT|718.70|Developmental dislocation of joint, site unspecified
C1176349|ICD9CM|AB|718.70|Dev dislocat jt site NOS
C1176350|ICD9CM|PT|718.71|Developmental dislocation of joint, shoulder region
C1176350|ICD9CM|AB|718.71|Dev dislocat joint-shldr
C1176351|ICD9CM|PT|718.72|Developmental dislocation of joint, upper arm
C1176351|ICD9CM|AB|718.72|Dev dislocat jt-up/arm
C1176352|ICD9CM|PT|718.73|Developmental dislocation of joint, forearm
C1176352|ICD9CM|AB|718.73|Dev dislocat jt-forearm
C1176353|ICD9CM|PT|718.74|Developmental dislocation of joint, hand
C1176353|ICD9CM|AB|718.74|Dev dislocat joint-hand
C1176354|ICD9CM|PT|718.75|Developmental dislocation of joint, pelvic region and thigh
C1176354|ICD9CM|AB|718.75|Dev dis jt-pelvic/thigh
C1176355|ICD9CM|PT|718.76|Developmental dislocation of joint, lower leg
C1176355|ICD9CM|AB|718.76|Dev disloc jt-lower leg
C1176356|ICD9CM|PT|718.77|Developmental dislocation of joint, ankle and foot
C1176356|ICD9CM|AB|718.77|Dev disloc jt-ankle/foot
C1176357|ICD9CM|PT|718.78|Developmental dislocation of joint, other specified sites
C1176357|ICD9CM|AB|718.78|Dev disloc jt-site NEC
C1176358|ICD9CM|PT|718.79|Developmental dislocation of joint, multiple sites
C1176358|ICD9CM|AB|718.79|Dev disloc jt-mult sites
C1176359|ICD9CM|PT|823.40|Torus fracture, tibia alone
C1176359|ICD9CM|AB|823.40|Torus fracture of tibia
C1176360|ICD9CM|PT|823.41|Torus fracture, fibula alone
C1176360|ICD9CM|AB|823.41|Torus fracture of fibula
C1176361|ICD9CM|PT|823.42|Torus fracture, fibula with tibia
C1176361|ICD9CM|AB|823.42|Torus fx tibia/fibula
C1253936|ICD9CM|HT|719.0|Effusion of joint
C1253936|ICD9CM|PT|719.00|Effusion of joint, site unspecified
C1253936|ICD9CM|AB|719.00|Joint effusion-unspec
C1254389|ICD9CM|AB|90.22|Culture-eye
C1254389|ICD9CM|PT|90.22|Microscopic examination of specimen from eye, culture
C1258666|ICD9CM|AB|727.43|Ganglion NOS
C1258666|ICD9CM|PT|727.43|Ganglion, unspecified
C1260368|ICD9CM|PT|00.15|High-dose infusion interleukin-2 [IL-2]
C1260368|ICD9CM|AB|00.15|High-dose infusion IL-2
C1260369|ICD9CM|HT|37.5|Heart replacement procedures
C1260376|ICD9CM|PT|37.54|Replacement or repair of other implantable component of (total) replacement heart system
C1260376|ICD9CM|AB|37.54|Repl/rep oth tot hrt sys
C1260379|ICD9CM|PT|68.31|Laparoscopic supracervical hysterectomy [LSH]
C1260379|ICD9CM|AB|68.31|Lap scervic hysterectomy
C1260381|ICD9CM|PT|81.62|Fusion or refusion of 2-3 vertebrae
C1260381|ICD9CM|AB|81.62|Fus/refus 2-3 vertebrae
C1260382|ICD9CM|PT|81.63|Fusion or refusion of 4-8 vertebrae
C1260382|ICD9CM|AB|81.63|Fus/refus 4-8 vertebrae
C1260383|ICD9CM|PT|81.64|Fusion or refusion of 9 or more vertebrae
C1260383|ICD9CM|AB|81.64|Fus/refus 9 vertebrae
C1260386|ICD9CM|PT|255.11|Glucocorticoid-remediable aldosteronism
C1260386|ICD9CM|AB|255.11|Glucrtcod-rem aldsternsm
C1260387|ICD9CM|PT|255.14|Other secondary aldosteronism
C1260387|ICD9CM|AB|255.14|Secondry aldosternsm NEC
C1260391|ICD9CM|PT|277.83|Iatrogenic carnitine deficiency
C1260391|ICD9CM|AB|277.83|Iatrogenic carnitine def
C1260392|ICD9CM|PT|277.84|Other secondary carnitine deficiency
C1260392|ICD9CM|AB|277.84|Sec carnitine defncy NEC
C1260393|ICD9CM|PT|282.41|Sickle-cell thalassemia without crisis
C1260393|ICD9CM|AB|282.41|Thlasema Hb-S w/o crisis
C1260398|ICD9CM|PT|282.64|Sickle-cell/Hb-C disease with crisis
C1260398|ICD9CM|AB|282.64|Hb-S/Hb-C dis w crisis
C1260401|ICD9CM|PT|282.68|Other sickle-cell disease without crisis
C1260401|ICD9CM|AB|282.68|Hb-S dis w/o crisis NEC
C1260402|ICD9CM|AB|289.52|Splenic sequestration
C1260402|ICD9CM|PT|289.52|Splenic sequestration
C1260404|ICD9CM|PT|289.81|Primary hypercoagulable state
C1260404|ICD9CM|AB|289.81|Prim hypercoagulable st
C1260406|ICD9CM|PT|331.19|Other frontotemporal dementia
C1260406|ICD9CM|AB|331.19|Frontotemp dementia NEC
C1260408|ICD9CM|AB|348.39|Encephalopathy NEC
C1260408|ICD9CM|PT|348.39|Other encephalopathy
C1260409|ICD9CM|PT|358.00|Myasthenia gravis without (acute) exacerbation
C1260409|ICD9CM|AB|358.00|Mysthna grvs w/o ac exac
C1260413|ICD9CM|PT|458.21|Hypotension of hemodialysis
C1260413|ICD9CM|AB|458.21|Hemododialysis hypotensn
C1260414|ICD9CM|PT|458.29|Other iatrogenic hypotension
C1260414|ICD9CM|AB|458.29|Iatrogenc hypotnsion NEC
C1260415|ICD9CM|PT|480.3|Pneumonia due to SARS-associated coronavirus
C1260415|ICD9CM|AB|480.3|Pneumonia due to SARS
C1260416|ICD9CM|HT|493.8|Other forms of asthma
C1260417|ICD9CM|PT|530.20|Ulcer of esophagus without bleeding
C1260417|ICD9CM|AB|530.20|Ulc esophagus w/o bleed
C1260419|ICD9CM|PT|600.01|Hypertrophy (benign) of prostate with urinary obstruction and other lower urinary tract symptoms (LUTS)
C1260419|ICD9CM|AB|600.01|BPH w urinary obs/LUTS
C1260421|ICD9CM|PT|600.10|Nodular prostate without urinary obstruction
C1260421|ICD9CM|AB|600.10|Nod prostate w/o ur obst
C1260422|ICD9CM|PT|600.11|Nodular prostate with urinary obstruction
C1260422|ICD9CM|AB|600.11|Nod prostate w ur obst
C1260424|ICD9CM|PT|600.21|Benign localized hyperplasia of prostate with urinary obstruction and other lower urinary tract symptoms (LUTS)
C1260424|ICD9CM|AB|600.21|BPH loc w urin obs/LUTS
C1260426|ICD9CM|PT|600.91|Hyperplasia of prostate, unspecified, with urinary obstruction and other lower urinary symptoms (LUTS)
C1260426|ICD9CM|AB|600.91|BPH NOS w ur obs/LUTS
C1260427|ICD9CM|PT|674.50|Peripartum cardiomyopathy, unspecified as to episode of care or not applicable
C1260427|ICD9CM|AB|674.50|Peripart cardiomy-unspec
C1260428|ICD9CM|PT|674.51|Peripartum cardiomyopathy, delivered, with or without mention of antepartum condition
C1260428|ICD9CM|AB|674.51|Peripartum cardiomy-del
C1260429|ICD9CM|PT|674.52|Peripartum cardiomyopathy, delivered, with mention of postpartum condition
C1260429|ICD9CM|AB|674.52|Peripart card del w p/p
C1260430|ICD9CM|PT|674.53|Peripartum cardiomyopathy, antepartum condition or complication
C1260430|ICD9CM|AB|674.53|Peripartum card-antepart
C1260431|ICD9CM|PT|674.54|Peripartum cardiomyopathy, postpartum condition or complication
C1260431|ICD9CM|AB|674.54|Peripartum card-postpart
C1260432|ICD9CM|AB|752.81|Scrotal transposition
C1260432|ICD9CM|PT|752.81|Scrotal transposition
C1260437|ICD9CM|PT|767.19|Other injuries to scalp
C1260437|ICD9CM|AB|767.19|Injuries to scalp NEC
C1260438|ICD9CM|PT|779.83|Delayed separation of umbilical cord
C1260438|ICD9CM|AB|779.83|Delay separate umbl cord
C1260443|ICD9CM|PT|790.29|Other abnormal glucose
C1260443|ICD9CM|AB|790.29|Abnormal glucose NEC
C1260444|ICD9CM|PT|850.11|Concussion, with loss of consciousness of 30 minutes or less
C1260444|ICD9CM|AB|850.11|Concus-brief coma <31 mn
C1260445|ICD9CM|PT|850.12|Concussion, with loss of consciousness from 31 to 59 minutes
C1260445|ICD9CM|AB|850.12|Concus-brf coma 31-59 mn
C1260446|ICD9CM|PT|959.12|Other injury of abdomen
C1260446|ICD9CM|AB|959.12|Injury of abdomen NEC
C1260447|ICD9CM|PT|959.13|Fracture of corpus cavernosum penis
C1260447|ICD9CM|AB|959.13|Fx corpus cavrnosm penis
C1260449|ICD9CM|PT|959.19|Other injury of other sites of trunk
C1260449|ICD9CM|AB|959.19|Trunk injury-sites NEC
C1260451|ICD9CM|AB|V01.82|Exposure to SARS
C1260451|ICD9CM|PT|V01.82|Exposure to SARS-associated coronavirus
C1260452|ICD9CM|PT|V04.81|Need for prophylactic vaccination and inoculation against influenza
C1260452|ICD9CM|AB|V04.81|Vaccin for influenza
C1260453|ICD9CM|PT|V04.82|Need for prophylactic vaccination and inoculation against respiratory syncytial virus (RSV)
C1260453|ICD9CM|AB|V04.82|Vaccination for RSV
C1260454|ICD9CM|HT|V04.8|Need for prophylactic vaccination and inoculation against other viral diseases
C1260454|ICD9CM|PT|V04.89|Need for prophylactic vaccination and inoculation against other viral diseases
C1260454|ICD9CM|AB|V04.89|Vaccn/inoc viral dis NEC
C1260455|ICD9CM|PT|V15.87|History of extracorporeal membrane oxygenation (ECMO)
C1260455|ICD9CM|AB|V15.87|Hx of ECMO
C1260457|ICD9CM|PT|V25.03|Encounter for emergency contraceptive counseling and prescription
C1260457|ICD9CM|AB|V25.03|Contracept mgmt-emergncy
C1260458|ICD9CM|PT|V43.22|Organ or tissue replaced by other means, fully implantable artificial heart
C1260458|ICD9CM|AB|V43.22|Artficial heart replace
C1260459|ICD9CM|AB|V45.85|Insulin pump status
C1260459|ICD9CM|PT|V45.85|Insulin pump status
C1260460|ICD9CM|PT|V53.91|Fitting and adjustment of insulin pump
C1260460|ICD9CM|AB|V53.91|Fit/adjust insulin pump
C1260461|ICD9CM|PT|V54.01|Encounter for removal of internal fixation device
C1260461|ICD9CM|AB|V54.01|Removal int fixation dev
C1260462|ICD9CM|PT|V54.02|Encounter for lengthening/adjustment of growth rod
C1260462|ICD9CM|AB|V54.02|Length/adjust growth rod
C1260463|ICD9CM|PT|V54.09|Other aftercare involving internal fixation device
C1260463|ICD9CM|AB|V54.09|Aftrcre int fixation dev
C1260466|ICD9CM|PT|V58.65|Long-term (current) use of steroids
C1260466|ICD9CM|AB|V58.65|Long-term use steroids
C1260467|ICD9CM|PT|V64.41|Laparoscopic surgical procedure converted to open procedure
C1260467|ICD9CM|AB|V64.41|Lap surg convert to open
C1260468|ICD9CM|PT|V64.42|Thoracoscopic surgical procedure converted to open procedure
C1260468|ICD9CM|AB|V64.42|Thoracoscop conv to open
C1260469|ICD9CM|PT|V64.43|Arthroscopic surgical procedure converted to open procedure
C1260469|ICD9CM|AB|V64.43|Arthroscopc conv to open
C1260471|ICD9CM|PT|V65.19|Other person consulting on behalf of another person
C1260471|ICD9CM|AB|V65.19|Person consult for anoth
C1260472|ICD9CM|PT|V65.46|Encounter for insulin pump training
C1260472|ICD9CM|AB|V65.46|Insulin pump training
C1260473|ICD9CM|PT|E928.4|External constriction caused by hair
C1260473|ICD9CM|AB|E928.4|Ext constriction-hair
C1260474|ICD9CM|PT|E928.5|External constriction caused by other object
C1260474|ICD9CM|AB|E928.5|Ext constriction-obj NEC
C1260673|ICD9CM|PT|282.69|Other sickle-cell disease with crisis
C1260673|ICD9CM|AB|282.69|Hb-SS dis NEC w crisis
C1260873|ICD9CM|AB|424.1|Aortic valve disorder
C1260873|ICD9CM|PT|424.1|Aortic valve disorders
C1260873|ICD9CM|HT|395|Diseases of aortic valve
C1260908|ICD9CM|HT|956|Injury to peripheral nerve(s) of pelvic girdle and lower limb
C1260915|ICD9CM|PT|096|Late syphilis, latent
C1260915|ICD9CM|AB|096|Late syphilis latent
C1260922|ICD9CM|PT|786.00|Respiratory abnormality, unspecified
C1260922|ICD9CM|AB|786.00|Respiratory abnorm NOS
C1261016|ICD9CM|AB|65.92|Transplantation of ovary
C1261016|ICD9CM|PT|65.92|Transplantation of ovary
C1261176|ICD9CM|PT|751.1|Atresia and stenosis of small intestine
C1261176|ICD9CM|AB|751.1|Atresia small intestine
C1261251|ICD9CM|PT|752.45|Vaginal agenesis
C1261251|ICD9CM|AB|752.45|Vaginal agenesis
C1261262|ICD9CM|HT|642.9|Unspecified hypertension complicating pregnancy, childbirth, or the puerperium
C1261276|ICD9CM|PT|754.32|Congenital subluxation of hip, unilateral
C1261276|ICD9CM|AB|754.32|Cong hip sublux, unilat
C1261278|ICD9CM|AB|595.3|Trigonitis
C1261278|ICD9CM|PT|595.3|Trigonitis
C1261281|ICD9CM|PT|996.81|Complications of transplanted kidney
C1261281|ICD9CM|AB|996.81|Compl kidney transplant
C1261282|ICD9CM|PT|996.82|Complications of transplanted liver
C1261282|ICD9CM|AB|996.82|Compl liver transplant
C1261289|ICD9CM|PT|77.45|Biopsy of bone, femur
C1261289|ICD9CM|AB|77.45|Femoral biopsy
C1261292|ICD9CM|PT|35.42|Creation of septal defect in heart
C1261292|ICD9CM|AB|35.42|Create septal defect
C1261295|ICD9CM|PT|52.11|Closed [aspiration] [needle] [percutaneous] biopsy of pancreas
C1261295|ICD9CM|AB|52.11|Closed pancreatic biopsy
C1261297|ICD9CM|PT|58.92|Excision of periurethral tissue
C1261297|ICD9CM|AB|58.92|Periurethral excision
C1261298|ICD9CM|AB|64.44|Reconstruction of penis
C1261298|ICD9CM|PT|64.44|Reconstruction of penis
C1261299|ICD9CM|PT|70.77|Vaginal suspension and fixation
C1261299|ICD9CM|AB|70.77|Vaginal suspens & fixat
C1261300|ICD9CM|PT|70.51|Repair of cystocele
C1261300|ICD9CM|AB|70.51|Cystocele repair
C1261304|ICD9CM|PT|10.0|Removal of embedded foreign body from conjunctiva by incision
C1261304|ICD9CM|AB|10.0|Incise/remov conjunct FB
C1261307|ICD9CM|PT|15.21|Lengthening procedure on one extraocular muscle
C1261307|ICD9CM|AB|15.21|Lengthen 1 extraoc musc
C1261308|ICD9CM|PT|15.22|Shortening procedure on one extraocular muscle
C1261308|ICD9CM|AB|15.22|Shorten 1 extraoc musc
C1261309|ICD9CM|PT|34.23|Biopsy of chest wall
C1261309|ICD9CM|AB|34.23|Chest wall biopsy
C1261311|ICD9CM|PT|99.23|Injection of steroid
C1261311|ICD9CM|AB|99.23|Inject steroid
C1261312|ICD9CM|PT|99.35|Vaccination against tularemia
C1261312|ICD9CM|AB|99.35|Tularemia vaccination
C1261318|ICD9CM|PT|115.05|Infection by Histoplasma capsulatum, pneumonia
C1261318|ICD9CM|AB|115.05|Histoplasm caps pneumon
C1261319|ICD9CM|PT|635.92|Legally induced abortion, without mention of complication, complete
C1261319|ICD9CM|AB|635.92|Legal abort uncompl-comp
C1261324|ICD9CM|PT|V67.2|Follow-up examination, following chemotherapy
C1261324|ICD9CM|AB|V67.2|Chemotherapy follow-up
C1261325|ICD9CM|PT|V16.3|Family history of malignant neoplasm of breast
C1261325|ICD9CM|AB|V16.3|Family hx-breast malig
C1261328|ICD9CM|HT|V18.6|Family history of kidney diseases
C1261331|ICD9CM|AB|362.54|Macular cyst or hole
C1261331|ICD9CM|PT|362.54|Macular cyst, hole, or pseudohole
C1261332|ICD9CM|PT|03.02|Reopening of laminectomy site
C1261332|ICD9CM|AB|03.02|Reopen laminectomy site
C1261378|ICD9CM|HT|V16|Family history of malignant neoplasm
C1261378|ICD9CM|PT|V16.9|Family history of unspecified malignant neoplasm
C1261378|ICD9CM|AB|V16.9|Family hx-malignancy NOS
C1261514|ICD9CM|AB|86.65|Heterograft to skin
C1261514|ICD9CM|PT|86.65|Heterograft to skin
C1261518|ICD9CM|AB|46.97|Transplant of intestine
C1261518|ICD9CM|PT|46.97|Transplant of intestine
C1262477|ICD9CM|AB|783.21|Abnormal loss of weight
C1262477|ICD9CM|PT|783.21|Loss of weight
C1262481|ICD9CM|PT|558.41|Eosinophilic gastroenteritis
C1262481|ICD9CM|AB|558.41|Eosinophilic gastroent
C1263817|ICD9CM|HT|637.2|Unspecified abortion complicated by damage to pelvic organs or tissues
C1263817|ICD9CM|PT|637.20|Unspecified abortion, complicated by damage to pelvic organs or tissues, unspecified
C1263817|ICD9CM|AB|637.20|Ab NOS w pelv damag-unsp
C1263846|ICD9CM|PT|314.01|Attention deficit disorder with hyperactivity
C1263846|ICD9CM|HT|314|Hyperkinetic syndrome of childhood
C1263846|ICD9CM|PT|314.9|Unspecified hyperkinetic syndrome
C1263846|ICD9CM|AB|314.9|Hyperkinetic synd NOS
C1263846|ICD9CM|AB|314.01|Attn deficit w hyperact
C1263961|ICD9CM|PT|251.9|Unspecified disorder of pancreatic internal secretion
C1263961|ICD9CM|AB|251.9|Pancreatic disorder NOS
C1264275|ICD9CM|PT|834.02|Closed dislocation of interphalangeal (joint), hand
C1264275|ICD9CM|AB|834.02|Disl interphaln hand-cl
C1264623|ICD9CM|PT|053.10|Herpes zoster with unspecified nervous system complication
C1264623|ICD9CM|AB|053.10|H zoster nerv syst NOS
C1266194|ICD9CM|HT|201.4|Hodgkin's disease, lymphocytic-histiocytic predominance
C1269750|ICD9CM|PT|290.20|Senile dementia with delusional features
C1269750|ICD9CM|AB|290.20|Senile delusion
C1270937|ICD9CM|AB|96.14|Vaginal packing
C1270937|ICD9CM|PT|96.14|Vaginal packing
C1271437|ICD9CM|AB|70.21|Vaginoscopy
C1271437|ICD9CM|PT|70.21|Vaginoscopy
C1272092|ICD9CM|AB|790.21|Impaired fasting glucose
C1272092|ICD9CM|PT|790.21|Impaired fasting glucose
C1274184|ICD9CM|AB|698.4|Dermatitis factitia
C1274184|ICD9CM|PT|698.4|Dermatitis factitia [artefacta]
C1274259|ICD9CM|PT|173.01|Basal cell carcinoma of skin of lip
C1274259|ICD9CM|AB|173.01|Basal cell ca skin lip
C1274329|ICD9CM|PT|058.12|Roseola infantum due to human herpesvirus 7
C1274329|ICD9CM|AB|058.12|Roseola infant d/t HHV-7
C1275737|ICD9CM|AB|19.52|Type 2 tympanoplasty
C1275737|ICD9CM|PT|19.52|Type II tympanoplasty
C1275806|ICD9CM|HT|664.3|Fourth-degree perineal laceration during delivery
C1275806|ICD9CM|PT|664.31|Fourth-degree perineal laceration, delivered, with or without mention of antepartum condition
C1275806|ICD9CM|AB|664.31|Del w 4 deg lacerat-del
C1278558|ICD9CM|PT|E918|Caught accidentally in or between objects
C1278558|ICD9CM|AB|E918|Caught between objects
C1278561|ICD9CM|AB|E978|Legal execution
C1278561|ICD9CM|PT|E978|Legal execution
C1278681|ICD9CM|PT|48.82|Excision of perirectal tissue
C1278681|ICD9CM|AB|48.82|Perirectal excision
C1278807|ICD9CM|PT|099.41|Other nongonococcal urethritis, chlamydia trachomatis
C1278807|ICD9CM|AB|099.41|Chlmyd trachomatis ureth
C1279224|ICD9CM|PT|009.0|Infectious colitis, enteritis, and gastroenteritis
C1279224|ICD9CM|AB|009.0|Infectious enteritis NOS
C1279258|ICD9CM|PT|182.0|Malignant neoplasm of corpus uteri, except isthmus
C1279258|ICD9CM|AB|182.0|Malig neo corpus uteri
C1279296|ICD9CM|HT|208.1|Leukemia of unspecified cell type, chronic
C1279396|ICD9CM|HT|533.7|Chronic peptic ulcer of unspecified site without mention of hemorrhage or perforation
C1279412|ICD9CM|PT|359.3|Periodic paralysis
C1279412|ICD9CM|AB|359.3|Periodic paralysis
C1279573|ICD9CM|PT|890.0|Open wound of hip and thigh, without mention of complication
C1279573|ICD9CM|AB|890.0|Open wound of hip/thigh
C1279739|ICD9CM|AB|83.81|Tendon graft
C1279739|ICD9CM|PT|83.81|Tendon graft
C1279945|ICD9CM|PT|516.33|Acute interstitial pneumonitis
C1279945|ICD9CM|AB|516.33|Acute interstitial pneum
C1280859|ICD9CM|PT|77.46|Biopsy of bone, patella
C1280859|ICD9CM|AB|77.46|Patellar biopsy
C1281543|ICD9CM|AB|94.23|Neuroleptic therapy
C1281543|ICD9CM|PT|94.23|Neuroleptic therapy
C1281603|ICD9CM|AB|94.21|Narcoanalysis
C1281603|ICD9CM|PT|94.21|Narcoanalysis
C1281729|ICD9CM|PT|836.0|Tear of medial cartilage or meniscus of knee, current
C1281729|ICD9CM|AB|836.0|Tear med menisc knee-cur
C1281794|ICD9CM|PT|836.1|Tear of lateral cartilage or meniscus of knee, current
C1281794|ICD9CM|AB|836.1|Tear lat menisc knee-cur
C1282883|ICD9CM|PT|52.81|Reimplantation of pancreatic tissue
C1282883|ICD9CM|AB|52.81|Reimplant pancreatic tis
C1282912|ICD9CM|PT|732.4|Juvenile osteochondrosis of lower extremity, excluding foot
C1282912|ICD9CM|AB|732.4|Juv osteochondrosis leg
C1282937|ICD9CM|PT|46.71|Suture of laceration of duodenum
C1282937|ICD9CM|AB|46.71|Duodenal lacerat suture
C1282983|ICD9CM|PT|082.41|Ehrlichiosis chafeensis [E. chafeensis]
C1282983|ICD9CM|AB|082.41|Ehrlichiosis chafeensis
C1283021|ICD9CM|PT|80.78|Synovectomy, foot and toe
C1283021|ICD9CM|AB|80.78|Foot synovectomy
C1285368|ICD9CM|HT|776|Hematological disorders of newborn
C1288279|ICD9CM|PT|354.2|Lesion of ulnar nerve
C1288279|ICD9CM|AB|354.2|Ulnar nerve lesion
C1290220|ICD9CM|PT|738.10|Unspecified acquired deformity of head
C1290220|ICD9CM|AB|738.10|Unspf acq deformity head
C1290744|ICD9CM|AB|525.61|Open restoration margins
C1290744|ICD9CM|PT|525.61|Open restoration margins
C1290810|ICD9CM|PT|070.1|Viral hepatitis A without mention of hepatic coma
C1290810|ICD9CM|AB|070.1|Hepatitis A w/o coma
C1291056|ICD9CM|PT|524.54|Insufficient anterior guidance
C1291056|ICD9CM|AB|524.54|Insuff anterior guidance
C1292772|ICD9CM|HT|205.2|Myeloid leukemia, subacute
C1292779|ICD9CM|PT|238.74|Myelodysplastic syndrome with 5q deletion
C1292779|ICD9CM|AB|238.74|Myelodyspls syn w 5q del
C1292969|ICD9CM|HT|00.6|Procedures on blood vessels
C1293003|ICD9CM|PT|71.9|Other operations on female genital organs
C1293003|ICD9CM|AB|71.9|Other female genital ops
C1293256|ICD9CM|AB|84.04|Disarticulation of wrist
C1293256|ICD9CM|PT|84.04|Disarticulation of wrist
C1293595|ICD9CM|PT|41.33|Open biopsy of spleen
C1293595|ICD9CM|AB|41.33|Open spleen biopsy
C1293675|ICD9CM|PT|68.14|Open biopsy of uterine ligaments
C1293675|ICD9CM|AB|68.14|Open uterine ligament bx
C1297885|ICD9CM|HT|79.3|Open reduction of fracture with internal fixation
C1298685|ICD9CM|PT|338.4|Chronic pain syndrome
C1298685|ICD9CM|AB|338.4|Chronic pain syndrome
C1298714|ICD9CM|PT|753.21|Congenital obstruction of ureteropelvic junction
C1298714|ICD9CM|AB|753.21|Congen obst urtroplv jnc
C1299558|ICD9CM|HT|637.8|Unspecified abortion with unspecified complication
C1299558|ICD9CM|PT|637.80|Unspecified abortion, with unspecified complication, unspecified
C1299558|ICD9CM|AB|637.80|Ab NOS w compl NOS-unsp
C1299919|ICD9CM|AB|007.2|Coccidiosis
C1299919|ICD9CM|PT|007.2|Coccidiosis
C1300133|ICD9CM|PT|375.03|Chronic enlargement of lacrimal gland
C1300133|ICD9CM|AB|375.03|Ch enlargmnt lacrim glnd
C1300597|ICD9CM|PT|02.01|Opening of cranial suture
C1300597|ICD9CM|AB|02.01|Linear craniectomy
C1301937|ICD9CM|AB|754.70|Talipes NOS
C1301937|ICD9CM|PT|754.70|Talipes, unspecified
C1302169|ICD9CM|PT|99.39|Administration of diphtheria-tetanus-pertussis, combined
C1302169|ICD9CM|AB|99.39|Dpt administration
C1302325|ICD9CM|PT|355.4|Lesion of medial popliteal nerve
C1302325|ICD9CM|AB|355.4|Med popliteal nerve les
C1302752|ICD9CM|AB|521.20|Abrasion NOS
C1302752|ICD9CM|PT|521.20|Abrasion, unspecified
C1304542|ICD9CM|PT|83.84|Release of clubfoot, not elsewhere classified
C1304542|ICD9CM|AB|83.84|Clubfoot release NEC
C1304652|ICD9CM|HT|82.7|Plastic operation on hand with graft or implant
C1304679|ICD9CM|PT|35.61|Repair of atrial septal defect with tissue graft
C1304679|ICD9CM|AB|35.61|Graft repair atrial def
C1304875|ICD9CM|PT|67.32|Destruction of lesion of cervix by cauterization
C1304875|ICD9CM|AB|67.32|Cervical les cauterizat
C1304878|ICD9CM|PT|80.26|Arthroscopy, knee
C1304878|ICD9CM|AB|80.26|Knee arthroscopy
C1305122|ICD9CM|PT|441.6|Thoracoabdominal aneurysm, ruptured
C1305122|ICD9CM|AB|441.6|Thoracoabd aneurysm rupt
C1305875|ICD9CM|AB|610.2|Fibroadenosis of breast
C1305875|ICD9CM|PT|610.2|Fibroadenosis of breast
C1305927|ICD9CM|HT|758.8|Other conditions due to chromosome anomalies
C1305927|ICD9CM|PT|758.89|Other conditions due to chromosome anomalies
C1305927|ICD9CM|AB|758.89|Oth con d/t chrm anm NEC
C1305934|ICD9CM|HT|610|Benign mammary dysplasias
C1305934|ICD9CM|AB|610.9|Benign mamm dysplas NOS
C1305934|ICD9CM|PT|610.9|Benign mammary dysplasia, unspecified
C1305964|ICD9CM|PT|753.6|Atresia and stenosis of urethra and bladder neck
C1305964|ICD9CM|AB|753.6|Congen urethral stenosis
C1306015|ICD9CM|PT|940.0|Chemical burn of eyelids and periocular area
C1306015|ICD9CM|AB|940.0|Chemical burn periocular
C1306068|ICD9CM|HT|366.5|After-cataract
C1306068|ICD9CM|AB|366.50|After-cataract NOS
C1306068|ICD9CM|PT|366.50|After-cataract, unspecified
C1306110|ICD9CM|PT|840.3|Infraspinatus (muscle) (tendon) sprain
C1306110|ICD9CM|AB|840.3|Sprain infraspinatus
C1306122|ICD9CM|PT|368.61|Congenital night blindness
C1306122|ICD9CM|AB|368.61|Congen night blindness
C1306154|ICD9CM|PT|811.13|Open fracture of glenoid cavity and neck of scapula
C1306154|ICD9CM|AB|811.13|Fx scap, glen cav/nck-op
C1306246|ICD9CM|PT|345.40|Localization-related (focal) (partial) epilepsy and epileptic syndromes with complex partial seizures, without mention of intractable epilepsy
C1306246|ICD9CM|AB|345.40|Psymotr epil w/o int epi
C1306306|ICD9CM|PT|718.45|Contracture of joint, pelvic region and thigh
C1306306|ICD9CM|AB|718.45|Jt contracture-pelvis
C1306315|ICD9CM|PT|83.75|Tendon transfer or transplantation
C1306315|ICD9CM|AB|83.75|Tendon trnsfr/transplant
C1306506|ICD9CM|PT|04.02|Division of trigeminal nerve
C1306506|ICD9CM|AB|04.02|Trigeminal nerv division
C1306539|ICD9CM|PT|31.71|Suture of laceration of trachea
C1306539|ICD9CM|AB|31.71|Suture of tracheal lacer
C1306540|ICD9CM|PT|33.41|Suture of laceration of bronchus
C1306540|ICD9CM|AB|33.41|Bronchial lacerat suture
C1306585|ICD9CM|HT|79.2|Open reduction of fracture without internal fixation
C1306605|ICD9CM|HT|156|Malignant neoplasm of gallbladder and extrahepatic bile ducts
C1306638|ICD9CM|PT|201.93|Hodgkin's disease, unspecified type, intra-abdominal lymph nodes
C1306638|ICD9CM|AB|201.93|Hodgkins dis NOS abdom
C1306794|ICD9CM|PT|040.42|Wound botulism
C1306794|ICD9CM|AB|040.42|Wound botulism
C1306822|ICD9CM|PT|396.2|Mitral valve insufficiency and aortic valve stenosis
C1306822|ICD9CM|AB|396.2|Mitral insuf/aort stenos
C1306848|ICD9CM|AB|072.9|Mumps uncomplicated
C1306848|ICD9CM|PT|072.9|Mumps without mention of complication
C1306873|ICD9CM|HT|993|Effects of air pressure
C1306891|ICD9CM|PT|V69.0|Lack of physical exercise
C1306891|ICD9CM|AB|V69.0|Lack of physical exercse
C1313860|ICD9CM|PT|V61.6|Illegitimacy or illegitimate pregnancy
C1313860|ICD9CM|AB|V61.6|Illegitimate pregnancy
C1313863|ICD9CM|AB|908.9|Late effect injury NOS
C1313863|ICD9CM|PT|908.9|Late effect of unspecified injury
C1313876|ICD9CM|HT|764.0|"Light-for-dates" without mention of fetal malnutrition
C1313885|ICD9CM|AB|757.0|Hereditary edema of legs
C1313885|ICD9CM|PT|757.0|Hereditary edema of legs
C1313895|ICD9CM|HT|V30|Single liveborn
C1313895|ICD9CM|PT|V27.0|Outcome of delivery, single liveborn
C1313895|ICD9CM|AB|V27.0|Deliver-single liveborn
C1313896|ICD9CM|PT|V27.1|Outcome of delivery, single stillborn
C1313896|ICD9CM|AB|V27.1|Deliver-single stillborn
C1313924|ICD9CM|PT|V73.4|Screening examination for yellow fever
C1313924|ICD9CM|AB|V73.4|Screening-yellow fever
C1313933|ICD9CM|AB|V59.2|Bone donor
C1313933|ICD9CM|PT|V59.2|Bone donors
C1313934|ICD9CM|AB|V59.3|Bone marrow donor
C1313934|ICD9CM|PT|V59.3|Bone marrow donors
C1313935|ICD9CM|AB|V59.4|Kidney donor
C1313935|ICD9CM|PT|V59.4|Kidney donors
C1313951|ICD9CM|HT|V59.0|Blood donors
C1314803|ICD9CM|HT|360-379.99|DISORDERS OF THE EYE AND ADNEXA
C1314803|ICD9CM|HT|379.9|Unspecified disorder of eye and adnexa
C1314968|ICD9CM|AB|694.3|Impetigo herpetiformis
C1314968|ICD9CM|PT|694.3|Impetigo herpetiformis
C1318464|ICD9CM|AB|93.83|Occupational therapy
C1318464|ICD9CM|PT|93.83|Occupational therapy
C1318500|ICD9CM|PT|241.9|Unspecified nontoxic nodular goiter
C1318500|ICD9CM|HT|241|Nontoxic nodular goiter
C1318500|ICD9CM|AB|241.9|Nontox nodul goiter NOS
C1318512|ICD9CM|PT|862.22|Injury to esophagus without mention of open wound into cavity
C1318512|ICD9CM|AB|862.22|Esophagus injury-closed
C1318514|ICD9CM|PT|674.14|Disruption of cesarean wound, postpartum condition or complication
C1318514|ICD9CM|AB|674.14|Disrupt c-sect-postpart
C1318533|ICD9CM|AB|289.0|Secondary polycythemia
C1318533|ICD9CM|PT|289.0|Polycythemia, secondary
C1318543|ICD9CM|PT|727.02|Giant cell tumor of tendon sheath
C1318543|ICD9CM|AB|727.02|Giant cell tumor tendon
C1318552|ICD9CM|PT|432.0|Nontraumatic extradural hemorrhage
C1318552|ICD9CM|AB|432.0|Nontraum extradural hem
C1318565|ICD9CM|AB|006.6|Amebic skin ulceration
C1318565|ICD9CM|PT|006.6|Amebic skin ulceration
C1320634|ICD9CM|PT|98.27|Removal of foreign body without incision from upper limb, except hand
C1320634|ICD9CM|AB|98.27|Removal FB from arm
C1320640|ICD9CM|HT|362.6|Peripheral retinal degenerations
C1320640|ICD9CM|PT|362.60|Peripheral retinal degeneration, unspecified
C1320640|ICD9CM|AB|362.60|Periph retina degen NOS
C1321345|ICD9CM|PT|364.82|Plateau iris syndrome
C1321345|ICD9CM|AB|364.82|Plateau iris syndrome
C1321831|ICD9CM|HT|V46.1|Dependence on respirator [Ventilator]
C1321896|ICD9CM|AB|956.3|Injury peroneal nerve
C1321896|ICD9CM|PT|956.3|Injury to peroneal nerve
C1321898|ICD9CM|AB|578.1|Blood in stool
C1321898|ICD9CM|PT|578.1|Blood in stool
C1321926|ICD9CM|PT|951.0|Injury to oculomotor nerve
C1321926|ICD9CM|AB|951.0|Injury oculomotor nerve
C1328252|ICD9CM|PT|085.5|Mucocutaneous leishmaniasis, (American)
C1328252|ICD9CM|AB|085.5|Mucocutan leishmaniasis
C1328333|ICD9CM|PT|372.34|Pingueculitis
C1328333|ICD9CM|AB|372.34|Pingueculitis
C1328479|ICD9CM|PT|157.4|Malignant neoplasm of islets of langerhans
C1328479|ICD9CM|AB|157.4|Mal neo islet langerhans
C1328840|ICD9CM|PT|279.41|Autoimmune lymphoproliferative syndrome
C1328840|ICD9CM|AB|279.41|Autoimmun lymphprof synd
C1328971|ICD9CM|PT|722.2|Displacement of intervertebral disc, site unspecified, without myelopathy
C1328971|ICD9CM|AB|722.2|Disc displacement NOS
C1331611|ICD9CM|PT|905.1|Late effect of fracture of spine and trunk without mention of spinal cord lesion
C1331611|ICD9CM|AB|905.1|Late eff spine/trunk fx
C1333139|ICD9CM|PT|621.32|Complex endometrial hyperplasia without atypia
C1333139|ICD9CM|AB|621.32|Comp endo hyper w/o atyp
C1335929|ICD9CM|PT|237.73|Schwannomatosis
C1335929|ICD9CM|AB|237.73|Schwannomatosis
C1335967|ICD9CM|PT|621.31|Simple endometrial hyperplasia without atypia
C1335967|ICD9CM|AB|621.31|Simp endo hyper w/o atyp
C1336746|ICD9CM|PT|209.22|Malignant carcinoid tumor of the thymus
C1336746|ICD9CM|AB|209.22|Malig carcinoid thymus
C1363843|ICD9CM|PT|362.13|Changes in vascular appearance of retina
C1363843|ICD9CM|AB|362.13|Retinal vascular changes
C1363999|ICD9CM|PT|006.0|Acute amebic dysentery without mention of abscess
C1363999|ICD9CM|AB|006.0|Ac amebiasis w/o abscess
C1366330|ICD9CM|PT|896.0|Traumatic amputation of foot (complete) (partial), unilateral, without mention of complication
C1366330|ICD9CM|AB|896.0|Amputation foot, unilat
C1367654|ICD9CM|HT|200.3|Marginal zone lymphoma
C1367972|ICD9CM|HT|451|Phlebitis and thrombophlebitis
C1367972|ICD9CM|PT|451.9|Phlebitis and thrombophlebitis of unspecified site
C1367972|ICD9CM|AB|451.9|Thrombophlebitis NOS
C1367974|ICD9CM|PT|694.60|Benign mucous membrane pemphigoid without mention of ocular involvement
C1367974|ICD9CM|AB|694.60|Bn mucous memb pemph NOS
C1370824|ICD9CM|AB|518.1|Interstitial emphysema
C1370824|ICD9CM|PT|518.1|Interstitial emphysema
C1370867|ICD9CM|PT|986|Toxic effect of carbon monoxide
C1370867|ICD9CM|AB|986|Tox eff carbon monoxide
C1377996|ICD9CM|AB|70.61|Vaginal construction
C1377996|ICD9CM|PT|70.61|Vaginal construction
C1384485|ICD9CM|AB|650|Normal delivery
C1384485|ICD9CM|PT|650|Normal delivery
C1384500|ICD9CM|PT|E858.7|Accidental poisoning by agents primarily affecting skin and mucous membrane, ophthalmological, otorhinolaryngological, and dental drugs
C1384500|ICD9CM|AB|E858.7|Acc poisn-skin/eent agnt
C1384514|ICD9CM|AB|255.12|Conn's syndrome
C1384514|ICD9CM|PT|255.12|Conn's syndrome
C1384584|ICD9CM|HT|715.0|Osteoarthrosis, generalized
C1384584|ICD9CM|PT|715.09|Osteoarthrosis, generalized, multiple sites
C1384584|ICD9CM|AB|715.09|General osteoarthrosis
C1384587|ICD9CM|PT|543.0|Hyperplasia of appendix (lymphoid)
C1384587|ICD9CM|AB|543.0|Hyperplasia of appendix
C1384591|ICD9CM|HT|73.0|Artificial rupture of membranes
C1384593|ICD9CM|PT|89.34|Digital examination of rectum
C1384593|ICD9CM|AB|89.34|Digital rectal exam
C1384594|ICD9CM|AB|593.0|Nephroptosis
C1384594|ICD9CM|PT|593.0|Nephroptosis
C1384596|ICD9CM|AB|22.2|Intranasal antrotomy
C1384596|ICD9CM|PT|22.2|Intranasal antrotomy
C1384631|ICD9CM|HT|534|Gastrojejunal ulcer
C1384666|ICD9CM|HT|389|Hearing loss
C1384666|ICD9CM|AB|389.9|Hearing loss NOS
C1384666|ICD9CM|PT|389.9|Unspecified hearing loss
C1384683|ICD9CM|PT|V42.5|Cornea replaced by transplant
C1384683|ICD9CM|AB|V42.5|Cornea transplant status
C1384687|ICD9CM|PT|126.0|Ancylostomiasis due to ancylostoma duodenale
C1384687|ICD9CM|AB|126.0|Ancylostoma duodenale
C1386808|ICD9CM|HT|V88.1|Acquired absence of pancreas
C1390180|ICD9CM|PT|772.6|Cutaneous hemorrhage of fetus or newborn
C1390180|ICD9CM|AB|772.6|NB cutaneous hemorrhage
C1395264|ICD9CM|PT|110.6|Deep seated dermatophytosis
C1395264|ICD9CM|AB|110.6|Deep dermatophytosis
C1399001|ICD9CM|PT|V21.0|Period of rapid growth in childhood
C1399001|ICD9CM|AB|V21.0|Rapid childhood growth
C1399262|ICD9CM|PT|V75.7|Screening examination for intestinal helminthiasis
C1399262|ICD9CM|AB|V75.7|Screen for helminthiasis
C1401143|ICD9CM|AB|V45.3|Intestinal bypass status
C1401143|ICD9CM|PT|V45.3|Intestinal bypass or anastomosis status
C1403891|ICD9CM|PT|036.3|Waterhouse-Friderichsen syndrome, meningococcal
C1403891|ICD9CM|AB|036.3|Meningococc adrenal synd
C1404542|ICD9CM|AB|359.24|Drug induced myotonia
C1404542|ICD9CM|PT|359.24|Drug- induced myotonia
C1410098|ICD9CM|PT|779.85|Cardiac arrest of newborn
C1410098|ICD9CM|AB|779.85|NB cardiac arrest
C1439344|ICD9CM|PT|996.90|Complications of unspecified reattached extremity
C1439344|ICD9CM|AB|996.90|Comp reattach extrem NOS
C1442831|ICD9CM|HT|716|Other and unspecified arthropathies
C1442831|ICD9CM|HT|719|Other and unspecified disorders of joint
C1442839|ICD9CM|PT|278.4|Hypervitaminosis D
C1442839|ICD9CM|AB|278.4|Hypervitaminosis d
C1442861|ICD9CM|AB|921.0|Black eye NOS
C1442861|ICD9CM|PT|921.0|Black eye, not otherwise specified
C1442902|ICD9CM|HT|726|Peripheral enthesopathies and allied syndromes
C1442903|ICD9CM|PT|726.91|Exostosis of unspecified site
C1442903|ICD9CM|AB|726.91|Exostosis, site NOS
C1442952|ICD9CM|PT|723.4|Brachial neuritis or radiculitis NOS
C1442952|ICD9CM|AB|723.4|Brachial neuritis NOS
C1442967|ICD9CM|PT|533.10|Acute peptic ulcer of unspecified site with perforation, without mention of obstruction
C1442967|ICD9CM|AB|533.10|Ac peptic ulcer w perfor
C1442980|ICD9CM|PT|552.21|Incisional ventral hernia with obstruction
C1442980|ICD9CM|AB|552.21|Obstr incisional hernia
C1442981|ICD9CM|AB|571.3|Alcohol liver damage NOS
C1442981|ICD9CM|PT|571.3|Alcoholic liver damage, unspecified
C1443010|ICD9CM|PT|944.37|Full-thickness skin loss [third degree, not otherwise specified] of wrist
C1443010|ICD9CM|AB|944.37|3rd deg burn wrist
C1443011|ICD9CM|PT|944.27|Blisters, epidermal loss [second degree] of wrist
C1443011|ICD9CM|AB|944.27|2nd deg burn wrist
C1443030|ICD9CM|HT|965.0|Poisoning by opiates and related narcotics
C1443291|ICD9CM|PT|354.4|Causalgia of upper limb
C1443291|ICD9CM|AB|354.4|Causalgia upper limb
C1443352|ICD9CM|PT|73.01|Induction of labor by artificial rupture of membranes
C1443352|ICD9CM|AB|73.01|Induct labor-rupt memb
C1443381|ICD9CM|AB|362.23|Retinoph prematr,stage 1
C1443381|ICD9CM|PT|362.23|Retinopathy of prematurity, stage 1
C1443382|ICD9CM|PT|362.24|Retinopathy of prematurity, stage 2
C1443382|ICD9CM|AB|362.24|Retinoph prematr,stage 2
C1443383|ICD9CM|AB|362.25|Retinoph prematr,stage 3
C1443383|ICD9CM|PT|362.25|Retinopathy of prematurity, stage 3
C1443384|ICD9CM|PT|362.26|Retinopathy of prematurity, stage 4
C1443384|ICD9CM|AB|362.26|Retinoph prematr.stage 4
C1443385|ICD9CM|AB|362.27|Retinoph prematr,stage 5
C1443385|ICD9CM|PT|362.27|Retinopathy of prematurity, stage 5
C1443972|ICD9CM|AB|600.3|Cyst of prostate
C1443972|ICD9CM|PT|600.3|Cyst of prostate
C1443978|ICD9CM|PT|733.14|Pathologic fracture of neck of femur
C1443978|ICD9CM|AB|733.14|Path fx neck of femur
C1444204|ICD9CM|PT|831.12|Open posterior dislocation of humerus
C1444204|ICD9CM|AB|831.12|Post disloc humerus-open
C1444208|ICD9CM|HT|330-337.99|HEREDITARY AND DEGENERATIVE DISEASES OF THE CENTRAL NERVOUS SYSTEM
C1449721|ICD9CM|PT|778.7|Breast engorgement in newborn
C1449721|ICD9CM|AB|778.7|NB breast engorgement
C1455742|ICD9CM|HT|381.2|Chronic mucoid otitis media
C1455742|ICD9CM|PT|381.20|Chronic mucoid otitis media, simple or unspecified
C1455742|ICD9CM|AB|381.20|Chr mucoid OM simp/NOS
C1455852|ICD9CM|PT|89.49|Automatic implantable cardioverter/defibrillator (AICD) check
C1455852|ICD9CM|AB|89.49|AICD check
C1455856|ICD9CM|HT|89.4|Cardiac stress tests and pacemaker and defibrillator checks
C1455876|ICD9CM|PT|79.02|Closed reduction of fracture without internal fixation, radius and ulna
C1455876|ICD9CM|AB|79.02|Cl fx reduc-radius/ulna
C1455877|ICD9CM|PT|79.03|Closed reduction of fracture without internal fixation, carpals and metacarpals
C1455877|ICD9CM|AB|79.03|Cl fx reduc-metacar/car
C1455878|ICD9CM|PT|79.04|Closed reduction of fracture without internal fixation, phalanges of hand
C1455878|ICD9CM|AB|79.04|Cl fx reduc-finger
C1455879|ICD9CM|PT|79.05|Closed reduction of fracture without internal fixation, femur
C1455879|ICD9CM|AB|79.05|Cl fx reduc-femur
C1455880|ICD9CM|PT|79.06|Closed reduction of fracture without internal fixation, tibia and fibula
C1455880|ICD9CM|AB|79.06|Cl fx reduc-tibia/fibula
C1455881|ICD9CM|PT|79.07|Closed reduction of fracture without internal fixation, tarsals and metatarsals
C1455881|ICD9CM|AB|79.07|Cl fx reduc-metatar/tar
C1455882|ICD9CM|PT|79.08|Closed reduction of fracture without internal fixation, phalanges of foot
C1455882|ICD9CM|AB|79.08|Cl fx reduc-toe
C1455883|ICD9CM|PT|79.09|Closed reduction of fracture without internal fixation, other specified bone
C1455883|ICD9CM|AB|79.09|Closed fx reduction NEC
C1455884|ICD9CM|PT|790.95|Elevated C-reactive protein (CRP)
C1455884|ICD9CM|AB|790.95|Elev C-reactive protein
C1455885|ICD9CM|PT|795.00|Abnormal glandular Papanicolaou smear of cervix
C1455885|ICD9CM|AB|795.00|Abn glandular pap smear
C1455889|ICD9CM|PT|795.01|Papanicolaou smear of cervix with atypical squamous cells of undetermined significance (ASC-US)
C1455889|ICD9CM|AB|795.01|Pap smear (ASC-US)
C1455890|ICD9CM|PT|795.02|Papanicolaou smear of cervix with atypical squamous cells cannot exclude high grade squamous intraepithelial lesion (ASC-H)
C1455890|ICD9CM|AB|795.02|Pap smear (ASC-H)
C1455891|ICD9CM|PT|795.03|Papanicolaou smear of cervix with low grade squamous intraepithelial lesion (LGSIL)
C1455891|ICD9CM|AB|795.03|Pap smear cervix w LGSIL
C1455892|ICD9CM|PT|795.04|Papanicolaou smear of cervix with high grade squamous intraepithelial lesion (HGSIL)
C1455892|ICD9CM|AB|795.04|Pap smear cervix w HGSIL
C1455894|ICD9CM|PT|795.05|Cervical high risk human papillomavirus (HPV) DNA test positive
C1455894|ICD9CM|AB|795.05|Cervical (HPV) DNA pos
C1455897|ICD9CM|PT|795.09|Other abnormal Papanicolaou smear of cervix and cervical HPV
C1455897|ICD9CM|AB|795.09|Abn pap cervix HPV NEC
C1455899|ICD9CM|HT|795.0|Abnormal Papanicolaou smear of cervix and cervical HPV
C1455902|ICD9CM|HT|795|Other and nonspecific abnormal cytological, histological, immunological and DNA test findings
C1455903|ICD9CM|AB|796.6|Abnorm neonate screening
C1455903|ICD9CM|PT|796.6|Abnormal findings on neonatal screening
C1455904|ICD9CM|AB|99.78|Aquapheresis
C1455904|ICD9CM|PT|99.78|Aquapheresis
C1455908|ICD9CM|PT|84.53|Implantation of internal limb lengthening device with kinetic distraction
C1455908|ICD9CM|AB|84.53|Imp limb length kinetic
C1455909|ICD9CM|PT|84.54|Implantation of other internal limb lengthening device
C1455909|ICD9CM|AB|84.54|Impl other limb length
C1455910|ICD9CM|PT|84.55|Insertion of bone void filler
C1455910|ICD9CM|AB|84.55|Ins bone void filler
C1455915|ICD9CM|PT|84.59|Insertion of other spinal devices
C1455915|ICD9CM|AB|84.59|Insert othr spin device
C1455916|ICD9CM|PT|84.60|Insertion of spinal disc prosthesis, not otherwise specified
C1455916|ICD9CM|AB|84.60|Insert disc pros NOS
C1455918|ICD9CM|PT|84.61|Insertion of partial spinal disc prosthesis, cervical
C1455918|ICD9CM|AB|84.61|Ins part disc pros cerv
C1455922|ICD9CM|PT|84.62|Insertion of total spinal disc prosthesis, cervical
C1455922|ICD9CM|AB|84.62|Ins tot disc prost cerv
C1455926|ICD9CM|PT|84.63|Insertion of spinal disc prosthesis, thoracic
C1455926|ICD9CM|AB|84.63|Ins spin disc pros thor
C1455930|ICD9CM|PT|84.64|Insertion of partial spinal disc prosthesis, lumbosacral
C1455930|ICD9CM|AB|84.64|Ins part disc pros lumb
C1455934|ICD9CM|PT|84.65|Insertion of total spinal disc prosthesis, lumbosacral
C1455934|ICD9CM|AB|84.65|Ins totl disc pros lumb
C1455938|ICD9CM|PT|84.66|Revision or replacement of artificial spinal disc prosthesis, cervical
C1455938|ICD9CM|AB|84.66|Revise disc prost cerv
C1455942|ICD9CM|PT|84.67|Revision or replacement of artificial spinal disc prosthesis, thoracic
C1455942|ICD9CM|AB|84.67|Revise disc prost thora
C1455946|ICD9CM|PT|84.68|Revision or replacement of artificial spinal disc prosthesis, lumbosacral
C1455946|ICD9CM|AB|84.68|Revise disc prosth lumb
C1455950|ICD9CM|PT|84.69|Revision or replacement of artificial spinal disc prosthesis, not otherwise specified
C1455950|ICD9CM|AB|84.69|Revise disc prosth NOS
C1455954|ICD9CM|HT|84.6|Replacement of spinal disc
C1455955|ICD9CM|PT|86.05|Incision with removal of foreign body or device from skin and subcutaneous tissue
C1455955|ICD9CM|AB|86.05|Removal fb/dev from skin
C1455966|ICD9CM|PT|86.96|Insertion or replacement of other neurostimulator pulse generator
C1455966|ICD9CM|AB|86.96|Insert/repl oth neurost
C1455968|ICD9CM|PT|V01.71|Contact with or exposure to varicella
C1455968|ICD9CM|AB|V01.71|Varicella contact/exp
C1455969|ICD9CM|PT|V01.83|Contact with or exposure to escherichia coli (E. coli)
C1455969|ICD9CM|AB|V01.83|E. coli contact/exp
C1455970|ICD9CM|PT|V01.84|Contact with or exposure to meningococcus
C1455970|ICD9CM|AB|V01.84|Meningococcus contact
C1455974|ICD9CM|PT|V46.11|Dependence on respirator, status
C1455974|ICD9CM|AB|V46.11|Respirator depend status
C1455975|ICD9CM|PT|V46.12|Encounter for respirator dependence during power failure
C1455975|ICD9CM|AB|V46.12|Resp depend-powr failure
C1455976|ICD9CM|PT|V49.83|Awaiting organ transplant status
C1455976|ICD9CM|AB|V49.83|Await organ transplnt st
C1455977|ICD9CM|PT|V58.44|Aftercare following organ transplant
C1455977|ICD9CM|AB|V58.44|Aftercare organ transplt
C1455979|ICD9CM|PT|V58.67|Long-term (current) use of insulin
C1455979|ICD9CM|AB|V58.67|Long-term use of insulin
C1455980|ICD9CM|AB|V69.4|Lack of adequate sleep
C1455980|ICD9CM|PT|V69.4|Lack of adequate sleep
C1455982|ICD9CM|PT|V72.31|Routine gynecological examination
C1455982|ICD9CM|AB|V72.31|Routine gyn examination
C1455985|ICD9CM|PT|V72.32|Encounter for Papanicolaou cervical smear to confirm findings of recent normal smear following initial abnormal smear
C1455985|ICD9CM|AB|V72.32|Pap smear confirmation
C1455986|ICD9CM|HT|V72.3|Special investigations and examinations - Gynecological examination
C1455988|ICD9CM|PT|V72.41|Pregnancy examination or test, negative result
C1455988|ICD9CM|AB|V72.41|Pregnancy test negative
C1455989|ICD9CM|HT|V72.4|Pregnancy examination or test
C1455990|ICD9CM|PT|V84.01|Genetic susceptibility to malignant neoplasm of breast
C1455990|ICD9CM|AB|V84.01|Genetc sus mal neo brest
C1455991|ICD9CM|PT|V84.02|Genetic susceptibility to malignant neoplasm of ovary
C1455991|ICD9CM|AB|V84.02|Genetc sus mal neo ovary
C1455992|ICD9CM|PT|V84.03|Genetic susceptibility to malignant neoplasm of prostate
C1455992|ICD9CM|AB|V84.03|Genetc sus mal neo prost
C1455993|ICD9CM|PT|V84.04|Genetic susceptibility to malignant neoplasm of endometrium
C1455993|ICD9CM|AB|V84.04|Genetc susc mal neo endo
C1455994|ICD9CM|PT|V84.09|Genetic susceptibility to other malignant neoplasm
C1455994|ICD9CM|AB|V84.09|Genetic susc mal neo NEC
C1455995|ICD9CM|HT|V84.0|Genetic susceptibility to malignant neoplasm
C1455996|ICD9CM|HT|V84.8|Genetic susceptibility to other disease
C1455996|ICD9CM|PT|V84.89|Genetic susceptibility to other disease
C1455996|ICD9CM|AB|V84.89|Genetic suscept dis NEC
C1456000|ICD9CM|PT|00.16|Pressurized treatment of venous bypass graft [conduit] with pharmaceutical substance
C1456000|ICD9CM|AB|00.16|Pressurized treat graft
C1456003|ICD9CM|PT|00.17|Infusion of vasopressor agent
C1456003|ICD9CM|AB|00.17|Infusion of vasopressor
C1456004|ICD9CM|PT|00.21|Intravascular imaging of extracranial cerebral vessels
C1456004|ICD9CM|AB|00.21|IVUS extracran cereb ves
C1456007|ICD9CM|PT|00.22|Intravascular imaging of intrathoracic vessels
C1456007|ICD9CM|AB|00.22|IVUS intrathoracic ves
C1456012|ICD9CM|PT|00.23|Intravascular imaging of peripheral vessels
C1456012|ICD9CM|AB|00.23|IVUS peripheral vessels
C1456016|ICD9CM|PT|00.24|Intravascular imaging of coronary vessels
C1456016|ICD9CM|AB|00.24|IVUS coronary vessels
C1456018|ICD9CM|PT|00.25|Intravascular imaging of renal vessels
C1456018|ICD9CM|AB|00.25|IVUS renal vessels
C1456021|ICD9CM|PT|00.28|Intravascular imaging, other specified vessel(s)
C1456021|ICD9CM|AB|00.28|Intravascul imaging NEC
C1456022|ICD9CM|PT|00.29|Intravascular imaging, unspecified vessel(s)
C1456022|ICD9CM|AB|00.29|Intravascul imaging NOS
C1456023|ICD9CM|HT|00.2|Intravascular imaging of blood vessels
C1456026|ICD9CM|PT|00.31|Computer assisted surgery with CT/CTA
C1456026|ICD9CM|AB|00.31|CAS w CT/CTA
C1456027|ICD9CM|PT|00.32|Computer assisted surgery with MR/MRA
C1456027|ICD9CM|AB|00.32|CAS w MR/MRA
C1456028|ICD9CM|PT|00.33|Computer assisted surgery with fluoroscopy
C1456028|ICD9CM|AB|00.33|CAS w fluoroscopy
C1456029|ICD9CM|PT|00.34|Imageless computer assisted surgery
C1456029|ICD9CM|AB|00.34|Imageless comp asst surg
C1456030|ICD9CM|PT|00.35|Computer assisted surgery with multiple datasets
C1456030|ICD9CM|AB|00.35|CAS w multiple datasets
C1456031|ICD9CM|PT|00.39|Other computer assisted surgery
C1456031|ICD9CM|AB|00.39|Other CAS
C1456032|ICD9CM|HT|00.3|Computer assisted surgery [CAS]
C1456042|ICD9CM|PT|00.62|Percutaneous angioplasty of intracranial vessel(s)
C1456042|ICD9CM|AB|00.62|Perc angio intracran ves
C1456043|ICD9CM|PT|00.63|Percutaneous insertion of carotid artery stent(s)
C1456043|ICD9CM|AB|00.63|Perc ins carotid stent
C1456045|ICD9CM|PT|00.64|Percutaneous insertion of other extracranial artery stent(s)
C1456045|ICD9CM|AB|00.64|Perc ins extracran stent
C1456048|ICD9CM|PT|00.65|Percutaneous insertion of intracranial vascular stent(s)
C1456048|ICD9CM|AB|00.65|Perc ins intracran stent
C1456049|ICD9CM|PT|00.91|Transplant from live related donor
C1456049|ICD9CM|AB|00.91|Trnsplnt live rel donor
C1456050|ICD9CM|PT|00.92|Transplant from live non-related donor
C1456050|ICD9CM|AB|00.92|Trnsplnt live nonrel don
C1456051|ICD9CM|PT|00.93|Transplant from cadaver
C1456051|ICD9CM|AB|00.93|Transplant cadaver donor
C1456052|ICD9CM|HT|00.9|Other procedures and interventions
C1456053|ICD9CM|PT|01.22|Removal of intracranial neurostimulator lead(s)
C1456053|ICD9CM|AB|01.22|Removal brain stim lead
C1456059|ICD9CM|PT|629.21|Female genital mutilation Type I status
C1456059|ICD9CM|AB|629.21|Genital mutilatn type I
C1456061|ICD9CM|PT|629.22|Female genital mutilation Type II status
C1456061|ICD9CM|AB|629.22|Genital mutilatn type II
C1456063|ICD9CM|PT|629.23|Female genital mutilation Type III status
C1456063|ICD9CM|AB|629.23|Genital muilatn type III
C1456066|ICD9CM|PT|477.2|Allergic rhinitis due to animal (cat) (dog) hair and dander
C1456066|ICD9CM|AB|477.2|Allerg rhinitis-cat/dog
C1456074|ICD9CM|PT|37.66|Insertion of implantable heart assist system
C1456074|ICD9CM|AB|37.66|Implantable hrt assist
C1456082|ICD9CM|PT|37.68|Insertion of percutaneous external heart assist device
C1456082|ICD9CM|AB|37.68|Percutan hrt assist syst
C1456086|ICD9CM|HT|37.6|Implantation of heart and circulatory assist system(s)
C1456087|ICD9CM|PT|37.90|Insertion of left atrial appendage device
C1456087|ICD9CM|AB|37.90|Ins left atr append dev
C1456093|ICD9CM|PT|39.50|Angioplasty of other non-coronary vessel(s)
C1456093|ICD9CM|AB|39.50|Angio oth non-coronary
C1456094|ICD9CM|PT|41.08|Allogeneic hematopoietic stem cell transplant with purging
C1456094|ICD9CM|AB|41.08|Allo hem stem ct w purg
C1456095|ICD9CM|PT|414.07|Coronary atherosclerosis of bypass graft (artery) (vein) of transplanted heart
C1456095|ICD9CM|AB|414.07|Cor ath bps graft tp hrt
C1456097|ICD9CM|PT|44.67|Laparoscopic procedures for creation of esophagogastric sphincteric competence
C1456097|ICD9CM|AB|44.67|Lap creat esoph sphinct
C1456099|ICD9CM|PT|44.68|Laparoscopic gastroplasty
C1456099|ICD9CM|AB|44.68|Laparoscop gastroplasty
C1456102|ICD9CM|PT|44.95|Laparoscopic gastric restrictive procedure
C1456102|ICD9CM|AB|44.95|Lap gastric restric proc
C1456104|ICD9CM|PT|44.96|Laparoscopic revision of gastric restrictive procedure
C1456104|ICD9CM|AB|44.96|Lap rev gast restri proc
C1456107|ICD9CM|PT|44.97|Laparoscopic removal of gastric restrictive device(s)
C1456107|ICD9CM|AB|44.97|Lap rem gast restric dev
C1456111|ICD9CM|PT|44.98|(Laparoscopic) adjustment of size of adjustable gastric restrictive device
C1456111|ICD9CM|AB|44.98|Adjust gast restrict dev
C1456114|ICD9CM|PT|692.84|Contact dermatitis and other eczema due to animal (cat) (dog) dander
C1456114|ICD9CM|AB|692.84|Contact drmatitis-animal
C1456131|ICD9CM|PT|491.22|Obstructive chronic bronchitis with acute bronchitis
C1456131|ICD9CM|AB|491.22|Obs chr bronc w ac bronc
C1456132|ICD9CM|PT|705.21|Primary focal hyperhidrosis
C1456132|ICD9CM|AB|705.21|Primary focal hyprhidros
C1456136|ICD9CM|PT|705.22|Secondary focal hyperhidrosis
C1456136|ICD9CM|AB|705.22|Sec focal hyperhidrosis
C1456139|ICD9CM|PT|707.02|Pressure ulcer, upper back
C1456139|ICD9CM|AB|707.02|Pressure ulcer, upr back
C1456141|ICD9CM|AB|707.03|Pressure ulcer, low back
C1456141|ICD9CM|PT|707.03|Pressure ulcer, lower back
C1456142|ICD9CM|PT|707.09|Pressure ulcer, other site
C1456142|ICD9CM|AB|707.09|Pressure ulcer, site NEC
C1456144|ICD9CM|PT|521.06|Dental caries pit and fissure
C1456144|ICD9CM|AB|521.06|Dentl caries-pit/fissure
C1456145|ICD9CM|PT|521.07|Dental caries of smooth surface
C1456145|ICD9CM|AB|521.07|Dentl caries-smooth surf
C1456147|ICD9CM|PT|521.10|Excessive attrition, unspecified
C1456147|ICD9CM|AB|521.10|Excessive attrition NOS
C1456148|ICD9CM|PT|521.11|Excessive attrition, limited to enamel
C1456148|ICD9CM|AB|521.11|Excess attrition-enamel
C1456149|ICD9CM|PT|521.12|Excessive attrition, extending into dentine
C1456149|ICD9CM|AB|521.12|Excess attrition-dentine
C1456150|ICD9CM|PT|521.13|Excessive attrition, extending into pulp
C1456150|ICD9CM|AB|521.13|Excessive attrition-pulp
C1456151|ICD9CM|PT|521.14|Excessive attrition, localized
C1456151|ICD9CM|AB|521.14|Excess attrition-local
C1456152|ICD9CM|PT|521.15|Excessive attrition, generalized
C1456152|ICD9CM|AB|521.15|Excess attrition-general
C1456153|ICD9CM|HT|521.1|Excessive dental attrition [approximal wear] [occlusal wear]
C1456155|ICD9CM|PT|521.21|Abrasion, limited to enamel
C1456155|ICD9CM|AB|521.21|Abrasion-enamel
C1456156|ICD9CM|PT|521.22|Abrasion, extending into dentine
C1456156|ICD9CM|AB|521.22|Abrasion-dentine
C1456157|ICD9CM|PT|521.23|Abrasion, extending into pulp
C1456157|ICD9CM|AB|521.23|Abrasion-pulp
C1456158|ICD9CM|PT|521.24|Abrasion, localized
C1456158|ICD9CM|AB|521.24|Abrasion-localized
C1456159|ICD9CM|PT|521.25|Abrasion, generalized
C1456159|ICD9CM|AB|521.25|Abrasion-generalized
C1456160|ICD9CM|AB|521.30|Erosion NOS
C1456160|ICD9CM|PT|521.30|Erosion, unspecified
C1456162|ICD9CM|PT|521.32|Erosion, extending into dentine
C1456162|ICD9CM|AB|521.32|Erosion-dentine
C1456163|ICD9CM|PT|521.33|Erosion, extending into pulp
C1456163|ICD9CM|AB|521.33|Erosion-pulp
C1456164|ICD9CM|PT|521.34|Erosion, localized
C1456164|ICD9CM|AB|521.34|Erosion-localized
C1456165|ICD9CM|AB|521.35|Erosion-generalized
C1456165|ICD9CM|PT|521.35|Erosion, generalized
C1456166|ICD9CM|PT|521.40|Pathological resorption, unspecified
C1456166|ICD9CM|AB|521.40|Path resorption NOS
C1456167|ICD9CM|PT|521.41|Pathological resorption, internal
C1456167|ICD9CM|AB|521.41|Path resorption-internal
C1456169|ICD9CM|PT|521.49|Other pathological resorption
C1456169|ICD9CM|AB|521.49|Path resorption NEC
C1456170|ICD9CM|PT|521.7|Intrinsic posteruptive color changes
C1456170|ICD9CM|AB|521.7|Intrin posteruptv color
C1456171|ICD9CM|PT|523.21|Gingival recession, minimal
C1456171|ICD9CM|AB|523.21|Gingival recess-minimal
C1456172|ICD9CM|PT|523.22|Gingival recession, moderate
C1456172|ICD9CM|AB|523.22|Gingival recess-moderate
C1456173|ICD9CM|PT|523.23|Gingival recession, severe
C1456173|ICD9CM|AB|523.23|Gingival recess-severe
C1456175|ICD9CM|PT|524.07|Excessive tuberosity of jaw
C1456175|ICD9CM|AB|524.07|Excessive tuberosity-jaw
C1456181|ICD9CM|PT|524.25|Open posterior occlusal relationship
C1456181|ICD9CM|AB|524.25|Open posterior occlusion
C1456182|ICD9CM|PT|524.26|Excessive horizontal overlap
C1456182|ICD9CM|AB|524.26|Excess horizontl overlap
C1456183|ICD9CM|AB|524.27|Reverse articulation
C1456183|ICD9CM|PT|524.27|Reverse articulation
C1456186|ICD9CM|PT|524.28|Anomalies of interarch distance
C1456186|ICD9CM|AB|524.28|Anom interarch distance
C1456189|ICD9CM|PT|524.29|Other anomalies of dental arch relationship
C1456189|ICD9CM|AB|524.29|Anomaly dental arch NEC
C1456191|ICD9CM|PT|524.32|Excessive spacing of teeth
C1456191|ICD9CM|AB|524.32|Excessive spacing-teeth
C1456192|ICD9CM|PT|524.33|Horizontal displacement of teeth
C1456192|ICD9CM|AB|524.33|Horizontl displace-teeth
C1456194|ICD9CM|PT|524.34|Vertical displacement of teeth
C1456194|ICD9CM|AB|524.34|Vertical displace-teeth
C1456197|ICD9CM|PT|524.36|Insufficient interocclusal distance of teeth (ridge)
C1456197|ICD9CM|AB|524.36|Insuf interocclusl-teeth
C1456198|ICD9CM|PT|524.37|Excessive interocclusal distance of teeth
C1456198|ICD9CM|AB|524.37|Exces interocclusl-teeth
C1456200|ICD9CM|PT|524.39|Other anomalies of tooth position
C1456200|ICD9CM|AB|524.39|Tooth position anom NEC
C1456201|ICD9CM|HT|524.3|Anomalies of tooth position of fully erupted teeth
C1456203|ICD9CM|PT|524.53|Deviation in opening and closing of the mandible
C1456203|ICD9CM|AB|524.53|Dev open/close mandible
C1456205|ICD9CM|PT|524.55|Centric occlusion maximum intercuspation discrepancy
C1456205|ICD9CM|AB|524.55|Centric occl intrcsp dis
C1456207|ICD9CM|PT|524.57|Lack of posterior occlusal support
C1456207|ICD9CM|AB|524.57|Lack post occlsl support
C1456208|ICD9CM|PT|524.59|Other dentofacial functional abnormalities
C1456208|ICD9CM|AB|524.59|Dentofac funct abnor NEC
C1456213|ICD9CM|PT|524.64|Temporomandibular joint sounds on opening and/or closing the jaw
C1456213|ICD9CM|AB|524.64|TMJ sounds opn/close jaw
C1456214|ICD9CM|PT|524.75|Vertical displacement of alveolus and teeth
C1456214|ICD9CM|AB|524.75|Vertical displace teeth
C1456216|ICD9CM|AB|524.76|Occlusal plane deviation
C1456216|ICD9CM|PT|524.76|Occlusal plane deviation
C1456217|ICD9CM|PT|524.81|Anterior soft tissue impingement
C1456217|ICD9CM|AB|524.81|Anterior soft tiss impg
C1456218|ICD9CM|PT|524.82|Posterior soft tissue impingement
C1456218|ICD9CM|AB|524.82|Posterior soft tiss impg
C1456219|ICD9CM|PT|525.20|Unspecified atrophy of edentulous alveolar ridge
C1456219|ICD9CM|AB|525.20|Atrophy alvlar ridge NOS
C1456221|ICD9CM|AB|525.21|Atrophy mandible-minimal
C1456221|ICD9CM|PT|525.21|Minimal atrophy of the mandible
C1456222|ICD9CM|PT|525.22|Moderate atrophy of the mandible
C1456222|ICD9CM|AB|525.22|Atrophy mandible-modrate
C1456223|ICD9CM|AB|525.23|Atrophy mandible-severe
C1456223|ICD9CM|PT|525.23|Severe atrophy of the mandible
C1456224|ICD9CM|AB|525.24|Atrophy maxilla-minimal
C1456224|ICD9CM|PT|525.24|Minimal atrophy of the maxilla
C1456225|ICD9CM|AB|525.25|Atrophy maxilla-moderate
C1456225|ICD9CM|PT|525.25|Moderate atrophy of the maxilla
C1456226|ICD9CM|AB|525.26|Atrophy maxilla-severe
C1456226|ICD9CM|PT|525.26|Severe atrophy of the maxilla
C1456227|ICD9CM|PT|528.71|Minimal keratinized residual ridge mucosa
C1456227|ICD9CM|AB|528.71|Keratin ridge mucosa-min
C1456228|ICD9CM|PT|528.72|Excessive keratinized residual ridge mucosa
C1456228|ICD9CM|AB|528.72|Keratin ridge muc-excess
C1456233|ICD9CM|AB|530.86|Esophagostomy infection
C1456233|ICD9CM|PT|530.86|Infection of esophagostomy
C1456234|ICD9CM|PT|530.87|Mechanical complication of esophagostomy
C1456234|ICD9CM|AB|530.87|Mech comp esophagostomy
C1456238|ICD9CM|PT|03.93|Implantation or replacement of spinal neurostimulator lead(s)
C1456238|ICD9CM|AB|03.93|Imp/repl spine stim lead
C1456239|ICD9CM|PT|03.94|Removal of spinal neurostimulator lead(s)
C1456239|ICD9CM|AB|03.94|Removal spine stim lead
C1456240|ICD9CM|PT|347.00|Narcolepsy, without cataplexy
C1456240|ICD9CM|AB|347.00|Narcolepsy w/o cataplexy
C1456241|ICD9CM|PT|347.10|Narcolepsy in conditions classified elsewhere, without cataplexy
C1456241|ICD9CM|AB|347.10|Narclpsy w/o cat oth dis
C1456242|ICD9CM|PT|347.11|Narcolepsy in conditions classified elsewhere, with cataplexy
C1456242|ICD9CM|AB|347.11|Narcolepsy w cat oth dis
C1456243|ICD9CM|HT|347.1|Narcolepsy in conditions classified elsewhere
C1456244|ICD9CM|PT|04.92|Implantation or replacement of peripheral neurostimulator lead(s)
C1456244|ICD9CM|AB|04.92|Imp/repl peri stim lead
C1456245|ICD9CM|PT|04.93|Removal of peripheral neurostimulator lead(s)
C1456245|ICD9CM|AB|04.93|Removal peri stim lead
C1456246|ICD9CM|AB|041.82|Bacteroides fragilis
C1456246|ICD9CM|PT|041.82|Bacteroides fragilis
C1456247|ICD9CM|PT|618.00|Unspecified prolapse of vaginal walls
C1456247|ICD9CM|AB|618.00|Vaginal wall prolpse NOS
C1456248|ICD9CM|AB|618.01|Cystocele, midline
C1456248|ICD9CM|PT|618.01|Cystocele, midline
C1456251|ICD9CM|AB|618.05|Perineocele
C1456251|ICD9CM|PT|618.05|Perineocele
C1456252|ICD9CM|PT|618.09|Other prolapse of vaginal walls without mention of uterine prolapse
C1456252|ICD9CM|AB|618.09|Cystourethrocele
C1456253|ICD9CM|PT|618.81|Incompetence or weakening of pubocervical tissue
C1456253|ICD9CM|AB|618.81|Incomptnce pubocerv tiss
C1456254|ICD9CM|PT|618.82|Incompetence or weakening of rectovaginal tissue
C1456254|ICD9CM|AB|618.82|Incomptnce rectovag tiss
C1456255|ICD9CM|AB|618.83|Pelvic muscle wasting
C1456255|ICD9CM|PT|618.83|Pelvic muscle wasting
C1456259|ICD9CM|PT|066.42|West Nile Fever with other neurologic manifestation
C1456259|ICD9CM|AB|066.42|West Nile neuro man NEC
C1456260|ICD9CM|PT|066.49|West Nile Fever with other complications
C1456260|ICD9CM|AB|066.49|West Nile w complic NEC
C1456261|ICD9CM|PT|070.41|Acute hepatitis C with hepatic coma
C1456261|ICD9CM|AB|070.41|Hpt C acute w hepat Coma
C1456262|ICD9CM|PT|070.51|Acute hepatitis C without mention of hepatic coma
C1456262|ICD9CM|AB|070.51|Hpt C acute wo hpat coma
C1456263|ICD9CM|PT|070.70|Unspecified viral hepatitis C without hepatic coma
C1456263|ICD9CM|AB|070.70|Hpt C w/o hepat coma NOS
C1456265|ICD9CM|PT|070.71|Unspecified viral hepatitis C with hepatic coma
C1456265|ICD9CM|AB|070.71|Hpt C w hepatic coma NOS
C1456268|ICD9CM|PT|252.02|Secondary hyperparathyroidism, non-renal
C1456268|ICD9CM|AB|252.02|Sec hyprprthyrd nonrenal
C1456269|ICD9CM|PT|27.64|Insertion of palatal implant
C1456269|ICD9CM|AB|27.64|Insert palatal implant
C1456270|ICD9CM|PT|277.85|Disorders of fatty acid oxidation
C1456270|ICD9CM|AB|277.85|Disorders acid oxidation
C1456275|ICD9CM|PT|277.87|Disorders of mitochondrial metabolism
C1456275|ICD9CM|AB|277.87|Dis mitochondrial metab
C1456282|ICD9CM|PT|289.82|Secondary hypercoagulable state
C1456282|ICD9CM|AB|289.82|Sec hypercoagulable st
C1456283|ICD9CM|PT|291.89|Other alcohol-induced mental disorders
C1456283|ICD9CM|HT|291.8|Other specified alcohol-induced mental disorders
C1456283|ICD9CM|AB|291.89|Alcohol mental disor NEC
C1456285|ICD9CM|HT|291|Alcohol-induced mental disorders
C1456286|ICD9CM|PT|292.11|Drug-induced psychotic disorder with delusions
C1456286|ICD9CM|AB|292.11|Drug psych disor w delus
C1456288|ICD9CM|PT|292.82|Drug-induced persisting dementia
C1456288|ICD9CM|AB|292.82|Drug persisting dementia
C1456289|ICD9CM|PT|292.83|Drug-induced persisting amnestic disorder
C1456289|ICD9CM|AB|292.83|Drug persist amnestc dis
C1456292|ICD9CM|PT|292.85|Drug induced sleep disorders
C1456292|ICD9CM|AB|292.85|Drug induced sleep disor
C1456296|ICD9CM|PT|293.0|Delirium due to conditions classified elsewhere
C1456296|ICD9CM|AB|293.0|Delirium d/t other cond
C1456297|ICD9CM|PT|293.81|Psychotic disorder with delusions in conditions classified elsewhere
C1456297|ICD9CM|AB|293.81|Psy dis w delus oth dis
C1456298|ICD9CM|PT|293.83|Mood disorder in conditions classified elsewhere
C1456298|ICD9CM|AB|293.83|Mood disorder other dis
C1456299|ICD9CM|PT|293.84|Anxiety disorder in conditions classified elsewhere
C1456299|ICD9CM|AB|293.84|Anxiety disorder oth dis
C1456301|ICD9CM|HT|293.8|Other specified transient mental disorders due to conditions classified elsewhere
C1456302|ICD9CM|PT|293.9|Unspecified transient mental disorder in conditions classified elsewhere
C1456302|ICD9CM|AB|293.9|Transient mental dis NOS
C1456303|ICD9CM|HT|293|Transient mental disorders due to conditions classified elsewhere
C1456304|ICD9CM|HT|296.4|Bipolar I disorder, most recent episode (or current) manic
C1456305|ICD9CM|HT|296.5|Bipolar I disorder, most recent episode (or current) depressed
C1456306|ICD9CM|HT|296.6|Bipolar I disorder, most recent episode (or current) mixed
C1456307|ICD9CM|PT|296.7|Bipolar I disorder, most recent episode (or current) unspecified
C1456307|ICD9CM|AB|296.7|Bipolor I current NOS
C1456308|ICD9CM|PT|296.89|Other bipolar disorders
C1456308|ICD9CM|AB|296.89|Bipolar disorder NEC
C1456309|ICD9CM|HT|296.8|Other and unspecified bipolar disorders
C1456310|ICD9CM|PT|296.99|Other specified episodic mood disorder
C1456310|ICD9CM|AB|296.99|Episodic mood disord NEC
C1456311|ICD9CM|HT|296.9|Other and unspecified episodic mood disorder
C1456313|ICD9CM|HT|299.8|Other specified pervasive developmental disorders
C1456314|ICD9CM|HT|300.1|Dissociative, conversion and factitious disorders
C1456315|ICD9CM|PT|300.29|Other isolated or specific phobias
C1456315|ICD9CM|AB|300.29|Isolated/spec phobia NEC
C1456316|ICD9CM|HT|300|Anxiety, dissociative and somatoform disorders
C1456319|ICD9CM|AB|302.74|Male orgasmic disorder
C1456319|ICD9CM|PT|302.74|Male orgasmic disorder
C1456321|ICD9CM|PT|307.89|Other pain disorders related to psychological factors
C1456321|ICD9CM|AB|307.89|Psychogenic pain NEC
C1456322|ICD9CM|HT|307.8|Pain disorders related to psychological factors
C1456323|ICD9CM|PT|310.1|Personality change due to conditions classified elsewhere
C1456323|ICD9CM|AB|310.1|Personality chg oth dis
C1456324|ICD9CM|HT|310|Specific nonpsychotic mental disorders due to brain damage
C1456326|ICD9CM|AB|313.23|Selective mutism
C1456326|ICD9CM|PT|313.23|Selective mutism
C1456424|ICD9CM|PT|751.60|Unspecified anomaly of gallbladder, bile ducts, and liver
C1456424|ICD9CM|AB|751.60|Biliary & liver anom NOS
C1456428|ICD9CM|PT|294.9|Unspecified persistent mental disorders due to conditions classified elsewhere
C1456428|ICD9CM|AB|294.9|Mental disor NOS oth dis
C1456434|ICD9CM|HT|296|Episodic mood disorders
C1456434|ICD9CM|PT|296.90|Unspecified episodic mood disorder
C1456434|ICD9CM|AB|296.90|Episodic mood disord NOS
C1456732|ICD9CM|PT|292.12|Drug-induced psychotic disorder with hallucinations
C1456732|ICD9CM|AB|292.12|Drug psy dis w hallucin
C1456783|ICD9CM|HT|297|Paranoid states (Delusional disorders)
C1456786|ICD9CM|AB|297.9|Paranoid state NOS
C1456786|ICD9CM|PT|297.9|Unspecified paranoid state
C1456876|ICD9CM|HT|635|Legally induced abortion
C1457882|ICD9CM|PT|96.58|Irrigation of wound catheter
C1457882|ICD9CM|AB|96.58|Wound catheter irrigat
C1457887|ICD9CM|HT|780-789.99|SYMPTOMS
C1457889|ICD9CM|PT|290.9|Unspecified senile psychotic condition
C1457889|ICD9CM|AB|290.9|Senile psychot cond NOS
C1457897|ICD9CM|PT|279.04|Congenital hypogammaglobulinemia
C1457897|ICD9CM|AB|279.04|Cong hypogammaglobulinem
C1504340|ICD9CM|HT|349.3|Dural tear
C1504394|ICD9CM|PT|33.42|Closure of bronchial fistula
C1504394|ICD9CM|AB|33.42|Bronchial fistula clos
C1504514|ICD9CM|PT|058.82|Human herpesvirus 7 infection
C1504514|ICD9CM|AB|058.82|Human herpesvirus 7 infc
C1510449|ICD9CM|HT|364.1|Chronic iridocyclitis
C1510449|ICD9CM|PT|364.10|Chronic iridocyclitis, unspecified
C1510449|ICD9CM|AB|364.10|Chr iridocyclitis NOS
C1510455|ICD9CM|AB|755.55|Acrocephalosyndactyly
C1510455|ICD9CM|PT|755.55|Acrocephalosyndactyly
C1510471|ICD9CM|AB|269.2|Vitamin Deficiency NOS
C1510471|ICD9CM|PT|269.2|Unspecified vitamin deficiency
C1510472|ICD9CM|HT|304|Drug dependence
C1510472|ICD9CM|HT|304.9|Unspecified drug dependence
C1510475|ICD9CM|HT|562|Diverticula of intestine
C1510479|ICD9CM|AB|353.5|Neuralgic amyotrophy
C1510479|ICD9CM|PT|353.5|Neuralgic amyotrophy
C1510504|ICD9CM|HT|764.2|Fetal malnutrition without mention of "light-for-dates"
C1527169|ICD9CM|HT|V59|Donors
C1527344|ICD9CM|AB|784.42|Dysphonia
C1527344|ICD9CM|PT|784.42|Dysphonia
C1527368|ICD9CM|AB|101|Vincent's angina
C1527368|ICD9CM|PT|101|Vincent's angina
C1532320|ICD9CM|PT|V16.42|Family history of malignant neoplasm of prostate
C1532320|ICD9CM|AB|V16.42|Fm hx prostate malig
C1532368|ICD9CM|PT|205.12|Chronic myeloid leukemia, in relapse
C1532368|ICD9CM|AB|205.12|Chr myel leuk in relapse
C1532669|ICD9CM|HT|552.2|Ventral hernia with obstruction
C1532669|ICD9CM|PT|552.20|Ventral, unspecified, hernia with obstruction
C1532669|ICD9CM|AB|552.20|Obstr ventral hernia NOS
C1533166|ICD9CM|PT|967.3|Poisoning by bromine compounds
C1533166|ICD9CM|AB|967.3|Poisoning-bromine compnd
C1533173|ICD9CM|PT|09.82|Conjunctivocystorhinostomy
C1533173|ICD9CM|AB|09.82|Conjunctivocystorhinost
C1533614|ICD9CM|HT|30-34.99|OPERATIONS ON THE RESPIRATORY SYSTEM
C1533618|ICD9CM|AB|958.1|Fat embolism
C1533618|ICD9CM|PT|958.1|Fat embolism
C1533626|ICD9CM|HT|647.3|Tuberculosis complicating pregnancy, childbirth, or the puerperium
C1533651|ICD9CM|HT|279.1|Deficiency of cell-mediated immunity
C1533659|ICD9CM|HT|361|Retinal detachments and defects
C1533661|ICD9CM|PT|80.23|Arthroscopy, wrist
C1533661|ICD9CM|AB|80.23|Wrist arthroscopy
C1533664|ICD9CM|PT|48.41|Soave submucosal resection of rectum
C1533664|ICD9CM|AB|48.41|Soave submuc rect resect
C1533665|ICD9CM|HT|56.8|Repair of ureter
C1533667|ICD9CM|AB|70.76|Hymenorrhaphy
C1533667|ICD9CM|PT|70.76|Hymenorrhaphy
C1533669|ICD9CM|PT|08.11|Biopsy of eyelid
C1533669|ICD9CM|AB|08.11|Eyelid biopsy
C1533670|ICD9CM|PT|08.33|Repair of blepharoptosis by resection or advancement of levator muscle or aponeurosis
C1533670|ICD9CM|AB|08.33|Ptosis rep-levat mus adv
C1533671|ICD9CM|HT|13.6|Other cataract extraction
C1533671|ICD9CM|PT|13.69|Other cataract extraction
C1533671|ICD9CM|AB|13.69|Cataract extraction NEC
C1533672|ICD9CM|HT|E942|Agents primarily affecting the cardiovascular system causing adverse effects in therapeutic use
C1533674|ICD9CM|HT|365.0|Borderline glaucoma [glaucoma suspect]
C1533675|ICD9CM|HT|377|Disorders of optic nerve and visual pathways
C1533675|ICD9CM|PT|377.9|Unspecified disorder of optic nerve and visual pathways
C1533675|ICD9CM|AB|377.9|Optic nerve disorder NOS
C1534555|ICD9CM|PT|93.77|Training in braille or moon
C1534555|ICD9CM|AB|93.77|Braille or moon training
C1535481|ICD9CM|PT|E865.3|Accidental poisoning from berries and seeds
C1535481|ICD9CM|AB|E865.3|Acc poison-berries/seeds
C1535939|ICD9CM|AB|136.3|Pneumocystosis
C1535939|ICD9CM|PT|136.3|Pneumocystosis
C1536114|ICD9CM|PT|338.0|Central pain syndrome
C1536114|ICD9CM|AB|338.0|Central pain syndrome
C1536381|ICD9CM|AB|81.96|Other repair of joint
C1536381|ICD9CM|PT|81.96|Other repair of joint
C1536686|ICD9CM|PT|953.1|Injury to dorsal nerve root
C1536686|ICD9CM|AB|953.1|Dorsal root injury
C1536863|ICD9CM|PT|60.82|Excision of periprostatic tissue
C1536863|ICD9CM|AB|60.82|Periprostatic excision
C1536867|ICD9CM|PT|68.13|Open biopsy of uterus
C1536867|ICD9CM|AB|68.13|Open uterine biopsy
C1536871|ICD9CM|PT|75.62|Repair of current obstetric laceration of rectum and sphincter ani
C1536871|ICD9CM|AB|75.62|Repair ob lac rect/anus
C1541850|ICD9CM|PT|447.0|Arteriovenous fistula, acquired
C1541850|ICD9CM|AB|447.0|Acq arterioven fistula
C1541919|ICD9CM|PT|414.10|Aneurysm of heart (wall)
C1541919|ICD9CM|AB|414.10|Aneurysm of heart
C1541963|CCS|XM|NOCODE|ICD9CM_2005 to CCS2005 Mappings
C1542178|ICD9CM|HT|820-829.99|FRACTURE OF LOWER LIMB
C1542327|ICD9CM|PT|760.71|Alcohol affecting fetus or newborn via placenta or breast milk
C1542327|ICD9CM|AB|760.71|Maternl alc aff NB/fetus
C1561612|MTH|PN|NOCODE|Other diseases of larynx, NEC in ICD9CM
C1561612|ICD9CM|HT|478.7|Other diseases of larynx, not elsewhere classified
C1561612|ICD9CM|PT|478.79|Other diseases of larynx, not elsewhere classified
C1561612|ICD9CM|AB|478.79|Disease of larynx NEC
C1561613|ICD9CM|HT|525.4|Complete edentulism
C1561613|ICD9CM|AB|525.40|Complete edentulism NOS
C1561613|ICD9CM|PT|525.40|Complete edentulism, unspecified
C1561614|ICD9CM|PT|525.41|Complete edentulism, class I
C1561614|ICD9CM|AB|525.41|Comp edentulism,class I
C1561615|ICD9CM|PT|525.42|Complete edentulism, class II
C1561615|ICD9CM|AB|525.42|Comp edentulism,class II
C1561616|ICD9CM|PT|525.43|Complete edentulism, class III
C1561616|ICD9CM|AB|525.43|Comp edentulsm,class III
C1561617|ICD9CM|PT|525.44|Complete edentulism, class IV
C1561617|ICD9CM|AB|525.44|Comp edentulism,class IV
C1561619|ICD9CM|HT|525.5|Partial edentulism
C1561619|ICD9CM|AB|525.50|Partial edentulism NOS
C1561619|ICD9CM|PT|525.50|Partial edentulism, unspecified
C1561620|ICD9CM|PT|525.51|Partial edentulism, class I
C1561620|ICD9CM|AB|525.51|Part edentulism,class I
C1561621|ICD9CM|PT|525.52|Partial edentulism, class II
C1561621|ICD9CM|AB|525.52|Part edentulism,class II
C1561622|ICD9CM|PT|525.53|Partial edentulism, class III
C1561622|ICD9CM|AB|525.53|Part edentulsm,class III
C1561623|ICD9CM|PT|525.54|Partial edentulism, class IV
C1561623|ICD9CM|AB|525.54|Part edentulism,class IV
C1561633|ICD9CM|PT|567.38|Other retroperitoneal abscess
C1561633|ICD9CM|AB|567.38|Retroperiton abscess NEC
C1561634|ICD9CM|PT|567.39|Other retroperitoneal infections
C1561634|ICD9CM|AB|567.39|Retroperiton infect NEC
C1561637|ICD9CM|HT|567|Peritonitis and retroperitoneal infections
C1561638|ICD9CM|PT|585.1|Chronic kidney disease, Stage I
C1561638|ICD9CM|AB|585.1|Chro kidney dis stage I
C1561639|ICD9CM|PT|585.2|Chronic kidney disease, Stage II (mild)
C1561639|ICD9CM|AB|585.2|Chro kidney dis stage II
C1561640|ICD9CM|PT|585.3|Chronic kidney disease, Stage III (moderate)
C1561640|ICD9CM|AB|585.3|Chr kidney dis stage III
C1561641|ICD9CM|PT|585.4|Chronic kidney disease, Stage IV (severe)
C1561641|ICD9CM|AB|585.4|Chr kidney dis stage IV
C1561642|ICD9CM|PT|585.5|Chronic kidney disease, Stage V
C1561642|ICD9CM|AB|585.5|Chron kidney dis stage V
C1561643|ICD9CM|HT|585|Chronic kidney disease (CKD)
C1561643|ICD9CM|PT|585.9|Chronic kidney disease, unspecified
C1561643|ICD9CM|AB|585.9|Chronic kidney dis NOS
C1561646|ICD9CM|PT|599.69|Urinary obstruction, not elsewhere classified
C1561646|ICD9CM|AB|599.69|Urinary obstruction NEC
C1561647|ICD9CM|PT|651.70|Multiple gestation following (elective) fetal reduction, unspecified as to episode of care or not applicable
C1561647|ICD9CM|AB|651.70|Mul gest-fet reduct unsp
C1561648|ICD9CM|PT|651.71|Multiple gestation following (elective) fetal reduction,delivered, with or without mention of antepartum condition
C1561648|ICD9CM|AB|651.71|Mult gest-fet reduct del
C1561649|ICD9CM|PT|651.73|Multiple gestation following (elective) fetal reduction, antepartum condition or complication
C1561649|ICD9CM|AB|651.73|Mul gest-fet reduct ante
C1561650|ICD9CM|HT|651.7|Multiple gestation following (elective) fetal reduction
C1561653|MTH|PN|NOCODE|Other specified adverse effects, NEC in ICD9CM_2014
C1561653|ICD9CM|AB|995.89|Adverse effect NEC
C1561653|ICD9CM|HT|995.8|Other specified adverse effects, not elsewhere classified
C1561653|ICD9CM|PT|995.89|Other specified adverse effects, not elsewhere classified
C1561654|ICD9CM|PT|996.40|Unspecified mechanical complication of internal orthopedic device, implant, and graft
C1561654|ICD9CM|AB|996.40|Cmp int orth dev/gft NOS
C1561655|ICD9CM|PT|996.41|Mechanical loosening of prosthetic joint
C1561655|ICD9CM|AB|996.41|Mech loosening pros jt
C1561661|ICD9CM|PT|996.44|Peri-prosthetic fracture around prosthetic joint
C1561661|ICD9CM|AB|996.44|Periprosthetc fx-pros jt
C1561664|ICD9CM|PT|996.47|Other mechanical complication of prosthetic joint implant
C1561664|ICD9CM|AB|996.47|Mech com pros jt implant
C1561666|ICD9CM|PT|996.49|Other mechanical complication of other internal orthopedic device, implant, and graft
C1561666|ICD9CM|AB|996.49|Mech com orth dev NEC
C1561673|ICD9CM|PT|V46.13|Encounter for weaning from respirator [ventilator]
C1561673|ICD9CM|AB|V46.13|Weaning from respirator
C1561674|ICD9CM|PT|V46.14|Mechanical complication of respirator [ventilator]
C1561674|ICD9CM|AB|V46.14|Mech comp respirator
C1561676|ICD9CM|AB|V49.84|Bed confinement status
C1561676|ICD9CM|PT|V49.84|Bed confinement status
C1561677|ICD9CM|PT|V58.11|Encounter for antineoplastic chemotherapy
C1561677|ICD9CM|AB|V58.11|Antineoplastic chemo enc
C1561678|ICD9CM|PT|V58.12|Encounter for antineoplastic immunotherapy
C1561678|ICD9CM|AB|V58.12|Immunotherapy encounter
C1561680|ICD9CM|PT|V59.71|Egg (oocyte) (ovum) donor, under age 35, anonymous recipient
C1561680|ICD9CM|AB|V59.71|Egg donor age <35 anon
C1561683|ICD9CM|PT|V59.73|Egg (oocyte) (ovum) donor, age 35 and over, anonymous recipient
C1561683|ICD9CM|AB|V59.73|Egg donor age 35+ anon
C1561686|ICD9CM|HT|V59.7|Egg (oocyte) (ovum)
C1561694|ICD9CM|PT|V64.04|Vaccination not carried out because of allergy to vaccine or component
C1561694|ICD9CM|AB|V64.04|No vaccin-allergy to vac
C1561695|ICD9CM|PT|V64.05|Vaccination not carried out because of caregiver refusal
C1561695|ICD9CM|AB|V64.05|No vaccin-caregiv refuse
C1561696|ICD9CM|PT|V64.06|Vaccination not carried out because of patient refusal
C1561696|ICD9CM|AB|V64.06|No vaccination-pt refuse
C1561697|ICD9CM|PT|V64.07|Vaccination not carried out for religious reasons
C1561697|ICD9CM|AB|V64.07|No vaccination-religion
C1561698|ICD9CM|PT|V64.08|Vaccination not carried out because patient had disease being vaccinated against
C1561698|ICD9CM|AB|V64.08|No vaccin-prev disease
C1561709|ICD9CM|PT|V72.86|Encounter for blood typing
C1561709|ICD9CM|AB|V72.86|Blood typing encounter
C1561710|ICD9CM|PT|V85.0|Body Mass Index less than 19, adult
C1561710|ICD9CM|AB|V85.0|BMI less than 19,adult
C1561711|ICD9CM|PT|V85.1|Body Mass Index between 19-24, adult
C1561711|ICD9CM|AB|V85.1|BMI between 19-24,adult
C1561717|ICD9CM|HT|V85.2|Body Mass Index between 25-29, adult
C1561728|ICD9CM|HT|V85.3|Body Mass Index between 30-39, adult
C1561729|ICD9CM|HT|V85.4|Body Mass Index 40 and over, adult
C1561739|ICD9CM|PT|00.40|Procedure on single vessel
C1561739|ICD9CM|AB|00.40|Procedure-one vessel
C1561741|ICD9CM|PT|00.41|Procedure on two vessels
C1561741|ICD9CM|AB|00.41|Procedure-two vessels
C1561742|ICD9CM|PT|00.42|Procedure on three vessels
C1561742|ICD9CM|AB|00.42|Procedure-three vessels
C1561743|ICD9CM|PT|00.43|Procedure on four or more vessels
C1561743|ICD9CM|AB|00.43|Procedure-four+ vessels
C1561744|ICD9CM|PT|00.45|Insertion of one vascular stent
C1561744|ICD9CM|AB|00.45|Insert 1 vascular stent
C1561746|ICD9CM|PT|00.46|Insertion of two vascular stents
C1561746|ICD9CM|AB|00.46|Insert 2 vascular stents
C1561747|ICD9CM|PT|00.47|Insertion of three vascular stents
C1561747|ICD9CM|AB|00.47|Insert 3 vascular stents
C1561748|ICD9CM|PT|00.48|Insertion of four or more vascular stents
C1561748|ICD9CM|AB|00.48|Insert 4+ vasculr stents
C1561749|ICD9CM|HT|00.4|Adjunct Vascular System Procedures
C1561753|ICD9CM|PT|00.70|Revision of hip replacement, both acetabular and femoral components
C1561753|ICD9CM|AB|00.70|Rev hip repl-acetab/fem
C1561755|ICD9CM|PT|00.71|Revision of hip replacement, acetabular component
C1561755|ICD9CM|AB|00.71|Rev hip repl-acetab comp
C1561759|ICD9CM|PT|00.72|Revision of hip replacement, femoral component
C1561759|ICD9CM|AB|00.72|Rev hip repl-fem comp
C1561763|ICD9CM|PT|00.73|Revision of hip replacement, acetabular liner and/or femoral head only
C1561763|ICD9CM|AB|00.73|Rev hip repl-liner/head
C1561767|ICD9CM|HT|00.7|Other hip procedures
C1561768|ICD9CM|PT|00.80|Revision of knee replacement, total (all components)
C1561768|ICD9CM|AB|00.80|Rev knee replacemt-total
C1561770|ICD9CM|PT|00.81|Revision of knee replacement, tibial component
C1561770|ICD9CM|AB|00.81|Rev knee repl-tibia comp
C1561772|ICD9CM|PT|00.82|Revision of knee replacement, femoral component
C1561772|ICD9CM|AB|00.82|Rev knee repl-femur comp
C1561774|ICD9CM|PT|00.83|Revision of knee replacement, patellar component
C1561774|ICD9CM|AB|00.83|Rev knee replace-patella
C1561775|ICD9CM|PT|00.84|Revision of total knee replacement, tibial insert (liner)
C1561775|ICD9CM|AB|00.84|Rev knee repl-tibia lin
C1561781|ICD9CM|PT|760.77|Anticonvulsants affecting fetus or newborn via placenta or breast milk
C1561781|ICD9CM|AB|760.77|Mat anticonv aff NB/fet
C1561786|ICD9CM|PT|760.78|Antimetabolic agents affecting fetus or newborn via placenta or breast milk
C1561786|ICD9CM|AB|760.78|Mat antimetabol aff NB
C1561790|ICD9CM|AB|763.84|Meconium dur del aff NB
C1561790|ICD9CM|PT|763.84|Meconium passage during delivery
C1561791|ICD9CM|PT|770.10|Fetal and newborn aspiration, unspecified
C1561791|ICD9CM|AB|770.10|Fetal & newborn asp NOS
C1561792|ICD9CM|PT|770.11|Meconium aspiration without respiratory symptoms
C1561792|ICD9CM|AB|770.11|Meconium asp wo resp sym
C1561793|ICD9CM|PT|770.12|Meconium aspiration with respiratory symptoms
C1561793|ICD9CM|AB|770.12|Meconium asp w resp symp
C1561794|ICD9CM|PT|770.13|Aspiration of clear amniotic fluid without respiratory symptoms
C1561794|ICD9CM|AB|770.13|Amniotc asp w/o resp sym
C1561796|ICD9CM|PT|770.14|Aspiration of clear amniotic fluid with respiratory symptoms
C1561796|ICD9CM|AB|770.14|Amniotic asp w resp sym
C1561799|ICD9CM|PT|770.15|Aspiration of blood without respiratory symptoms
C1561799|ICD9CM|AB|770.15|Blood asp w/o resp sympt
C1561800|ICD9CM|PT|770.16|Aspiration of blood with respiratory symptoms
C1561800|ICD9CM|AB|770.16|Blood asp w resp sympt
C1561801|ICD9CM|PT|770.17|Other fetal and newborn aspiration without respiratory symptoms
C1561801|ICD9CM|AB|770.17|NB asp w/o resp symp NEC
C1561802|ICD9CM|PT|770.18|Other fetal and newborn aspiration with respiratory symptoms
C1561802|ICD9CM|AB|770.18|NB asp w resp symp NEC
C1561805|ICD9CM|HT|770.1|Fetal and newborn aspiration
C1561806|ICD9CM|PT|770.85|Aspiration of postnatal stomach contents without respiratory symptoms
C1561806|ICD9CM|AB|770.85|Stomch cont asp w/o resp
C1561808|ICD9CM|PT|770.86|Aspiration of postnatal stomach contents with respiratory symptoms
C1561808|ICD9CM|AB|770.86|Stomach cont asp w resp
C1561811|ICD9CM|HT|78.1|Application of external fixator device
C1561813|ICD9CM|PT|780.51|Insomnia with sleep apnea, unspecified
C1561813|ICD9CM|AB|780.51|Insomn w sleep apnea NOS
C1561815|ICD9CM|PT|780.53|Hypersomnia with sleep apnea, unspecified
C1561815|ICD9CM|AB|780.53|Hypersom w slp apnea NOS
C1561817|ICD9CM|PT|780.55|Disruption of 24 hour sleep wake cycle, unspecified
C1561817|ICD9CM|AB|780.55|Irreg sleep-wake rhy NOS
C1561818|ICD9CM|PT|780.58|Sleep related movement disorder, unspecified
C1561818|ICD9CM|AB|780.58|Sleep rel move disor NOS
C1561822|ICD9CM|HT|799.0|Asphyxia and hypoxemia
C1561826|ICD9CM|HT|278.0|Overweight and obesity
C1561827|ICD9CM|HT|278|Overweight, obesity and other hyperalimentation
C1561828|ICD9CM|PT|285.21|Anemia in chronic kidney disease
C1561828|ICD9CM|AB|285.21|Anemia in chr kidney dis
C1561830|ICD9CM|PT|287.30|Primary thrombocytopenia,unspecified
C1561830|ICD9CM|AB|287.30|Prim thrombocytopen NOS
C1561831|ICD9CM|PT|287.33|Congenital and hereditary thrombocytopenic purpura
C1561831|ICD9CM|AB|287.33|Cong/herid thromb purpra
C1561844|ICD9CM|PT|307.45|Circadian rhythm sleep disorder of nonorganic origin
C1561844|ICD9CM|AB|307.45|Nonorganic circadian rhy
C1561849|ICD9CM|PT|327.01|Insomnia due to medical condition classified elsewhere
C1561849|ICD9CM|AB|327.01|Insomnia in other dis
C1561850|ICD9CM|PT|327.02|Insomnia due to mental disorder
C1561850|ICD9CM|AB|327.02|Insomnia dt mental disor
C1561851|ICD9CM|PT|327.09|Other organic insomnia
C1561851|ICD9CM|AB|327.09|Organic insomnia NEC
C1561852|ICD9CM|HT|327.0|Organic disorders of initiating and maintaining sleep [Organic insomnia]
C1561855|ICD9CM|PT|327.12|Idiopathic hypersomnia without long sleep time
C1561855|ICD9CM|AB|327.12|Idio hypersom-no lng slp
C1561857|ICD9CM|PT|327.14|Hypersomnia due to medical condition classified elsewhere
C1561857|ICD9CM|AB|327.14|Hypersomnia in other dis
C1561858|ICD9CM|PT|327.15|Hypersomnia due to mental disorder
C1561858|ICD9CM|AB|327.15|Hypersom dt mental disor
C1561859|ICD9CM|PT|327.19|Other organic hypersomnia
C1561859|ICD9CM|AB|327.19|Organic hypersomnia NEC
C1561860|ICD9CM|HT|327.1|Organic disorder of excessive somnolence [Organic hypersomnia]
C1561861|ICD9CM|HT|327.2|Organic sleep apnea
C1561861|ICD9CM|AB|327.20|Organic sleep apnea NOS
C1561861|ICD9CM|PT|327.20|Organic sleep apnea, unspecified
C1561862|ICD9CM|PT|327.22|High altitude periodic breathing
C1561862|ICD9CM|AB|327.22|High altitude breathing
C1561866|ICD9CM|PT|327.25|Congenital central alveolar hypoventilation syndrome
C1561866|ICD9CM|AB|327.25|Cong cntrl hypovent synd
C1561867|ICD9CM|PT|327.26|Sleep related hypoventilation/hypoxemia in conditions classifiable elsewhere
C1561867|ICD9CM|AB|327.26|Sleep hypovent oth dis
C1561868|ICD9CM|PT|327.27|Central sleep apnea in conditions classified elsewhere
C1561868|ICD9CM|AB|327.27|Cntrl sleep apnea ot dis
C1561869|ICD9CM|PT|327.29|Other organic sleep apnea
C1561869|ICD9CM|AB|327.29|Organic sleep apnea NEC
C1561871|ICD9CM|PT|327.30|Circadian rhythm sleep disorder, unspecified
C1561871|ICD9CM|AB|327.30|Circadian rhym sleep NOS
C1561874|ICD9CM|PT|327.33|Circadian rhythm sleep disorder, irregular sleep-wake type
C1561874|ICD9CM|AB|327.33|Circadian rhym-irreg slp
C1561878|ICD9CM|PT|327.37|Circadian rhythm sleep disorder in conditions classified elsewhere
C1561878|ICD9CM|AB|327.37|Circadian rhym oth dis
C1561879|ICD9CM|PT|327.39|Other circadian rhythm sleep disorder
C1561879|ICD9CM|AB|327.39|Circadian rhym sleep NEC
C1561882|ICD9CM|HT|327.4|Organic parasomnia
C1561882|ICD9CM|AB|327.40|Organic parasomnia NOS
C1561882|ICD9CM|PT|327.40|Organic parasomnia, unspecified
C1561883|ICD9CM|PT|327.43|Recurrent isolated sleep paralysis
C1561883|ICD9CM|AB|327.43|Recurrnt sleep paralysis
C1561885|ICD9CM|PT|327.49|Other organic parasomnia
C1561885|ICD9CM|AB|327.49|Organic parasomnia NEC
C1561888|ICD9CM|AB|327.52|Sleep related leg cramps
C1561888|ICD9CM|PT|327.52|Sleep related leg cramps
C1561889|ICD9CM|PT|327.59|Other organic sleep related movement disorders
C1561889|ICD9CM|AB|327.59|Organic sleep movemt NEC
C1561890|ICD9CM|HT|327.5|Organic sleep related movement disorders
C1561891|ICD9CM|PT|327.8|Other organic sleep disorders
C1561891|ICD9CM|AB|327.8|Sleep organic disord NEC
C1561892|ICD9CM|HT|327|Organic sleep disorders
C1561892|ICD9CM|HT|327-327.99|ORGANIC SLEEP DISORDERS
C1561895|ICD9CM|PT|37.41|Implantation of prosthetic cardiac support device around the heart
C1561895|ICD9CM|AB|37.41|Impl cardiac support dev
C1561900|ICD9CM|PT|37.49|Other repair of heart and pericardium
C1561900|ICD9CM|AB|37.49|Heart/pericard repr NEC
C1561901|ICD9CM|PT|37.79|Revision or relocation of cardiac device pocket
C1561901|ICD9CM|AB|37.79|Rev/reloc card dev pockt
C1561903|ICD9CM|PT|39.73|Endovascular implantation of graft in thoracic aorta
C1561903|ICD9CM|AB|39.73|Endo imp grft thor aorta
C1561927|ICD9CM|PT|81.18|Subtalar joint arthroereisis
C1561927|ICD9CM|AB|81.18|Subtalr jt arthroereisis
C1561928|ICD9CM|HT|81.1|Arthrodesis and arthroereisis of foot and ankle
C1561929|ICD9CM|PT|81.53|Revision of hip replacement, not otherwise specified
C1561929|ICD9CM|AB|81.53|Revise hip replacemt NOS
C1561931|ICD9CM|PT|81.55|Revision of knee replacement, not otherwise specified
C1561931|ICD9CM|AB|81.55|Revise knee replace NOS
C1561932|ICD9CM|PT|84.56|Insertion or replacement of (cement) spacer
C1561932|ICD9CM|AB|84.56|Ins or rep cement spacer
C1561934|ICD9CM|PT|84.57|Removal of (cement) spacer
C1561934|ICD9CM|AB|84.57|Removal of cement spacer
C1561937|ICD9CM|PT|84.71|Application of external fixator device, monoplanar system
C1561937|ICD9CM|AB|84.71|App ext fix dev-monoplan
C1561938|ICD9CM|PT|84.72|Application of external fixator device, ring system
C1561938|ICD9CM|AB|84.72|App ext fix dev-ring sys
C1561941|ICD9CM|PT|84.73|Application of hybrid external fixator device
C1561941|ICD9CM|AB|84.73|App hybrid ext fix dev
C1561943|ICD9CM|HT|84.7|Adjunct codes for external fixator devices
C1561944|ICD9CM|PT|86.94|Insertion or replacement of single array neurostimulator pulse generator, not specified as rechargeable
C1561944|ICD9CM|AB|86.94|Ins/repl single pul gen
C1561946|ICD9CM|PT|86.97|Insertion or replacement of single array rechargeable neurostimulator pulse generator
C1561946|ICD9CM|AB|86.97|Ins/rep 1 pul gen,rechrg
C1561950|ICD9CM|PT|92.20|Infusion of liquid brachytherapy radioisotope
C1561950|ICD9CM|AB|92.20|Inf liquid brachy isotop
C1562427|ICD9CM|PT|282.42|Sickle-cell thalassemia with crisis
C1562427|ICD9CM|AB|282.42|Thlassemia Hb-S w crisis
C1565171|ICD9CM|PT|339.03|Episodic paroxysmal hemicrania
C1565171|ICD9CM|AB|339.03|Episdc paroxyml hemicran
C1576412|ICD9CM|AB|360.43|Hemophthalmos
C1576412|ICD9CM|PT|360.43|Hemophthalmos, except current injury
C1608262|ICD9CM|PT|279.10|Immunodeficiency with predominant T-cell defect, unspecified
C1608262|ICD9CM|AB|279.10|Immundef t-cell def NOS
C1611187|ICD9CM|PT|008.65|Enteritis due to calicivirus
C1611187|ICD9CM|AB|008.65|Enteritis d/t calicivirs
C1611734|ICD9CM|AB|733.45|Aseptic necrosis of jaw
C1611734|ICD9CM|PT|733.45|Aseptic necrosis of bone, jaw
C1621349|ICD9CM|PT|601.4|Prostatitis in diseases classified elsewhere
C1621349|ICD9CM|AB|601.4|Prostatitis in oth dis
C1689951|ICD9CM|PT|330.2|Cerebral degeneration in generalized lipidoses
C1689951|ICD9CM|AB|330.2|Cereb degen in lipidosis
C1691215|ICD9CM|AB|752.61|Hypospadias
C1691215|ICD9CM|PT|752.61|Hypospadias
C1692323|ICD9CM|PT|716.50|Unspecified polyarthropathy or polyarthritis, site unspecified
C1692323|ICD9CM|HT|716.5|Unspecified polyarthropathy or polyarthritis
C1692323|ICD9CM|AB|716.50|Polyarthritis NOS-unspec
C1701940|ICD9CM|PT|997.31|Ventilator associated pneumonia
C1701940|ICD9CM|AB|997.31|Ventltr assoc pneumonia
C1704272|ICD9CM|HT|600.0|Hypertrophy (benign) of prostate
C1704274|ICD9CM|AB|621.5|Intrauterine synechiae
C1704274|ICD9CM|PT|621.5|Intrauterine synechiae
C1704300|ICD9CM|PT|779.6|Termination of pregnancy (fetus)
C1704300|ICD9CM|AB|779.6|Termination of pregnancy
C1704321|ICD9CM|AB|581.3|Minimal change nephrosis
C1704321|ICD9CM|PT|581.3|Nephrotic syndrome with lesion of minimal change glomerulonephritis
C1704330|ICD9CM|AB|525.9|Dental disorder NOS
C1704330|ICD9CM|PT|525.9|Unspecified disorder of the teeth and supporting structures
C1706492|ICD9CM|PT|238.79|Other lymphatic and hematopoietic tissues
C1706492|ICD9CM|AB|238.79|Lymph/hematpoitc tis NEC
C1718233|ICD9CM|HT|707.2|Pressure ulcer stages
C1719272|ICD9CM|PT|00.44|Procedure on vessel bifurcation
C1719272|ICD9CM|AB|00.44|Proc-vessel bifurcation
C1719280|ICD9CM|PT|00.56|Insertion or replacement of implantable pressure sensor with lead for intracardiac or great vessel hemodynamic monitoring
C1719280|ICD9CM|AB|00.56|Ins/rep sens-crd/vsl mtr
C1719281|ICD9CM|PT|00.57|Implantation or replacement of subcutaneous device for intracardiac or great vessel hemodynamic monitoring
C1719281|ICD9CM|AB|00.57|Imp/rep subcue card dev
C1719284|ICD9CM|PT|00.85|Resurfacing hip, total, acetabulum and femoral head
C1719284|ICD9CM|AB|00.85|Resrf hip,total-acet/fem
C1719286|ICD9CM|PT|00.86|Resurfacing hip, partial, femoral head
C1719286|ICD9CM|AB|00.86|Resrf hip,part-fem head
C1719289|ICD9CM|PT|00.87|Resurfacing hip, partial, acetabulum
C1719289|ICD9CM|AB|00.87|Resrf hip,part-acetablum
C1719290|ICD9CM|HT|00.8|Other knee and hip procedures
C1719291|ICD9CM|PT|01.27|Removal of catheter(s) from cranial cavity or tissue
C1719291|ICD9CM|AB|01.27|Rem cath cranial cav/tis
C1719292|ICD9CM|PT|01.28|Placement of intracerebral catheter(s) via burr hole(s)
C1719292|ICD9CM|AB|01.28|Intracereb cth-burr hole
C1719295|ICD9CM|PT|052.2|Postvaricella myelitis
C1719295|ICD9CM|AB|052.2|Postvaricella myelitis
C1719297|ICD9CM|PT|053.14|Herpes zoster myelitis
C1719297|ICD9CM|AB|053.14|Herpes zoster myelitis
C1719298|ICD9CM|PT|054.74|Herpes simplex myelitis
C1719298|ICD9CM|AB|054.74|Herpes simplex myelitis
C1719299|ICD9CM|PT|13.90|Operation on lens, not elsewhere classified
C1719299|ICD9CM|AB|13.90|Operation on lens NEC
C1719300|ICD9CM|PT|13.91|Implantation of intraocular telescope prosthesis
C1719300|ICD9CM|AB|13.91|Impl intraoc telesc pros
C1719305|ICD9CM|PT|238.72|Low grade myelodysplastic syndrome lesions
C1719305|ICD9CM|AB|238.72|Low grde myelody syn les
C1719308|ICD9CM|PT|238.73|High grade myelodysplastic syndrome lesions
C1719308|ICD9CM|AB|238.73|Hi grde myelodys syn les
C1719319|ICD9CM|PT|284.01|Constitutional red blood cell aplasia
C1719319|ICD9CM|AB|284.01|Constitution RBC aplasia
C1719322|ICD9CM|PT|284.09|Other constitutional aplastic anemia
C1719322|ICD9CM|AB|284.09|Const aplastc anemia NEC
C1719323|ICD9CM|HT|284|Aplastic anemia and other bone marrow failure syndromes
C1719324|ICD9CM|PT|285.29|Anemia of other chronic disease
C1719324|ICD9CM|AB|285.29|Anemia-other chronic dis
C1719330|ICD9CM|PT|288.59|Other decreased white blood cell count
C1719330|ICD9CM|AB|288.59|Decreased WBC count NEC
C1719337|ICD9CM|PT|288.61|Lymphocytosis (symptomatic)
C1719337|ICD9CM|AB|288.61|Lymphocytosis-symptomatc
C1719340|ICD9CM|PT|288.63|Monocytosis (symptomatic)
C1719340|ICD9CM|AB|288.63|Monocytosis-symptomatic
C1719341|ICD9CM|PT|288.69|Other elevated white blood cell count
C1719341|ICD9CM|AB|288.69|Elevated WBC count NEC
C1719342|ICD9CM|PT|32.23|Open ablation of lung lesion or tissue
C1719342|ICD9CM|AB|32.23|Open abltn lung les/tiss
C1719343|ICD9CM|PT|32.24|Percutaneous ablation of lung lesion or tissue
C1719343|ICD9CM|AB|32.24|Perc abltn lung les/tiss
C1719344|ICD9CM|PT|32.25|Thoracoscopic ablation of lung lesion or tissue
C1719344|ICD9CM|AB|32.25|Thor abltn lung les/tiss
C1719345|ICD9CM|PT|32.26|Other and unspecified ablation of lung lesion or tissue
C1719345|ICD9CM|AB|32.26|Abltn lung tiss NEC/NOS
C1719346|ICD9CM|PT|323.01|Encephalitis and encephalomyelitis in viral diseases classified elsewhere
C1719346|ICD9CM|AB|323.01|Enceph/encephmye oth dis
C1719347|ICD9CM|PT|323.02|Myelitis in viral diseases classified elsewhere
C1719347|ICD9CM|AB|323.02|Myelitis-oth viral dis
C1719348|ICD9CM|PT|323.1|Encephalitis, myelitis, and encephalomyelitis in rickettsial diseases classified elsewhere
C1719348|ICD9CM|AB|323.1|Rickettsial encephalitis
C1719349|ICD9CM|PT|323.2|Encephalitis, myelitis, and encephalomyelitis in protozoal diseases classified elsewhere
C1719349|ICD9CM|AB|323.2|Protozoal encephalitis
C1719350|ICD9CM|PT|323.41|Other encephalitis and encephalomyelitis due to other infections classified elsewhere
C1719350|ICD9CM|AB|323.41|Ot encph/mye ot inf else
C1719351|ICD9CM|PT|323.42|Other myelitis due to other infections classified elsewhere
C1719351|ICD9CM|AB|323.42|Oth myelitis ot inf else
C1719352|ICD9CM|HT|323.4|Other encephalitis, myelitis, and encephalomyelitis due to other infections classified elsewhere
C1719353|ICD9CM|PT|323.51|Encephalitis and encephalomyelitis following immunization procedures
C1719353|ICD9CM|AB|323.51|Enceph/myel folwg immune
C1719358|ICD9CM|HT|323.5|Encephalitis, myelitis, and encephalomyelitis following immunization procedures
C1719360|ICD9CM|PT|323.62|Other postinfectious encephalitis and encephalomyelitis
C1719360|ICD9CM|AB|323.62|Postinf encephalitis NEC
C1719361|ICD9CM|HT|323.6|Postinfectious encephalitis, myelitis, and encephalomyelitis
C1719362|ICD9CM|PT|323.71|Toxic encephalitis and encephalomyelitis
C1719362|ICD9CM|AB|323.71|Toxic encph & encephlomy
C1719364|ICD9CM|HT|323.7|Toxic encephalitis, myelitis, and encephalomyelitis
C1719365|ICD9CM|PT|323.81|Other causes of encephalitis and encephalomyelitis
C1719365|ICD9CM|AB|323.81|Enceph & encephlalo NEC
C1719367|ICD9CM|PT|323.82|Other causes of myelitis
C1719367|ICD9CM|AB|323.82|Myelitis cause NEC
C1719368|ICD9CM|HT|323.8|Other causes of encephalitis, myelitis, and encephalomyelitis
C1719369|ICD9CM|PT|323.9|Unspecified causes of encephalitis, myelitis, and encephalomyelitis
C1719369|ICD9CM|AB|323.9|Encephalitis NOS
C1719370|ICD9CM|PT|33.71|Endoscopic insertion or replacement of bronchial valve(s), single lobe
C1719370|ICD9CM|AB|33.71|Endo ins/re bron val,one
C1719373|ICD9CM|PT|33.78|Endoscopic removal of bronchial device(s) or substances
C1719373|ICD9CM|AB|33.78|Endo rem bronch devc/sub
C1719374|ICD9CM|PT|33.79|Endoscopic insertion of other bronchial device or substances
C1719374|ICD9CM|AB|33.79|Endo insrt bronc def/sub
C1719378|ICD9CM|PT|331.83|Mild cognitive impairment, so stated
C1719378|ICD9CM|AB|331.83|Mild cognitive impairemt
C1719381|ICD9CM|PT|333.79|Other acquired torsion dystonia
C1719381|ICD9CM|AB|333.79|Acq torsion dystonia NEC
C1719382|ICD9CM|HT|333.7|Acquired torsion dystonia
C1719389|ICD9CM|PT|338.11|Acute pain due to trauma
C1719389|ICD9CM|AB|338.11|Acute pain due to trauma
C1719390|ICD9CM|PT|338.12|Acute post-thoracotomy pain
C1719390|ICD9CM|AB|338.12|Acute post-thoracot pain
C1719392|ICD9CM|PT|338.18|Other acute postoperative pain
C1719392|ICD9CM|AB|338.18|Acute postop pain NEC
C1719393|ICD9CM|PT|338.21|Chronic pain due to trauma
C1719393|ICD9CM|AB|338.21|Chronc pain d/t trauma
C1719394|ICD9CM|PT|338.28|Other chronic postoperative pain
C1719394|ICD9CM|AB|338.28|Chronic postop pain NEC
C1719395|ICD9CM|PT|338.3|Neoplasm related pain (acute) (chronic)
C1719395|ICD9CM|AB|338.3|Neoplasm related pain
C1719403|ICD9CM|PT|341.21|Acute (transverse) myelitis in conditions classified elsewhere
C1719403|ICD9CM|AB|341.21|Acute myelitis oth cond
C1719404|ICD9CM|PT|341.22|Idiopathic transverse myelitis
C1719404|ICD9CM|AB|341.22|Idiopathc trans myelitis
C1719405|ICD9CM|HT|345.4|Localization-related (focal) (partial) epilepsy and epileptic syndromes with complex partial seizures
C1719407|ICD9CM|HT|345.5|Localization-related (focal) (partial) epilepsy and epileptic syndromes with simple partial seizures
C1719409|ICD9CM|HT|345.8|Other forms of epilepsy and recurrent seizures
C1719410|ICD9CM|HT|345|Epilepsy and recurrent seizures
C1719411|ICD9CM|PT|35.55|Repair of ventricular septal defect with prosthesis, closed technique
C1719411|ICD9CM|AB|35.55|Pros rep ventrc def-clos
C1719412|ICD9CM|PT|36.33|Endoscopic transmyocardial revascularization
C1719412|ICD9CM|AB|36.33|Endo transmyo revascular
C1719415|ICD9CM|PT|36.34|Percutaneous transmyocardial revascularization
C1719415|ICD9CM|AB|36.34|Perc transmyo revascular
C1719417|ICD9CM|PT|37.20|Noninvasive programmed electrical stimulation [NIPS]
C1719417|ICD9CM|AB|37.20|Noninvas elect stimulatn
C1719445|ICD9CM|PT|379.60|Inflammation (infection) of postprocedural bleb, unspecified
C1719445|ICD9CM|AB|379.60|Inflam postproc bleb NOS
C1719446|ICD9CM|PT|379.61|Inflammation (infection) of postprocedural bleb, stage 1
C1719446|ICD9CM|AB|379.61|Inflam postproc bleb, 1
C1719447|ICD9CM|PT|379.62|Inflammation (infection) of postprocedural bleb, stage 2
C1719447|ICD9CM|AB|379.62|Inflam postproc bleb, 2
C1719448|ICD9CM|PT|379.63|Inflammation (infection) of postprocedural bleb, stage 3
C1719448|ICD9CM|AB|379.63|Inflam postproc bleb, 3
C1719449|ICD9CM|HT|379.6|Inflammation (infection) of postprocedural bleb
C1719452|ICD9CM|PT|389.11|Sensory hearing loss, bilateral
C1719452|ICD9CM|AB|389.11|Sensry hearng loss,bilat
C1719455|ICD9CM|PT|389.16|Sensorineural hearing loss, asymmetrical
C1719455|ICD9CM|AB|389.16|Sensoneur hear loss asym
C1719460|ICD9CM|PT|403.00|Hypertensive chronic kidney disease, malignant, with chronic kidney disease stage I through stage IV, or unspecified
C1719460|ICD9CM|AB|403.00|Mal hy kid w cr kid I-IV
C1719461|ICD9CM|PT|403.01|Hypertensive chronic kidney disease, malignant, with chronic kidney disease stage V or end stage renal disease
C1719461|ICD9CM|AB|403.01|Mal hyp kid w cr kid V
C1719462|ICD9CM|HT|403.0|Hypertensive chronic kidney disease, malignant
C1719464|ICD9CM|PT|404.00|Hypertensive heart and chronic kidney disease, malignant, without heart failure and with chronic kidney disease stage I through stage IV, or unspecified
C1719464|ICD9CM|AB|404.00|Mal hy ht/kd I-IV w/o hf
C1719465|ICD9CM|PT|404.01|Hypertensive heart and chronic kidney disease, malignant, with heart failure and with chronic kidney disease stage I through stage IV, or unspecified
C1719465|ICD9CM|AB|404.01|Mal hyp ht/kd I-IV w hf
C1719466|ICD9CM|PT|404.02|Hypertensive heart and chronic kidney disease, malignant, without heart failure and with chronic kidney disease stage V or end stage renal disease
C1719466|ICD9CM|AB|404.02|Mal hy ht/kd st V w/o hf
C1719467|ICD9CM|PT|404.03|Hypertensive heart and chronic kidney disease, malignant, with heart failure and with chronic kidney disease stage V or end stage renal disease
C1719467|ICD9CM|AB|404.03|Mal hyp ht/kd stg V w hf
C1719468|ICD9CM|HT|404.0|Hypertensive heart and chronic kidney disease, malignant
C1719469|ICD9CM|HT|404|Hypertensive heart and chronic kidney disease
C1719478|ICD9CM|PT|50.23|Open ablation of liver lesion or tissue
C1719478|ICD9CM|AB|50.23|Opn abltn liver les/tiss
C1719479|ICD9CM|PT|50.24|Percutaneous ablation of liver lesion or tissue
C1719479|ICD9CM|AB|50.24|Perc abltn liver les/tis
C1719480|ICD9CM|PT|50.25|Laparoscopic ablation of liver lesion or tissue
C1719480|ICD9CM|AB|50.25|Lap abltn liver les/tiss
C1719481|ICD9CM|PT|50.26|Other and unspecified ablation of liver lesion or tissue
C1719481|ICD9CM|AB|50.26|Abltn liver les/tiss NEC
C1719483|ICD9CM|PT|519.19|Other diseases of trachea and bronchus
C1719483|ICD9CM|AB|519.19|Trachea & bronch dis NEC
C1719490|ICD9CM|PT|523.00|Acute gingivitis, plaque induced
C1719490|ICD9CM|AB|523.00|Acute gingititis, plaque
C1719491|ICD9CM|PT|523.01|Acute gingivitis, non-plaque induced
C1719491|ICD9CM|AB|523.01|Ac gingivitis,nonplaque
C1719492|ICD9CM|PT|523.11|Chronic gingivitis, non-plaque induced
C1719492|ICD9CM|AB|523.11|Chr gingivitis-nonplaque
C1719493|ICD9CM|PT|523.30|Aggressive periodontitis, unspecified
C1719493|ICD9CM|AB|523.30|Aggres periodontitis NOS
C1719494|ICD9CM|PT|523.31|Aggressive periodontitis, localized
C1719494|ICD9CM|AB|523.31|Aggres periodontitis,loc
C1719495|ICD9CM|PT|523.32|Aggressive periodontitis, generalized
C1719495|ICD9CM|AB|523.32|Aggres periodontitis,gen
C1719497|ICD9CM|PT|523.41|Chronic periodontitis, localized
C1719497|ICD9CM|AB|523.41|Chr periodontitis, local
C1719498|ICD9CM|PT|523.42|Chronic periodontitis, generalized
C1719498|ICD9CM|AB|523.42|Chron periodontitis,gen
C1719507|ICD9CM|PT|525.60|Unspecified unsatisfactory restoration of tooth
C1719507|ICD9CM|AB|525.60|Unsat restore tooth NOS
C1719512|ICD9CM|PT|525.63|Fractured dental restorative material without loss of material
C1719512|ICD9CM|AB|525.63|Fx dental mat w/o loss
C1719513|ICD9CM|PT|525.64|Fractured dental restorative material with loss of material
C1719513|ICD9CM|AB|525.64|Fx dentl material w loss
C1719514|ICD9CM|PT|525.65|Contour of existing restoration of tooth biologically incompatible with oral health
C1719514|ICD9CM|AB|525.65|Contour restore tooth
C1719517|ICD9CM|PT|525.67|Poor aesthetics of existing restoration
C1719517|ICD9CM|AB|525.67|Poor aesthetics restore
C1719518|ICD9CM|PT|525.69|Other unsatisfactory restoration of existing tooth
C1719518|ICD9CM|AB|525.69|Unsat restore tooth NEC
C1719519|ICD9CM|HT|525.6|Unsatisfactory restoration of tooth
C1719521|ICD9CM|PT|526.61|Perforation of root canal space
C1719521|ICD9CM|AB|526.61|Perfor root canal space
C1719522|ICD9CM|PT|526.62|Endodontic overfill
C1719522|ICD9CM|AB|526.62|Endodontic overfill
C1719523|ICD9CM|PT|526.63|Endodontic underfill
C1719523|ICD9CM|AB|526.63|Endodontic underfill
C1719524|ICD9CM|HT|526.6|Periradicular pathology associated with previous endodontic treatment
C1719526|ICD9CM|PT|528.01|Mucositis (ulcerative) due to antineoplastic therapy
C1719526|ICD9CM|AB|528.01|Mucosits d/t antineo rx
C1719527|ICD9CM|PT|528.02|Mucositis (ulcerative) due to other drugs
C1719527|ICD9CM|AB|528.02|Mucositis d/t drugs NEC
C1719528|ICD9CM|PT|528.09|Other stomatitis and mucositis (ulcerative)
C1719528|ICD9CM|HT|528.0|Stomatitis and mucositis (ulcerative)
C1719528|ICD9CM|AB|528.09|Stomatits & mucosits NEC
C1719533|ICD9CM|PT|55.32|Open ablation of renal lesion or tissue
C1719533|ICD9CM|AB|55.32|Opn abltn renal les/tiss
C1719534|ICD9CM|PT|55.33|Percutaneous ablation of renal lesion or tissue
C1719534|ICD9CM|AB|55.33|Perc abltn renl les/tiss
C1719535|ICD9CM|PT|55.34|Laparoscopic ablation of renal lesion or tissue
C1719535|ICD9CM|AB|55.34|Lap abltn renal les/tiss
C1719536|ICD9CM|PT|55.35|Other and unspecified ablation of renal lesion or tissue
C1719536|ICD9CM|AB|55.35|Abltn renal les/tiss NEC
C1719538|ICD9CM|PT|600.00|Hypertrophy (benign) of prostate without urinary obstruction and other lower urinary tract symptom (LUTS)
C1719538|ICD9CM|AB|600.00|BPH w/o urinary obs/LUTS
C1719539|ICD9CM|PT|600.20|Benign localized hyperplasia of prostate without urinary obstruction and other lower urinary tract symptoms (LUTS)
C1719539|ICD9CM|AB|600.20|BPH loc w/o ur obs/LUTS
C1719540|ICD9CM|PT|600.90|Hyperplasia of prostate, unspecified, without urinary obstruction and other lower urinary symptoms (LUTS)
C1719540|ICD9CM|AB|600.90|BPH NOS w/o ur obs/LUTS
C1719541|ICD9CM|PT|608.21|Extravaginal torsion of spermatic cord
C1719541|ICD9CM|AB|608.21|Extravag tors sperm cord
C1719542|ICD9CM|PT|608.22|Intravaginal torsion of spermatic cord
C1719542|ICD9CM|AB|608.22|Intravag tors sperm cord
C1719543|ICD9CM|PT|616.81|Mucositis (ulcerative) of cervix, vagina, and vulva
C1719543|ICD9CM|AB|616.81|Mucositis cerv,vag,vulva
C1719544|ICD9CM|PT|616.89|Other inflammatory disease of cervix, vagina and vulva
C1719544|ICD9CM|AB|616.89|Inflm cerv,vag,vulva NEC
C1719546|ICD9CM|PT|618.84|Cervical stump prolapse
C1719546|ICD9CM|AB|618.84|Cervical stump prolapse
C1719551|ICD9CM|PT|629.29|Other female genital mutilation status
C1719551|ICD9CM|AB|629.29|Fem genital mutilate NEC
C1719558|ICD9CM|PT|649.00|Tobacco use disorder complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C1719558|ICD9CM|AB|649.00|Tobacco use disord-unsp
C1719559|ICD9CM|PT|649.01|Tobacco use disorder complicating pregnancy, childbirth, or the puerperium, delivered, with or without mention of antepartum condition
C1719559|ICD9CM|AB|649.01|Tobacco use disor-delliv
C1719560|ICD9CM|PT|649.02|Tobacco use disorder complicating pregnancy, childbirth, or the puerperium, delivered, with mention of postpartum complication
C1719560|ICD9CM|AB|649.02|Tobacco use dis-del-p/p
C1719561|ICD9CM|PT|649.03|Tobacco use disorder complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C1719561|ICD9CM|AB|649.03|Tobacco use dis-antepart
C1719562|ICD9CM|PT|649.04|Tobacco use disorder complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication
C1719562|ICD9CM|AB|649.04|Tobacco use dis-postpart
C1719563|ICD9CM|HT|649.0|Tobacco use disorder complicating pregnancy, childbirth, or the puerperium
C1719565|ICD9CM|PT|649.10|Obesity complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C1719565|ICD9CM|AB|649.10|Obesity-unspecified
C1719566|ICD9CM|PT|649.11|Obesity complicating pregnancy, childbirth, or the puerperium, delivered, with or without mention of antepartum condition
C1719566|ICD9CM|AB|649.11|Obesity-delivered
C1719567|ICD9CM|PT|649.12|Obesity complicating pregnancy, childbirth, or the puerperium, delivered, with mention of postpartum complication
C1719567|ICD9CM|AB|649.12|Obesity-delivered w p/p
C1719568|ICD9CM|PT|649.13|Obesity complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C1719568|ICD9CM|AB|649.13|Obesity-antepartum
C1719569|ICD9CM|PT|649.14|Obesity complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication
C1719569|ICD9CM|AB|649.14|Obesity-postpartum
C1719570|ICD9CM|HT|649.1|Obesity complicating pregnancy, childbirth, or the puerperium
C1719571|ICD9CM|PT|649.20|Bariatric surgery status complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C1719571|ICD9CM|AB|649.20|Bariatric surg stat-unsp
C1719572|ICD9CM|PT|649.21|Bariatric surgery status complicating pregnancy, childbirth, or the puerperium, delivered, with or without mention of antepartum condition
C1719572|ICD9CM|AB|649.21|Bariatric surg stat-del
C1719573|ICD9CM|PT|649.22|Bariatric surgery status complicating pregnancy, childbirth, or the puerperium, delivered, with mention of postpartum complication
C1719573|ICD9CM|AB|649.22|Bariatric surg-del w p/p
C1719574|ICD9CM|PT|649.23|Bariatric surgery status complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C1719574|ICD9CM|AB|649.23|Bariatrc surg stat-antep
C1719575|ICD9CM|PT|649.24|Bariatric surgery status complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication
C1719575|ICD9CM|AB|649.24|Bariatrc surg stat w p/p
C1719576|ICD9CM|HT|649.2|Bariatric surgery status complicating pregnancy, childbirth, or the puerperium
C1719580|ICD9CM|PT|649.30|Coagulation defects complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C1719580|ICD9CM|AB|649.30|Coagulation def-unspec
C1719581|ICD9CM|PT|649.31|Coagulation defects complicating pregnancy, childbirth, or the puerperium, delivered, with or without mention of antepartum condition
C1719581|ICD9CM|AB|649.31|Coagulation def-deliv
C1719582|ICD9CM|PT|649.32|Coagulation defects complicating pregnancy, childbirth, or the puerperium, delivered, with mention of postpartum complication
C1719582|ICD9CM|AB|649.32|Coagulatn def-del w p/p
C1719583|ICD9CM|PT|649.33|Coagulation defects complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C1719583|ICD9CM|AB|649.33|Coagulation def-antepart
C1719584|ICD9CM|PT|649.34|Coagulation defects complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication
C1719584|ICD9CM|AB|649.34|Coagulation def-postpart
C1719585|ICD9CM|HT|649.3|Coagulation defects complicating pregnancy, childbirth, or the puerperium
C1719586|ICD9CM|PT|649.40|Epilepsy complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C1719586|ICD9CM|AB|649.40|Epilepsy-unspecified
C1719587|ICD9CM|PT|649.41|Epilepsy complicating pregnancy, childbirth, or the puerperium, delivered, with or without mention of antepartum condition
C1719587|ICD9CM|AB|649.41|Epilepsy-delivered
C1719588|ICD9CM|PT|649.42|Epilepsy complicating pregnancy, childbirth, or the puerperium, delivered, with mention of postpartum complication
C1719588|ICD9CM|AB|649.42|Epilepsy-delivered w p/p
C1719589|ICD9CM|PT|649.43|Epilepsy complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C1719589|ICD9CM|AB|649.43|Epilepsy-antepartum
C1719590|ICD9CM|PT|649.44|Epilepsy complicating pregnancy, childbirth, or the puerperium, postpartum condition or complication
C1719590|ICD9CM|AB|649.44|Epilepsy-postpartum
C1719591|ICD9CM|HT|649.4|Epilepsy complicating pregnancy, childbirth, or the puerperium
C1719592|ICD9CM|PT|649.50|Spotting complicating pregnancy, unspecified as to episode of care or not applicable
C1719592|ICD9CM|AB|649.50|Spotting-unspecified
C1719593|ICD9CM|PT|649.51|Spotting complicating pregnancy, delivered, with or without mention of antepartum condition
C1719593|ICD9CM|AB|649.51|Spotting-delivered
C1719594|ICD9CM|PT|649.53|Spotting complicating pregnancy, antepartum condition or complication
C1719594|ICD9CM|AB|649.53|Spotting-antepartum
C1719595|ICD9CM|HT|649.5|Spotting complicating pregnancy
C1719596|ICD9CM|PT|649.60|Uterine size date discrepancy, unspecified as to episode of care or not applicable
C1719596|ICD9CM|AB|649.60|Uterine size descrp-unsp
C1719597|ICD9CM|PT|649.61|Uterine size date discrepancy, delivered, with or without mention of antepartum condition
C1719597|ICD9CM|AB|649.61|Uterine size descrep-del
C1719598|ICD9CM|PT|649.62|Uterine size date discrepancy, delivered, with mention of postpartum complication
C1719598|ICD9CM|AB|649.62|Uterine size-del w p/p
C1719599|ICD9CM|PT|649.63|Uterine size date discrepancy, antepartum condition or complication
C1719599|ICD9CM|AB|649.63|Uterine size des-antepar
C1719600|ICD9CM|PT|649.64|Uterine size date discrepancy, postpartum condition or complication
C1719600|ICD9CM|AB|649.64|Uterine size descrep-p/p
C1719601|ICD9CM|HT|649.6|Uterine size date discrepancy
C1719602|ICD9CM|HT|649|Other conditions or status of the mother complicating pregnancy, childbirth, or the puerperium
C1719605|ICD9CM|PT|68.39|Other and unspecified subtotal abdominal hysterectomy
C1719605|ICD9CM|AB|68.39|Subtotl abd hyst NEC/NOS
C1719606|ICD9CM|PT|68.41|Laparoscopic total abdominal hysterectomy
C1719606|ICD9CM|AB|68.41|Lap total abdominal hyst
C1719609|ICD9CM|PT|68.59|Other and unspecified vaginal hysterectomy
C1719609|ICD9CM|AB|68.59|Vag hysterectomy NEC/NOS
C1719610|ICD9CM|PT|68.61|Laparoscopic radical abdominal hysterectomy
C1719610|ICD9CM|AB|68.61|Lap radical abdomnl hyst
C1719613|ICD9CM|PT|68.69|Other and unspecified radical abdominal hysterectomy
C1719613|ICD9CM|AB|68.69|Radical abd hyst NEC/NOS
C1719615|ICD9CM|PT|68.79|Other and unspecified radical vaginal hysterectomy
C1719615|ICD9CM|AB|68.79|Radical vag hyst NEC/NOS
C1719618|ICD9CM|PT|729.71|Nontraumatic compartment syndrome of upper extremity
C1719618|ICD9CM|AB|729.71|Nontraum comp syn-up ext
C1719620|ICD9CM|PT|729.72|Nontraumatic compartment syndrome of lower extremity
C1719620|ICD9CM|AB|729.72|Nontraum comp syn-low ex
C1719621|ICD9CM|PT|729.73|Nontraumatic compartment syndrome of abdomen
C1719621|ICD9CM|AB|729.73|Nontrauma comp syn-abd
C1719622|ICD9CM|PT|729.79|Nontraumatic compartment syndrome of other sites
C1719622|ICD9CM|AB|729.79|Nontrauma comp syn NEC
C1719623|ICD9CM|HT|729.7|Nontraumatic compartment syndrome
C1719624|ICD9CM|AB|731.3|Major osseous defects
C1719624|ICD9CM|PT|731.3|Major osseous defects
C1719625|ICD9CM|PT|768.3|Fetal distress first noted during labor and delivery, in liveborn infant
C1719625|ICD9CM|AB|768.3|Fetal distrs dur lab/del
C1719629|ICD9CM|PT|775.81|Other acidosis of newborn
C1719629|ICD9CM|AB|775.81|NB acidosis NEC
C1719633|ICD9CM|HT|775.8|Other neonatal endocrine and metabolic disturbances
C1719633|ICD9CM|PT|775.89|Other neonatal endocrine and metabolic disturbances
C1719633|ICD9CM|AB|775.89|Neonat endo/met dis NEC
C1719639|ICD9CM|PT|780.95|Excessive crying of child, adolescent, or adult
C1719639|ICD9CM|AB|780.95|Excs cry chld,adol,adult
C1719644|ICD9CM|PT|793.91|Image test inconclusive due to excess body fat
C1719644|ICD9CM|AB|793.91|Image test incon d/t fat
C1719645|ICD9CM|PT|793.99|Other nonspecific (abnormal) findings on radiological and other examinations of body structure
C1719645|ICD9CM|AB|793.99|Nonsp abn find-body NEC
C1719648|ICD9CM|PT|795.06|Papanicolaou smear of cervix with cytologic evidence of malignancy
C1719648|ICD9CM|AB|795.06|Pap smr cytol evid malig
C1719649|ICD9CM|PT|795.81|Elevated carcinoembryonic antigen [CEA]
C1719649|ICD9CM|AB|795.81|Elev ca-embryoic antigen
C1719650|ICD9CM|PT|795.89|Other abnormal tumor markers
C1719650|ICD9CM|AB|795.89|Abnorml tumor marker NEC
C1719651|ICD9CM|HT|795.8|Abnormal tumor markers
C1719657|ICD9CM|PT|958.91|Traumatic compartment syndrome of upper extremity
C1719657|ICD9CM|AB|958.91|Trauma comp synd up ext
C1719659|ICD9CM|PT|958.92|Traumatic compartment syndrome of lower extremity
C1719659|ICD9CM|AB|958.92|Trauma comp synd low ext
C1719660|ICD9CM|PT|958.93|Traumatic compartment syndrome of abdomen
C1719660|ICD9CM|AB|958.93|Trauma compart synd abd
C1719661|ICD9CM|PT|958.99|Traumatic compartment syndrome of other sites
C1719661|ICD9CM|AB|958.99|Trauma compart synd NEC
C1719662|ICD9CM|HT|958.9|Traumatic compartment syndrome
C1719666|ICD9CM|PT|995.20|Unspecified adverse effect of unspecified drug, medicinal and biological substance
C1719666|ICD9CM|AB|995.20|Adv eff med/biol sub NOS
C1719667|ICD9CM|PT|995.22|Unspecified adverse effect of anesthesia
C1719667|ICD9CM|AB|995.22|Adv eff anesthesia NOS
C1719668|ICD9CM|PT|995.23|Unspecified adverse effect of insulin
C1719668|ICD9CM|AB|995.23|Adverse eff insulin NOS
C1719669|ICD9CM|PT|995.27|Other drug allergy
C1719669|ICD9CM|AB|995.27|Drug allergy NEC
C1719670|ICD9CM|PT|995.29|Unspecified adverse effect of other drug, medicinal and biological substance
C1719670|ICD9CM|AB|995.29|Adv eff med/biol NEC/NOS
C1719672|ICD9CM|PT|995.92|Severe sepsis
C1719672|ICD9CM|AB|995.92|Severe sepsis
C1719676|ICD9CM|PT|995.93|Systemic inflammatory response syndrome due to noninfectious process without acute organ dysfunction
C1719676|ICD9CM|AB|995.93|SIRS-noninf w/o ac or ds
C1719677|ICD9CM|PT|995.94|Systemic inflammatory response syndrome due to noninfectious process with acute organ dysfunction
C1719677|ICD9CM|AB|995.94|SIRS-noninf w ac org dys
C1719681|ICD9CM|PT|V26.31|Testing of female for genetic disease carrier status
C1719681|ICD9CM|AB|V26.31|Fem genetic test dis car
C1719682|ICD9CM|PT|V26.32|Other genetic testing of female
C1719682|ICD9CM|AB|V26.32|Female genetic test NEC
C1719683|ICD9CM|PT|V26.34|Testing of male for genetic disease carrier status
C1719683|ICD9CM|AB|V26.34|Male genetc test dis car
C1719684|ICD9CM|PT|V26.39|Other genetic testing of male
C1719684|ICD9CM|AB|V26.39|Male genetic test NEC
C1719685|ICD9CM|HT|V28|Encounter for antenatal screening of mother
C1719686|ICD9CM|PT|V45.86|Bariatric surgery status
C1719686|ICD9CM|AB|V45.86|Bariatric surgery status
C1719690|ICD9CM|PT|V58.30|Encounter for change or removal of nonsurgical wound dressing
C1719690|ICD9CM|AB|V58.30|Attn rem nonsurg dressng
C1719692|ICD9CM|PT|V58.31|Encounter for change or removal of surgical wound dressing
C1719692|ICD9CM|AB|V58.31|Attn rem surg dressing
C1719693|ICD9CM|PT|V58.32|Encounter for removal of sutures
C1719693|ICD9CM|AB|V58.32|Attn removal of sutures
C1719694|ICD9CM|HT|V58.3|Attention to dressings and sutures
C1719697|ICD9CM|HT|V70-V82.99|PERSONS WITHOUT REPORTED DIAGNOSIS ENCOUNTERED DURING EXAMINATION AND INVESTIGATION OF INDIVIDUALS AND POPULATIONS
C1719698|ICD9CM|PT|V72.11|Encounter for hearing examination following failed hearing screening
C1719698|ICD9CM|AB|V72.11|Hearing exam-fail screen
C1719699|ICD9CM|PT|V72.19|Other examination of ears and hearing
C1719699|ICD9CM|AB|V72.19|Exam ears & hearing NEC
C1719700|ICD9CM|PT|V82.71|Screening for genetic disease carrier status
C1719700|ICD9CM|AB|V82.71|Screen-gentc dis carrier
C1719706|ICD9CM|PT|V86.0|Estrogen receptor positive status [ER+]
C1719706|ICD9CM|AB|V86.0|Estrogen recep pstv stat
C1719707|ICD9CM|PT|V86.1|Estrogen receptor negative status [ER-]
C1719707|ICD9CM|AB|V86.1|Estrogen recep neg stat
C1719710|ICD9CM|PT|338.22|Chronic post-thoracotomy pain
C1719710|ICD9CM|AB|338.22|Chron post-thoracot pain
C1719711|ICD9CM|PT|68.49|Other and unspecified total abdominal hysterectomy
C1719711|ICD9CM|AB|68.49|Total abd hyst NEC/NOS
C1719713|ICD9CM|PT|526.69|Other periradicular pathology associated with previous endodontic treatment
C1719713|ICD9CM|AB|526.69|Periradicular path NEC
C1719714|ICD9CM|PT|528.00|Stomatitis and mucositis, unspecified
C1719714|ICD9CM|AB|528.00|Stomatitis/mucositis NOS
C1719715|ICD9CM|PT|01.26|Insertion of catheter(s) into cranial cavity or tissue
C1719715|ICD9CM|AB|01.26|Ins cath cranial cav/tis
C1719716|ICD9CM|PT|39.74|Endovascular removal of obstruction from head and neck vessel(s)
C1719716|ICD9CM|AB|39.74|Endo rem obs hd/neck ves
C1719717|ICD9CM|PT|523.10|Chronic gingivitis, plaque induced
C1719717|ICD9CM|AB|523.10|Chronc gingititis,plaque
C1719719|ICD9CM|PT|525.66|Allergy to existing dental restorative material
C1719719|ICD9CM|AB|525.66|Allergy dental res mat
C1719722|ICD9CM|PT|323.61|Infectious acute disseminated encephalomyelitis (ADEM)
C1719722|ICD9CM|AB|323.61|Inf ac dis encephalomyel
C1719723|ICD9CM|PT|338.19|Other acute pain
C1719723|ICD9CM|AB|338.19|Acute pain NEC
C1719729|ICD9CM|PT|68.71|Laparoscopic radical vaginal hysterectomy [LRVH]
C1719729|ICD9CM|AB|68.71|Lap radical vaginal hyst
C1719811|ICD9CM|PT|707.23|Pressure ulcer, stage III
C1719811|ICD9CM|AB|707.23|Pressure ulcer,stage III
C1719910|ICD9CM|AB|707.24|Pressure ulcer, stage IV
C1719910|ICD9CM|PT|707.24|Pressure ulcer, stage IV
C1720363|ICD9CM|PT|707.25|Pressure ulcer, unstageable
C1720363|ICD9CM|AB|707.25|Pressure ulcer,unstagebl
C1720518|ICD9CM|AB|707.22|Pressure ulcer, stage II
C1720518|ICD9CM|PT|707.22|Pressure ulcer, stage II
C1720599|ICD9CM|AB|707.21|Pressure ulcer, stage I
C1720599|ICD9CM|PT|707.21|Pressure ulcer, stage I
C1720771|ICD9CM|HT|603|Hydrocele
C1720771|ICD9CM|AB|603.9|Hydrocele NOS
C1720771|ICD9CM|PT|603.9|Hydrocele, unspecified
C1735601|ICD9CM|PT|364.81|Floppy iris syndrome
C1735601|ICD9CM|AB|364.81|Floppy iris syndrome
C1739094|ICD9CM|PT|005.1|Botulism food poisoning
C1739094|ICD9CM|AB|005.1|Botulism food poisoning
C1739123|ICD9CM|PT|780.66|Febrile nonhemolytic transfusion reaction
C1739123|ICD9CM|AB|780.66|Feb nonhemo transf react
C1739395|ICD9CM|PT|429.83|Takotsubo syndrome
C1739395|ICD9CM|AB|429.83|Takotsubo syndrome
C1744615|ICD9CM|HT|884|Multiple and unspecified open wound of upper limb
C1744616|ICD9CM|HT|891|Open wound of knee, leg [except thigh], and ankle
C1744618|ICD9CM|PT|71.11|Biopsy of vulva
C1744618|ICD9CM|AB|71.11|Vulvar biopsy
C1744632|ICD9CM|HT|895|Traumatic amputation of toe(s) (complete) (partial)
C1761613|ICD9CM|AB|372.71|Hyperemia of conjunctiva
C1761613|ICD9CM|PT|372.71|Hyperemia of conjunctiva
C1800706|ICD9CM|PT|516.31|Idiopathic pulmonary fibrosis
C1800706|ICD9CM|AB|516.31|Idiopath pulmon fibrosis
C1812606|ICD9CM|HT|949|Burn, unspecified site
C1812609|ICD9CM|AB|050.0|Variola major
C1812609|ICD9CM|PT|050.0|Variola major
C1812610|ICD9CM|HT|010.9|Primary tuberculous infection, unspecified type
C1812611|ICD9CM|PT|010.90|Primary tuberculous infection, unspecified, unspecified
C1812611|ICD9CM|AB|010.90|Primary TB NOS-unspec
C1812612|ICD9CM|PT|010.00|Primary tuberculous infection, unspecified
C1812612|ICD9CM|AB|010.00|Prim TB complex-unspec
C1812613|ICD9CM|PT|894.0|Multiple and unspecified open wound of lower limb, without mention of complication
C1812613|ICD9CM|AB|894.0|Open wound of leg NEC
C1812614|ICD9CM|HT|942.0|Burn of trunk, unspecified degree
C1812615|ICD9CM|PT|942.00|Burn of unspecified degree of trunk, unspecified site
C1812615|ICD9CM|AB|942.00|Burn NOS trunk-unspec
C1812616|ICD9CM|PT|946.0|Burns of multiple specified sites, unspecified degree
C1812616|ICD9CM|AB|946.0|Burn NOS multiple site
C1812617|ICD9CM|PT|945.00|Burn of unspecified degree of lower limb [leg], unspecified site
C1812617|ICD9CM|AB|945.00|Burn NOS leg-unspec
C1812618|ICD9CM|HT|945.0|Burn of lower limb(s), unspecified degree
C1812619|ICD9CM|HT|944.0|Burn of wrist(s) and hand(s), unspecified degree
C1812620|ICD9CM|PT|657.00|Polyhydramnios, unspecified as to episode of care or not applicable
C1812620|ICD9CM|AB|657.00|Polyhydramnios-unspec
C1812621|ICD9CM|PT|672.00|Pyrexia of unknown origin during the puerperium, unspecified as to episode of care or not applicable
C1812621|ICD9CM|AB|672.00|Puerperal pyrexia-unspec
C1812623|ICD9CM|HT|373|Inflammation of eyelids
C1812624|ICD9CM|AB|305.01|Alcohol abuse-continuous
C1812624|ICD9CM|PT|305.01|Alcohol abuse, continuous
C1812625|ICD9CM|PT|665.03|Rupture of uterus before onset of labor, antepartum condition or complication
C1812625|ICD9CM|AB|665.03|Prelab rupt uter-antepar
C1812626|ICD9CM|PT|664.01|First-degree perineal laceration, delivered, with or without mention of antepartum condition
C1812626|ICD9CM|AB|664.01|Del w 1 deg lacerat-del
C1812627|ICD9CM|PT|674.04|Cerebrovascular disorders in the puerperium, postpartum condition or complication
C1812627|ICD9CM|AB|674.04|Cerebrovasc dis-postpart
C1827466|ICD9CM|PT|377.02|Papilledema associated with decreased ocular pressure
C1827466|ICD9CM|AB|377.02|Papilledema w decr press
C1830412|ICD9CM|AB|E013.1|Laundry
C1830412|ICD9CM|PT|E013.1|Activities involving laundry
C1841680|ICD9CM|PT|752.47|Longitudinal vaginal septum
C1841680|ICD9CM|AB|752.47|Longitud vaginal septum
C1856006|ICD9CM|PT|752.46|Transverse vaginal septum
C1856006|ICD9CM|AB|752.46|Transv vaginal septum
C1861783|ICD9CM|PT|447.4|Celiac artery compression syndrome
C1861783|ICD9CM|AB|447.4|Celiac art compress syn
C1868193|ICD9CM|PT|512.81|Primary spontaneous pneumothorax
C1868193|ICD9CM|AB|512.81|Prim spont pneumothorax
C1879322|ICD9CM|PT|28.0|Incision and drainage of tonsil and peritonsillar structures
C1879322|ICD9CM|AB|28.0|Peritonsillar i & d
C1879328|ICD9CM|PT|369.00|Profound impairment, both eyes, impairment level not further specified
C1879328|ICD9CM|AB|369.00|Both eyes blind-who def
C1955490|ICD9CM|PT|664.60|Anal sphincter tear complicating delivery, not associated with third-degree perineal laceration, unspecified as to episode of care or not applicable
C1955490|ICD9CM|AB|664.60|Anal sphincter tear NOS
C1955491|ICD9CM|PT|664.61|Anal sphincter tear complicating delivery, not associated with third-degree perineal laceration, delivered, with or without mention of antepartum condition
C1955491|ICD9CM|AB|664.61|Anal sphincter tear-del
C1955492|ICD9CM|PT|664.64|Anal sphincter tear complicating delivery, not associated with third-degree perineal laceration, postpartum condition or complication
C1955492|ICD9CM|AB|664.64|Anal sphinctr tear w p/p
C1955493|ICD9CM|HT|664.6|Anal sphincter tear complicating delivery, not associated with third-degree perineal laceration
C1955495|ICD9CM|PT|70.53|Repair of cystocele and rectocele with graft or prosthesis
C1955495|ICD9CM|AB|70.53|Cysto & recto w grf/pros
C1955496|ICD9CM|PT|70.54|Repair of cystocele with graft or prosthesis
C1955496|ICD9CM|AB|70.54|Rep cystocel w grft/pros
C1955498|ICD9CM|PT|70.55|Repair of rectocele with graft or prosthesis
C1955498|ICD9CM|AB|70.55|Rep rectocele w grf/pros
C1955499|ICD9CM|PT|70.63|Vaginal construction with graft or prosthesis
C1955499|ICD9CM|AB|70.63|Vaginal const w grf/pros
C1955500|ICD9CM|PT|70.64|Vaginal reconstruction with graft or prosthesis
C1955500|ICD9CM|AB|70.64|Vag reconst w grft/pros
C1955501|ICD9CM|PT|70.78|Vaginal suspension and fixation with graft or prosthesis
C1955501|ICD9CM|AB|70.78|Vag susp/fix w grft/pros
C1955502|ICD9CM|PT|70.93|Other operations on cul-de-sac with graft or prosthesis
C1955502|ICD9CM|AB|70.93|Cul-de-sac grf/pros NEC
C1955504|ICD9CM|PT|70.94|Insertion of biological graft
C1955504|ICD9CM|AB|70.94|Insert biological graft
C1955511|ICD9CM|PT|70.95|Insertion of synthetic graft or prosthesis
C1955511|ICD9CM|AB|70.95|Insert synth graft/prost
C1955516|ICD9CM|AB|787.23|Dysphagia, pharyngeal
C1955516|ICD9CM|PT|787.23|Dysphagia, pharyngeal phase
C1955517|ICD9CM|PT|787.24|Dysphagia, pharyngoesophageal phase
C1955517|ICD9CM|AB|787.24|Dysphagia,pharyngoesoph
C1955518|ICD9CM|PT|787.29|Other dysphagia
C1955518|ICD9CM|AB|787.29|Dysphagia NEC
C1955521|ICD9CM|PT|789.59|Other ascites
C1955521|ICD9CM|AB|789.59|Ascites NEC
C1955522|ICD9CM|PT|84.80|Insertion or replacement of interspinous process device(s)
C1955522|ICD9CM|AB|84.80|Ins/repl interspine dev
C1955525|ICD9CM|PT|84.81|Revision of interspinous process device(s)
C1955525|ICD9CM|AB|84.81|Rev interspine device
C1955527|ICD9CM|PT|84.82|Insertion or replacement of pedicle-based dynamic stabilization device(s)
C1955527|ICD9CM|AB|84.82|Ins/repl pdcl stabil dev
C1955528|ICD9CM|PT|84.83|Revision of pedicle-based dynamic stabilization device(s)
C1955528|ICD9CM|AB|84.83|Rev pedcl dyn stabil dev
C1955530|ICD9CM|PT|84.84|Insertion or replacement of facet replacement device(s)
C1955530|ICD9CM|AB|84.84|Ins/repl facet replc dev
C1955532|ICD9CM|PT|84.85|Revision of facet replacement device(s)
C1955532|ICD9CM|AB|84.85|Rev facet replace device
C1955534|ICD9CM|HT|84.8|Insertion, replacement and revision of posterior spinal motion preservation device(s)
C1955537|ICD9CM|PT|88.59|Intra-operative coronary fluorescence vascular angiography
C1955537|ICD9CM|AB|88.59|Intraop cor flr vas angi
C1955541|ICD9CM|PT|92.41|Intra-operative electron radiation therapy
C1955541|ICD9CM|AB|92.41|Intra-op electron rad rx
C1955543|ICD9CM|HT|92.4|Intra-operative radiation procedures
C1955545|ICD9CM|AB|999.31|Oth/uns inf-cen ven cath
C1955545|ICD9CM|PT|999.31|Other and unspecified infection due to central venous catheter
C1955550|ICD9CM|PT|999.39|Infection following other infusion, injection, transfusion, or vaccination
C1955550|ICD9CM|AB|999.39|Infect fol infus/inj/vac
C1955551|MTH|PN|NOCODE|VEHICLE ACCIDENTS NOT ELSEWHERE CLASSIFIABLE in ICD9CM
C1955551|ICD9CM|HT|E846-E848.9|VEHICLE ACCIDENTS NOT ELSEWHERE CLASSIFIABLE
C1955553|ICD9CM|HT|040.4|Other specified botulism
C1955556|ICD9CM|PT|E928.6|Environmental exposure to harmful algae and toxins
C1955556|ICD9CM|AB|E928.6|Envir expose algae/toxin
C1955565|ICD9CM|AB|E933.6|Oral bisphosphonates
C1955565|ICD9CM|PT|E933.6|Oral bisphosphonates
C1955566|ICD9CM|PT|E933.7|Intravenous bisphosphonates
C1955566|ICD9CM|AB|E933.7|IV bisphosphonates
C1955570|ICD9CM|AB|V12.54|Hx TIA/stroke w/o resid
C1955570|ICD9CM|PT|V12.54|Personal history of transient ischemic attack (TIA), and cerebral infarction without residual deficits
C1955573|ICD9CM|PT|V13.22|Personal history of cervical dysplasia
C1955573|ICD9CM|AB|V13.22|Hx of cervical dysplasia
C1955574|ICD9CM|PT|V16.52|Family history of malignant neoplasm, bladder
C1955574|ICD9CM|AB|V16.52|Fam hx-bladder malig
C1955576|ICD9CM|AB|V18.11|Fam hx MEN syndrome
C1955576|ICD9CM|PT|V18.11|Family history of multiple endocrine neoplasia [MEN] syndrome
C1955577|ICD9CM|HT|V18.1|Family history of other endocrine and metabolic diseases
C1955577|ICD9CM|PT|V18.19|Family history of other endocrine and metabolic diseases
C1955577|ICD9CM|AB|V18.19|Fm hx endo/metab dis NEC
C1955578|ICD9CM|AB|V25.04|Natrl fam pln-avoid preg
C1955578|ICD9CM|PT|V25.04|Counseling and instruction in natural family planning to avoid pregnancy
C1955579|ICD9CM|PT|V26.41|Procreative counseling and advice using natural family planning
C1955579|ICD9CM|AB|V26.41|Natrl family plan counsl
C1955580|MTH|PN|NOCODE|Encounter for procreative management counseling and advice in ICD9CM
C1955580|ICD9CM|PT|V26.49|Other procreative management counseling and advice
C1955580|ICD9CM|AB|V26.49|Procr mgmt cnsl/adv NEC
C1955581|ICD9CM|PT|V26.81|Encounter for assisted reproductive fertility procedure cycle
C1955581|ICD9CM|AB|V26.81|Assist repro fertility
C1955583|MTH|PN|NOCODE|PROCREATIVE MANAGEMT NEC in ICD9CM_2008
C1955583|ICD9CM|PT|V26.89|Other specified procreative management
C1955583|ICD9CM|AB|V26.89|Procreative managemt NEC
C1955592|ICD9CM|PT|V49.70|Unspecified level lower limb amputation status
C1955592|ICD9CM|AB|V49.70|Status amput lwr lmb NOS
C1955593|ICD9CM|PT|V49.71|Great toe amputation status
C1955593|ICD9CM|AB|V49.71|Status amput great toe
C1955594|ICD9CM|PT|V49.72|Other toe(s) amputation status
C1955594|ICD9CM|AB|V49.72|Status amput othr toe(s)
C1955595|ICD9CM|PT|V49.73|Foot amputation status
C1955595|ICD9CM|AB|V49.73|Status amput foot
C1955596|ICD9CM|PT|V49.74|Ankle amputation status
C1955596|ICD9CM|AB|V49.74|Status amput ankle
C1955599|ICD9CM|PT|V49.77|Hip amputation status
C1955599|ICD9CM|AB|V49.77|Status amput hip
C1955601|ICD9CM|HT|V49.7|Lower limb amputation status
C1955602|ICD9CM|PT|V49.85|Dual sensory impairment
C1955602|ICD9CM|AB|V49.85|Dual sensory impairment
C1955613|ICD9CM|AB|V68.01|Disability examination
C1955613|ICD9CM|PT|V68.01|Disability examination
C1955615|ICD9CM|PT|V72.12|Encounter for hearing conservation and treatment
C1955615|ICD9CM|AB|V72.12|Hearing conservatn/trtmt
C1955616|ICD9CM|HT|V73.8|Screening examination for other specified viral and chlamydial diseases
C1955618|ICD9CM|PT|V84.81|Genetic susceptibility to multiple endocrine neoplasia [MEN]
C1955618|ICD9CM|AB|V84.81|Genetc sus mult endo neo
C1955620|ICD9CM|PT|00.18|Infusion of immunosuppressive antibody therapy
C1955620|ICD9CM|AB|00.18|Infus immunosup antibody
C1955622|ICD9CM|PT|00.19|Disruption of blood brain barrier via infusion [BBBD]
C1955622|ICD9CM|AB|00.19|BBBD via infusion
C1955624|ICD9CM|PT|00.74|Hip bearing surface, metal-on-polyethylene
C1955624|ICD9CM|AB|00.74|Hip surface, metal/poly
C1955625|ICD9CM|AB|00.75|Hip surface, metal/metal
C1955625|ICD9CM|PT|00.75|Hip bearing surface, metal-on-metal
C1955626|ICD9CM|PT|00.76|Hip bearing surface, ceramic-on-ceramic
C1955626|ICD9CM|AB|00.76|Hip surface, cermc/cermc
C1955627|ICD9CM|PT|00.77|Hip bearing surface, ceramic-on-polyethylene
C1955627|ICD9CM|AB|00.77|Hip surface, cermc/poly
C1955628|ICD9CM|HT|058|Other human herpesvirus
C1955629|ICD9CM|PT|058.21|Human herpesvirus 6 encephalitis
C1955629|ICD9CM|AB|058.21|Human herpesvir 6 enceph
C1955630|ICD9CM|PT|058.29|Other human herpesvirus encephalitis
C1955630|ICD9CM|HT|058.2|Other human herpesvirus encephalitis
C1955630|ICD9CM|AB|058.29|Human herpesvr encph NEC
C1955633|ICD9CM|PT|058.89|Other human herpesvirus infection
C1955633|ICD9CM|HT|058.8|Other human herpesvirus infections
C1955633|ICD9CM|AB|058.89|Human herpesvirs inf NEC
C1955636|ICD9CM|HT|079.8|Other specified viral and chlamydial infections in conditions classified elsewhere and of unspecified site
C1955637|ICD9CM|PT|00.94|Intra-operative neurophysiologic monitoring
C1955637|ICD9CM|AB|00.94|Intra-op neurophys montr
C1955641|ICD9CM|PT|01.16|Intracranial oxygen monitoring
C1955641|ICD9CM|AB|01.16|Intracranial 02 monitor
C1955643|ICD9CM|PT|01.17|Brain temperature monitoring
C1955643|ICD9CM|AB|01.17|Brain temp monitoring
C1955644|ICD9CM|PT|07.81|Other partial excision of thymus
C1955644|ICD9CM|AB|07.81|Oth part excision thymus
C1955646|ICD9CM|PT|07.82|Other total excision of thymus
C1955646|ICD9CM|AB|07.82|Oth totl excision thymus
C1955648|ICD9CM|PT|07.83|Thoracoscopic partial excision of thymus
C1955648|ICD9CM|AB|07.83|Thorac part exisn thymus
C1955649|ICD9CM|PT|07.84|Thoracoscopic total excision of thymus
C1955649|ICD9CM|AB|07.84|Thorac total exc thymus
C1955650|ICD9CM|AB|07.92|Other incision of thymus
C1955650|ICD9CM|PT|07.92|Other incision of thymus
C1955652|ICD9CM|PT|07.95|Thoracoscopic incision of thymus
C1955652|ICD9CM|AB|07.95|Thorac incision thymus
C1955653|ICD9CM|PT|07.98|Other and unspecified thoracoscopic operations on thymus
C1955653|ICD9CM|AB|07.98|Oth thorac op thymus NOS
C1955654|ICD9CM|PT|07.99|Other and unspecified operations on thymus
C1955654|ICD9CM|AB|07.99|Other thymus ops NOS
C1955681|ICD9CM|PT|200.30|Marginal zone lymphoma, unspecified site, extranodal and solid organ sites
C1955681|ICD9CM|AB|200.30|Margnl zone lym xtrndl
C1955682|ICD9CM|PT|200.31|Marginal zone lymphoma, lymph nodes of head, face, and neck
C1955682|ICD9CM|AB|200.31|Margin zone lym head
C1955683|ICD9CM|PT|200.32|Marginal zone lymphoma, intrathoracic lymph nodes
C1955683|ICD9CM|AB|200.32|Margin zone lym thorax
C1955684|ICD9CM|PT|200.33|Marginal zone lymphoma, intraabdominal lymph nodes
C1955684|ICD9CM|AB|200.33|Margin zone lym abdom
C1955685|ICD9CM|PT|200.34|Marginal zone lymphoma, lymph nodes of axilla and upper limb
C1955685|ICD9CM|AB|200.34|Margin zone lym axilla
C1955686|ICD9CM|PT|200.35|Marginal zone lymphoma, lymph nodes of inguinal region and lower limb
C1955686|ICD9CM|AB|200.35|Margin zone lym inguin
C1955687|ICD9CM|PT|200.36|Marginal zone lymphoma, intrapelvic lymph nodes
C1955687|ICD9CM|AB|200.36|Margin zone lym pelvic
C1955689|ICD9CM|PT|200.38|Marginal zone lymphoma, lymph nodes of multiple sites
C1955689|ICD9CM|AB|200.38|Margin zone lymph multip
C1955691|ICD9CM|PT|200.40|Mantle cell lymphoma, unspecified site, extranodal and solid organ sites
C1955691|ICD9CM|AB|200.40|Mantle cell lym xtrrndl
C1955700|ICD9CM|PT|200.50|Primary central nervous system lymphoma, unspecified site, extranodal and solid organ sites
C1955700|ICD9CM|AB|200.50|Primary CNS lymph xtrndl
C1955701|ICD9CM|PT|200.51|Primary central nervous system lymphoma, lymph nodes of head, face, and neck
C1955701|ICD9CM|AB|200.51|Primary CNS lymph head
C1955702|ICD9CM|PT|200.52|Primary central nervous system lymphoma, intrathoracic lymph nodes
C1955702|ICD9CM|AB|200.52|Primary CNS lymph thorax
C1955703|ICD9CM|PT|200.53|Primary central nervous system lymphoma, intra-abdominal lymph nodes
C1955703|ICD9CM|AB|200.53|Primary CNS lymph abdom
C1955704|ICD9CM|PT|200.54|Primary central nervous system lymphoma, lymph nodes of axilla and upper limb
C1955704|ICD9CM|AB|200.54|Primary CNS lymph axilla
C1955705|ICD9CM|PT|200.55|Primary central nervous system lymphoma, lymph nodes of inguinal region and lower limb
C1955705|ICD9CM|AB|200.55|Primary CNS lym inguin
C1955706|ICD9CM|PT|200.56|Primary central nervous system lymphoma, intrapelvic lymph nodes
C1955706|ICD9CM|AB|200.56|Primary CNS lymph pelvic
C1955707|ICD9CM|PT|200.57|Primary central nervous system lymphoma, spleen
C1955707|ICD9CM|AB|200.57|Primary CNS lymph spleen
C1955708|ICD9CM|PT|200.58|Primary central nervous system lymphoma, lymph nodes of multiple sites
C1955708|ICD9CM|AB|200.58|Primary CNS lymph multip
C1955709|ICD9CM|PT|200.60|Anaplastic large cell lymphoma, unspecified site, extranodal and solid organ sites
C1955709|ICD9CM|AB|200.60|Anaplastic lymph xtrndl
C1955710|ICD9CM|PT|200.61|Anaplastic large cell lymphoma, lymph nodes of head, face, and neck
C1955710|ICD9CM|AB|200.61|Anaplastic lymph head
C1955711|ICD9CM|PT|200.62|Anaplastic large cell lymphoma, intrathoracic lymph nodes
C1955711|ICD9CM|AB|200.62|Anaplastic lymph thorax
C1955712|ICD9CM|PT|200.63|Anaplastic large cell lymphoma, intra-abdominal lymph nodes
C1955712|ICD9CM|AB|200.63|Anaplastic lymph abdom
C1955713|ICD9CM|PT|200.64|Anaplastic large cell lymphoma, lymph nodes of axilla and upper limb
C1955713|ICD9CM|AB|200.64|Anaplastic lymph axilla
C1955714|ICD9CM|PT|200.65|Anaplastic large cell lymphoma, lymph nodes of inguinal region and lower limb
C1955714|ICD9CM|AB|200.65|Anaplastic lymph inguin
C1955715|ICD9CM|PT|200.66|Anaplastic large cell lymphoma, intrapelvic lymph nodes
C1955715|ICD9CM|AB|200.66|Anaplastic lymph pelvic
C1955717|ICD9CM|PT|200.68|Anaplastic large cell lymphoma, lymph nodes of multiple sites
C1955717|ICD9CM|AB|200.68|Anaplastic lymph multip
C1955718|ICD9CM|PT|200.70|Large cell lymphoma, unspecified site, extranodal and solid organ sites
C1955718|ICD9CM|AB|200.70|Large cell lymph xtrndl
C1955719|ICD9CM|PT|200.71|Large cell lymphoma, lymph nodes of head, face, and neck
C1955719|ICD9CM|AB|200.71|Large cell lymphoma head
C1955720|ICD9CM|PT|200.72|Large cell lymphoma, intrathoracic lymph nodes
C1955720|ICD9CM|AB|200.72|Large cell lymph thorax
C1955721|ICD9CM|PT|200.73|Large cell lymphoma, intra-abdominal lymph nodes
C1955721|ICD9CM|AB|200.73|Large cell lymph abdom
C1955722|ICD9CM|PT|200.74|Large cell lymphoma, lymph nodes of axilla and upper limb
C1955722|ICD9CM|AB|200.74|Large cell lymph axilla
C1955723|ICD9CM|PT|200.75|Large cell lymphoma, lymph nodes of inguinal region and lower limb
C1955723|ICD9CM|AB|200.75|Large cell lymph inguin
C1955725|ICD9CM|PT|200.77|Large cell lymphoma, spleen
C1955725|ICD9CM|AB|200.77|Large cell lymph spleen
C1955726|ICD9CM|PT|200.78|Large cell lymphoma, lymph nodes of multiple sites
C1955726|ICD9CM|AB|200.78|Large cell lymph multip
C1955727|ICD9CM|HT|200|Lymphosarcoma and reticulosarcoma and other specified malignant tumors of lymphatic tissue
C1955728|ICD9CM|PT|202.70|Peripheral T cell lymphoma, unspecified site, extranodal and solid organ sites
C1955728|ICD9CM|AB|202.70|Periph T cell lym xtrndl
C1955730|ICD9CM|PT|202.72|Peripheral T cell lymphoma, intrathoracic lymph nodes
C1955730|ICD9CM|AB|202.72|Periph T cell lym thorax
C1955735|ICD9CM|PT|202.77|Peripheral T cell lymphoma, spleen
C1955735|ICD9CM|AB|202.77|Periph T cell lym spleen
C1955737|ICD9CM|PT|233.30|Carcinoma in situ, unspecified female genital organ
C1955737|ICD9CM|AB|233.30|Ca in situ fem gen NOS
C1955739|ICD9CM|PT|233.39|Carcinoma in situ, other female genital organ
C1955739|ICD9CM|AB|233.39|Ca in situ fem gen NEC
C1955741|ICD9CM|PT|255.41|Glucocorticoid deficiency
C1955741|ICD9CM|AB|255.41|Glucocorticoid deficient
C1955743|ICD9CM|PT|255.42|Mineralocorticoid deficiency
C1955743|ICD9CM|AB|255.42|Mineralcorticoid defcnt
C1955746|MTH|PN|NOCODE|APLASTIC ANEMIAS NEC in ICD9CM
C1955746|ICD9CM|AB|284.89|Aplastic anemias NEC
C1955746|ICD9CM|PT|284.89|Other specified aplastic anemias
C1955750|ICD9CM|PT|315.34|Speech and language developmental delay due to hearing loss
C1955750|ICD9CM|AB|315.34|Speech del d/t hear loss
C1955751|ICD9CM|PT|32.20|Thoracoscopic excision of lesion or tissue of lung
C1955751|ICD9CM|AB|32.20|Thorac exc lung lesion
C1955753|ICD9CM|PT|32.30|Thoracoscopic segmental resection of lung
C1955753|ICD9CM|AB|32.30|Thorac seg lung resect
C1955754|ICD9CM|PT|32.39|Other and unspecified segmental resection of lung
C1955754|ICD9CM|AB|32.39|Oth seg lung resect NOS
C1955755|ICD9CM|PT|32.49|Other lobectomy of lung
C1955755|ICD9CM|AB|32.49|Lobectomy of lung NEC
C1955756|ICD9CM|PT|32.59|Other and unspecified pneumonectomy
C1955756|ICD9CM|AB|32.59|Other pneumonectomy NOS
C1955760|ICD9CM|PT|331.5|Idiopathic normal pressure hydrocephalus (INPH)
C1955760|ICD9CM|AB|331.5|Norml pressure hydroceph
C1955761|ICD9CM|PT|34.06|Thoracoscopic drainage of pleural cavity
C1955761|ICD9CM|AB|34.06|Thorac drain pleurl cav
C1955763|MTH|PN|NOCODE|PLEURAL BIOPSY NEC in ICD9CM_2008
C1955763|ICD9CM|PT|34.24|Other pleural biopsy
C1955763|ICD9CM|AB|34.24|Pleural biopsy NEC
C1955764|ICD9CM|PT|34.52|Thoracoscopic decortication of lung
C1955764|ICD9CM|AB|34.52|Thoracoscopc decort lung
C1955771|ICD9CM|PT|388.45|Acquired auditory processing disorder
C1955771|ICD9CM|AB|388.45|Acq auditory process dis
C1955772|ICD9CM|PT|389.05|Conductive hearing loss, unilateral
C1955772|ICD9CM|AB|389.05|Condctv hear loss,unilat
C1955773|ICD9CM|PT|389.13|Neural hearing loss, unilateral
C1955773|ICD9CM|AB|389.13|Neural hear loss, unilat
C1955774|ICD9CM|PT|389.17|Sensory hearing loss, unilateral
C1955774|ICD9CM|AB|389.17|Sensory hear loss,unilat
C1955775|ICD9CM|PT|389.21|Mixed hearing loss, unilateral
C1955775|ICD9CM|AB|389.21|Mixed hearing loss,unilt
C1955777|ICD9CM|PT|389.7|Deaf, nonspeaking, not elsewhere classifiable
C1955777|ICD9CM|AB|389.7|Deaf, nonspeaking NEC
C1955779|ICD9CM|PT|414.2|Chronic total occlusion of coronary artery
C1955779|ICD9CM|AB|414.2|Chr tot occlus cor artry
C1955781|ICD9CM|PT|415.12|Septic pulmonary embolism
C1955781|ICD9CM|AB|415.12|Septic pulmonary embolsm
C1955783|ICD9CM|AB|440.4|Chr tot occl art extrem
C1955783|ICD9CM|PT|440.4|Chronic total occlusion of artery of the extremities
C1955786|ICD9CM|PT|449|Septic arterial embolism
C1955786|ICD9CM|AB|449|Septic arterial embolism
C1955790|ICD9CM|PT|50.13|Transjugular liver biopsy
C1955790|ICD9CM|AB|50.13|Transjugular liver bx
C1955799|ICD9CM|PT|525.72|Post-osseointegration biological failure of dental implant
C1955799|ICD9CM|AB|525.72|Post-osse biol fail impl
C1955807|ICD9CM|PT|525.73|Post-osseointegration mechanical failure of dental implant
C1955807|ICD9CM|AB|525.73|Post-osse mech fail impl
C1955810|ICD9CM|PT|525.79|Other endosseous dental implant failure
C1955810|ICD9CM|AB|525.79|Endos dentl imp fail NEC
C1955812|ICD9CM|HT|525.7|Endosseous dental implant failure
C1955814|ICD9CM|PT|569.43|Anal sphincter tear (healed) (old)
C1955814|ICD9CM|AB|569.43|Anal sphincter tear-old
C1955816|ICD9CM|PT|624.09|Other dystrophy of vulva
C1955816|ICD9CM|AB|624.09|Dystrophy of vulva NEC
C1959600|ICD9CM|PT|425.2|Obscure cardiomyopathy of Africa
C1959600|ICD9CM|AB|425.2|Obsc afric cardiomyopath
C1959635|ICD9CM|AB|079.83|Parvovirus B19
C1959635|ICD9CM|PT|079.83|Parvovirus B19
C1959639|ICD9CM|PT|V73.81|Special screening examination for Human papillomavirus (HPV)
C1959639|ICD9CM|AB|V73.81|Special screen exam HPV
C1961101|MTH|PN|NOCODE|BLADDER CALCULUS NEC in ICD9CM
C1961101|ICD9CM|PT|594.1|Other calculus in bladder
C1961101|ICD9CM|AB|594.1|Bladder calculus NEC
C1961111|MTH|PN|NOCODE|Tremor NEC in ICD9CM_2014
C1961111|ICD9CM|PT|333.1|Essential and other specified forms of tremor
C1961111|ICD9CM|AB|333.1|Tremor NEC
C1961116|ICD9CM|AB|V12.53|Hx sudden cardiac arrest
C1961116|ICD9CM|PT|V12.53|Personal history of sudden cardiac arrest
C1961121|ICD9CM|PT|743.58|Vascular anomalies
C1961121|ICD9CM|AB|743.58|Vascular anom post eye
C1961127|MTH|PN|NOCODE|Screening examination for venereal disease in ICD9CM_2008
C1961127|ICD9CM|PT|V74.5|Screening examination for venereal disease
C1961127|ICD9CM|AB|V74.5|Screen for veneral dis
C1961128|MTH|PN|NOCODE|Encounter for tuboplasty or vasoplasty after previous sterilization in ICD9CM_2008
C1961128|ICD9CM|PT|V26.0|Tuboplasty or vasoplasty after previous sterilization
C1961128|ICD9CM|AB|V26.0|Tuboplasty or vasoplasty
C1961134|MTH|PN|NOCODE|Encounter for examination of eyes and vision in ICD9CM_2008
C1961134|ICD9CM|PT|V72.0|Examination of eyes and vision
C1961134|ICD9CM|AB|V72.0|Eye & vision examination
C1961834|ICD9CM|PT|533.70|Chronic peptic ulcer of unspecified site without mention of hemorrhage or perforation, without mention of obstruction
C1961834|ICD9CM|AB|533.70|Chronic peptic ulcer NOS
C1961841|MTH|PN|NOCODE|MYELOPATHY NEC in ICD9CM
C1961841|ICD9CM|PT|336.8|Other myelopathy
C1961841|ICD9CM|AB|336.8|Myelopathy NEC
C1962919|MTH|PN|NOCODE|Encounter for screening for chromosomal anomalies by amniocentesis in ICD9CM
C1962919|ICD9CM|PT|V28.0|Antenatal screening for chromosomal anomalies by amniocentesis
C1962919|ICD9CM|AB|V28.0|Screening-chromosom anom
C1962929|MTH|PN|NOCODE|SLEEP DISTURBANCES NEC in ICD9CM
C1962929|ICD9CM|PT|780.59|Other sleep disturbances
C1962929|ICD9CM|AB|780.59|Sleep disturbances NEC
C1962938|MTH|PN|NOCODE|Need for prophylactic vaccination and inoculation against arthropod-borne viral encephalitis in ICD9CM (finding)
C1962938|ICD9CM|PT|V05.0|Need for prophylactic vaccination and inoculation against arthropod-borne viral encephalitis
C1962938|ICD9CM|AB|V05.0|Arbovirus enceph vaccin
C1962940|MTH|PN|NOCODE|Need for prophylactic vaccination and inoculation against poliomyelitis in ICD9CM
C1962940|ICD9CM|PT|V04.0|Need for prophylactic vaccination and inoculation against poliomyelitis
C1962940|ICD9CM|AB|V04.0|Vaccin for poliomyelitis
C1963536|ICD9CM|HT|747.6|Other congenital anomalies of peripheral vascular system
C1963544|ICD9CM|PT|718.57|Ankylosis of joint, ankle and foot
C1963544|ICD9CM|AB|718.57|Ankylosis-ankle
C1963546|ICD9CM|HT|825|Fracture of one or more tarsal and metatarsal bones
C1963551|ICD9CM|HT|68.6|Radical abdominal hysterectomy
C1963552|ICD9CM|PT|730.05|Acute osteomyelitis, pelvic region and thigh
C1963552|ICD9CM|AB|730.05|Ac osteomyelitis-pelvis
C1963664|ICD9CM|PT|718.47|Contracture of joint, ankle and foot
C1963664|ICD9CM|AB|718.47|Jt contracture-ankle
C1963706|MTH|PN|NOCODE|Family history of other cardiovascular diseases in ICD9CM
C1963706|ICD9CM|HT|V17.4|Family history of other cardiovascular diseases
C1963707|MTH|PN|NOCODE|Family history of other cardiovascular diseases NEC in ICD9CM
C1963707|ICD9CM|PT|V17.49|Family history of other cardiovascular diseases
C1963707|ICD9CM|AB|V17.49|Fam hx-cardiovas dis NEC
C1963710|MTH|PN|NOCODE|Antidotes and chelating agents, not elsewhere classified, causing adverse effects in therapeutic use in ICD9CM
C1963710|ICD9CM|PT|E947.2|Antidotes and chelating agents, not elsewhere classified, causing adverse effects in therapeutic use
C1963710|ICD9CM|AB|E947.2|Adv eff antidotes NEC
C1970956|ICD9CM|PT|20.01|Myringotomy with insertion of tube
C1970956|ICD9CM|AB|20.01|Myringotomy w intubation
C1970969|ICD9CM|HT|32|Excision of lung and bronchus
C1971612|MTH|PN|NOCODE|Encounter for occupational therapy in ICD9CM
C1971612|ICD9CM|PT|V57.21|Encounter for occupational therapy
C1971612|ICD9CM|AB|V57.21|Encntr occupatnal thrpy
C1971613|ICD9CM|PT|V50.2|Routine or ritual circumcision
C1971613|ICD9CM|AB|V50.2|Routine circumcision
C1971617|ICD9CM|PT|V52.2|Fitting and adjustment of artificial eye
C1971617|ICD9CM|AB|V52.2|Fitting artificial eye
C1971635|ICD9CM|HT|379.0|Scleritis and episcleritis
C1997588|ICD9CM|PT|323.52|Myelitis following immunization procedures
C1997588|ICD9CM|AB|323.52|Myelitis follwg immune
C1997777|ICD9CM|PT|608.24|Torsion of appendix epididymis
C1997777|ICD9CM|AB|608.24|Torsion appy epididymis
C1998428|ICD9CM|PT|292.84|Drug-induced mood disorder
C1998428|ICD9CM|AB|292.84|Drug-induced mood disord
C1998978|ICD9CM|PT|783.7|Adult failure to thrive
C1998978|ICD9CM|AB|783.7|Failure to thrive-adult
C2003945|ICD9CM|HT|768|Intrauterine hypoxia and birth asphyxia
C2004369|ICD9CM|PT|750.7|Other specified anomalies of stomach
C2004369|ICD9CM|AB|750.7|Gastric anomaly NEC
C2004376|ICD9CM|PT|727.05|Other tenosynovitis of hand and wrist
C2004376|ICD9CM|AB|727.05|Tenosynov hand/wrist NEC
C2004435|ICD9CM|HT|557|Vascular insufficiency of intestine
C2004435|ICD9CM|PT|557.9|Unspecified vascular insufficiency of intestine
C2004435|ICD9CM|AB|557.9|Vasc insuff intest NOS
C2004459|ICD9CM|HT|48.5|Abdominoperineal resection of rectum
C2004465|ICD9CM|PT|750.9|Unspecified anomaly of upper alimentary tract
C2004465|ICD9CM|AB|750.9|Upper GI anomaly NOS
C2004477|ICD9CM|PT|377.52|Disorders of optic chiasm associated with other neoplasms
C2004477|ICD9CM|AB|377.52|Opt chiasm dis/neopl NEC
C2004479|ICD9CM|HT|671.1|Varicose veins of vulva and perineum in pregnancy and the puerperium
C2004481|ICD9CM|PT|163.0|Malignant neoplasm of parietal pleura
C2004481|ICD9CM|AB|163.0|Mal neo parietal pleura
C2004482|ICD9CM|HT|941|Burn of face, head, and neck
C2004487|ICD9CM|AB|625.1|Vaginismus
C2004487|ICD9CM|PT|625.1|Vaginismus
C2004488|ICD9CM|AB|43.3|Pyloromyotomy
C2004488|ICD9CM|PT|43.3|Pyloromyotomy
C2004518|ICD9CM|HT|790-796.99|NONSPECIFIC ABNORMAL FINDINGS
C2018768|ICD9CM|PT|200.67|Anaplastic large cell lymphoma, spleen
C2018768|ICD9CM|AB|200.67|Anaplastic lymph spleen
C2018777|ICD9CM|PT|200.47|Mantle cell lymphoma, spleen
C2018777|ICD9CM|AB|200.47|Mantle cell lymph spleen
C2039668|ICD9CM|PT|090.3|Syphilitic interstitial keratitis
C2039668|ICD9CM|AB|090.3|Syphilitic keratitis
C2047520|ICD9CM|AB|272.2|Mixed hyperlipidemia
C2047520|ICD9CM|PT|272.2|Mixed hyperlipidemia
C2053058|ICD9CM|PT|81.66|Percutaneous vertebral augmentation
C2053058|ICD9CM|AB|81.66|Percut vertebral augment
C2053768|ICD9CM|PT|955.8|Injury to multiple nerves of shoulder girdle and upper limb
C2053768|ICD9CM|AB|955.8|Inj mult nerve shldr/arm
C2062527|ICD9CM|HT|209.0|Malignant carcinoid tumors of the small intestine
C2062529|ICD9CM|PT|209.11|Malignant carcinoid tumor of the appendix
C2062529|ICD9CM|AB|209.11|Malig carcinoid appendix
C2062573|ICD9CM|PT|209.23|Malignant carcinoid tumor of the stomach
C2062573|ICD9CM|AB|209.23|Malig carcinoid stomach
C2077104|ICD9CM|HT|E979|Terrorism
C2077104|ICD9CM|HT|E979-E979.9|TERRORISM
C2114658|ICD9CM|PT|658.91|Unspecified problem associated with amniotic cavity and membranes, delivered, with or without mention of antepartum condition
C2114658|ICD9CM|AB|658.91|Amniotic prob NOS-deliv
C2127287|ICD9CM|PT|789.45|Abdominal rigidity, periumbilic
C2127287|ICD9CM|AB|789.45|Abdmnal rgdt periumbilic
C2163761|ICD9CM|AB|12.72|Cyclocryotherapy
C2163761|ICD9CM|PT|12.72|Cyclocryotherapy
C2170463|ICD9CM|PT|37.53|Replacement or repair of thoracic unit of (total) replacement heart system
C2170463|ICD9CM|AB|37.53|Repl/rep thr unt tot hrt
C2183395|ICD9CM|PT|569.86|Dieulafoy lesion (hemorrhagic) of intestine
C2183395|ICD9CM|AB|569.86|Dieulafoy les, intestine
C2186390|ICD9CM|AB|V43.61|Joint replaced shoulder
C2186390|ICD9CM|PT|V43.61|Shoulder joint replacement
C2188200|ICD9CM|PT|525.62|Unrepairable overhanging of dental restorative materials
C2188200|ICD9CM|AB|525.62|Overhang dental restore
C2193446|ICD9CM|PT|13.41|Phacoemulsification and aspiration of cataract
C2193446|ICD9CM|AB|13.41|Catarac phacoemuls/aspir
C2197988|ICD9CM|PT|312.22|Socialized conduct disorder, moderate
C2197988|ICD9CM|AB|312.22|Social conduct dis-mod
C2205119|ICD9CM|PT|209.17|Malignant carcinoid tumor of the rectum
C2205119|ICD9CM|AB|209.17|Malig carcinoid rectum
C2223867|ICD9CM|AB|24.31|Gum lesion excision
C2223867|ICD9CM|PT|24.31|Excision of lesion or tissue of gum
C2227090|ICD9CM|AB|524.01|Maxillary hyperplasia
C2227090|ICD9CM|PT|524.01|Major anomalies of jaw size, maxillary hyperplasia
C2228890|ICD9CM|PT|996.57|Mechanical complication due to insulin pump
C2228890|ICD9CM|AB|996.57|Complcation-insulin pump
C2231357|ICD9CM|PT|312.21|Socialized conduct disorder, mild
C2231357|ICD9CM|AB|312.21|Social conduct dis-mild
C2231358|ICD9CM|PT|312.23|Socialized conduct disorder, severe
C2231358|ICD9CM|AB|312.23|Social conduct dis-sev
C2233848|ICD9CM|PT|611.81|Ptosis of breast
C2233848|ICD9CM|AB|611.81|Ptosis of breast
C2239098|ICD9CM|PT|736.73|Cavus deformity of foot, acquired
C2239098|ICD9CM|AB|736.73|Cavus deformity of foot
C2239106|ICD9CM|HT|363.2|Other and unspecified forms of chorioretinitis and retinochoroiditis
C2239133|ICD9CM|PT|57.33|Closed [transurethral] biopsy of bladder
C2239133|ICD9CM|AB|57.33|Clos transureth bladd bx
C2239162|ICD9CM|AB|84.47|Fit leg prosthesis NOS
C2239162|ICD9CM|PT|84.47|Fitting of prosthesis of leg, not otherwise specified
C2240369|ICD9CM|PT|V45.01|Cardiac pacemaker in situ
C2240369|ICD9CM|AB|V45.01|Status cardiac pacemaker
C2240388|ICD9CM|PT|058.11|Roseola infantum due to human herpesvirus 6
C2240388|ICD9CM|AB|058.11|Roseola infant d/t HHV-6
C2240395|ICD9CM|PT|909.9|Late effect of other and unspecified external causes
C2240395|ICD9CM|AB|909.9|Late eff exter cause NEC
C2240397|ICD9CM|PT|994.9|Other effects of external causes
C2240397|ICD9CM|AB|994.9|Effect external caus NEC
C2240398|ICD9CM|PT|996.96|Complication of reattached lower extremity, other and unspecified
C2240398|ICD9CM|AB|996.96|Compl reattached leg NEC
C2240399|ICD9CM|HT|V85-V85.99|BODY MASS INDEX
C2240399|ICD9CM|HT|V85|Body mass index [BMI]
C2242472|ICD9CM|HT|730.9|Unspecified infection of bone
C2242472|ICD9CM|PT|730.90|Unspecified infection of bone, site unspecified
C2242472|ICD9CM|AB|730.90|Bone infec NOS-unsp site
C2242475|ICD9CM|PT|730.94|Unspecified infection of bone, hand
C2242475|ICD9CM|AB|730.94|Bone infect NOS-hand
C2242765|ICD9CM|PT|738.4|Acquired spondylolisthesis
C2242765|ICD9CM|AB|738.4|Acq spondylolisthesis
C2242834|ICD9CM|AB|766.0|Exceptionally large baby
C2242834|ICD9CM|PT|766.0|Exceptionally large baby
C2242854|ICD9CM|PT|230.5|Carcinoma in situ of anal canal
C2242854|ICD9CM|AB|230.5|Ca in situ anal canal
C2243036|ICD9CM|PT|34.03|Reopening of recent thoracotomy site
C2243036|ICD9CM|AB|34.03|Reopen thoracotomy site
C2243087|ICD9CM|PT|535.01|Acute gastritis, with hemorrhage
C2243087|ICD9CM|AB|535.01|Acute gastritis w hmrhg
C2266788|ICD9CM|AB|704.42|Trichilemmal cyst
C2266788|ICD9CM|PT|704.42|Trichilemmal cyst
C2267227|ICD9CM|AB|307.51|Bulimia nervosa
C2267227|ICD9CM|PT|307.51|Bulimia nervosa
C2315695|ICD9CM|PT|389.12|Neural hearing loss, bilateral
C2315695|ICD9CM|AB|389.12|Neural hearng loss,bilat
C2315800|ICD9CM|PT|787.21|Dysphagia, oral phase
C2315800|ICD9CM|AB|787.21|Dysphagia, oral phase
C2316057|ICD9CM|PT|323.72|Toxic myelitis
C2316057|ICD9CM|AB|323.72|Toxic myelitis
C2316460|ICD9CM|AB|310.81|Pseudobulbar affect
C2316460|ICD9CM|PT|310.81|Pseudobulbar affect
C2316590|ICD9CM|AB|770.81|Primary apnea of newborn
C2316590|ICD9CM|PT|770.81|Primary apnea of newborn
C2316692|ICD9CM|PT|770.88|Hypoxemia of newborn
C2316692|ICD9CM|AB|770.88|NB hypoxia
C2317110|ICD9CM|PT|733.98|Stress fracture of pelvis
C2317110|ICD9CM|AB|733.98|Stress fx pelvis
C2349213|ICD9CM|PT|00.49|Supersaturated oxygen therapy
C2349213|ICD9CM|AB|00.49|SuperSat O2 therapy
C2349215|ICD9CM|PT|00.58|Insertion of intra-aneurysm sac pressure monitoring device (intraoperative)
C2349215|ICD9CM|AB|00.58|Ins intra-ansm pres mntr
C2349217|ICD9CM|PT|00.59|Intravascular pressure measurement of coronary arteries
C2349217|ICD9CM|AB|00.59|Intravasc msmnt cor art
C2349218|ICD9CM|PT|00.67|Intravascular pressure measurement of intrathoracic arteries
C2349218|ICD9CM|AB|00.67|Intravas msmnt thorc art
C2349221|ICD9CM|PT|00.68|Intravascular pressure measurement of peripheral arteries
C2349221|ICD9CM|AB|00.68|Intravas msmt periph art
C2349225|ICD9CM|PT|00.69|Intravascular pressure measurement, other specified and unspecified vessels
C2349225|ICD9CM|AB|00.69|Intravs msmt ves NEC/NOS
C2349230|ICD9CM|PT|136.21|Specific infection due to acanthamoeba
C2349230|ICD9CM|AB|136.21|Infectn d/t acanthamoeba
C2349231|ICD9CM|PT|136.29|Other specific infections by free-living amebae
C2349231|ICD9CM|AB|136.29|Infc free-liv amebae NEC
C2349232|ICD9CM|HT|17-17.99|OTHER MISCELLANEOUS DIAGNOSTIC AND THERAPEUTIC PROCEDURES
C2349233|ICD9CM|PT|17.11|Laparoscopic repair of direct inguinal hernia with graft or prosthesis
C2349233|ICD9CM|AB|17.11|Lap dir ing hern-graft
C2349235|ICD9CM|PT|17.12|Laparoscopic repair of indirect inguinal hernia with graft or prosthesis
C2349235|ICD9CM|AB|17.12|Lap indir ing hern-graft
C2349236|ICD9CM|PT|17.13|Laparoscopic repair of inguinal hernia with graft or prosthesis, not otherwise specified
C2349236|ICD9CM|AB|17.13|Lap ing hern-graft NOS
C2349237|ICD9CM|PT|17.21|Laparoscopic bilateral repair of direct inguinal hernia with graft or prosthesis
C2349237|ICD9CM|AB|17.21|Lap bil dir ing hrn-grft
C2349238|ICD9CM|PT|17.22|Laparoscopic bilateral repair of indirect inguinal hernia with graft or prosthesis
C2349238|ICD9CM|AB|17.22|Lap bi indir ing hrn-grf
C2349239|ICD9CM|PT|17.23|Laparoscopic bilateral repair of inguinal hernia, one direct and one indirect, with graft or prosthesis
C2349239|ICD9CM|AB|17.23|Lap bi dr/ind ing hrn-gr
C2349240|ICD9CM|PT|17.24|Laparoscopic bilateral repair of inguinal hernia with graft or prosthesis, not otherwise specified
C2349240|ICD9CM|AB|17.24|Lap bil ing hern-grf NOS
C2349241|ICD9CM|PT|17.31|Laparoscopic multiple segmental resection of large intestine
C2349241|ICD9CM|AB|17.31|Lap mul seg res lg intes
C2349242|ICD9CM|AB|17.32|Laparoscopic cecectomy
C2349242|ICD9CM|PT|17.32|Laparoscopic cecectomy
C2349243|ICD9CM|PT|17.34|Laparoscopic resection of transverse colon
C2349243|ICD9CM|AB|17.34|Lap res transverse colon
C2349244|ICD9CM|PT|17.35|Laparoscopic left hemicolectomy
C2349244|ICD9CM|AB|17.35|Lap left hemicolectomy
C2349246|ICD9CM|PT|17.39|Other laparoscopic partial excision of large intestine
C2349246|ICD9CM|AB|17.39|Lap pt ex lrg intest NEC
C2349247|ICD9CM|HT|17.3|Laparoscopic partial excision of large intestine
C2349248|ICD9CM|PT|17.41|Open robotic assisted procedure
C2349248|ICD9CM|AB|17.41|Open robotic assist proc
C2349249|ICD9CM|PT|17.42|Laparoscopic robotic assisted procedure
C2349249|ICD9CM|AB|17.42|Lap robotic assist proc
C2349250|ICD9CM|PT|17.43|Percutaneous robotic assisted procedure
C2349250|ICD9CM|AB|17.43|Perc robotic assist proc
C2349251|ICD9CM|PT|17.44|Endoscopic robotic assisted procedure
C2349251|ICD9CM|AB|17.44|Endo robotic assist proc
C2349252|ICD9CM|PT|17.45|Thoracoscopic robotic assisted procedure
C2349252|ICD9CM|AB|17.45|Thoraco robotic ast proc
C2349253|ICD9CM|PT|17.49|Other and unspecified robotic assisted procedure
C2349253|ICD9CM|AB|17.49|Robotic ast proc NEC/NOS
C2349254|ICD9CM|HT|17.4|Robotic assisted procedures
C2349259|ICD9CM|PT|199.2|Malignant neoplasm associated with transplant organ
C2349259|ICD9CM|AB|199.2|Malig neopl-transp organ
C2349260|ICD9CM|PT|203.00|Multiple myeloma, without mention of having achieved remission
C2349260|ICD9CM|AB|203.00|Mult mye w/o achv rmson
C2349261|ICD9CM|PT|203.02|Multiple myeloma, in relapse
C2349261|ICD9CM|AB|203.02|Mult myeloma in relapse
C2349262|ICD9CM|PT|203.10|Plasma cell leukemia, without mention of having achieved remission
C2349262|ICD9CM|AB|203.10|Pls cl leu w/o achv rmsn
C2349263|ICD9CM|PT|203.12|Plasma cell leukemia, in relapse
C2349263|ICD9CM|AB|203.12|Plsm cel leuk in relapse
C2349264|ICD9CM|PT|203.80|Other immunoproliferative neoplasms, without mention of having achieved remission
C2349264|ICD9CM|AB|203.80|Oth imno npl wo ach rmsn
C2349265|ICD9CM|PT|203.82|Other immunoproliferative neoplasms, in relapse
C2349265|ICD9CM|AB|203.82|Oth imnprlf neo-relapse
C2349266|ICD9CM|PT|204.00|Acute lymphoid leukemia, without mention of having achieved remission
C2349266|ICD9CM|AB|204.00|Ac lym leuk wo achv rmsn
C2349267|ICD9CM|PT|204.02|Acute lymphoid leukemia, in relapse
C2349267|ICD9CM|AB|204.02|Act lymp leuk in relapse
C2349268|ICD9CM|PT|204.10|Chronic lymphoid leukemia, without mention of having achieved remission
C2349268|ICD9CM|AB|204.10|Ch lym leuk wo achv rmsn
C2349269|ICD9CM|PT|204.20|Subacute lymphoid leukemia, without mention of having achieved remission
C2349269|ICD9CM|AB|204.20|Sbac lym leu wo ach rmsn
C2349270|ICD9CM|PT|204.22|Subacute lymphoid leukemia, in relapse
C2349270|ICD9CM|AB|204.22|Sbac lym leuk in relapse
C2349271|ICD9CM|PT|204.80|Other lymphoid leukemia, without mention of having achieved remission
C2349271|ICD9CM|AB|204.80|Oth lym leu wo achv rmsn
C2349272|ICD9CM|PT|204.82|Other lymphoid leukemia, in relapse
C2349272|ICD9CM|AB|204.82|Oth lym leuk in relapse
C2349273|ICD9CM|PT|204.90|Unspecified lymphoid leukemia, without mention of having achieved remission
C2349273|ICD9CM|AB|204.90|Uns lym leu wo ach rmsn
C2349274|ICD9CM|PT|204.92|Unspecified lymphoid leukemia, in relapse
C2349274|ICD9CM|AB|204.92|Lymp leuk NOS relapse
C2349275|ICD9CM|PT|205.00|Acute myeloid leukemia, without mention of having achieved remission
C2349275|ICD9CM|AB|205.00|Ac myl leuk wo achv rmsn
C2349276|ICD9CM|PT|205.02|Acute myeloid leukemia, in relapse
C2349276|ICD9CM|AB|205.02|Act myel leuk in relapse
C2349277|ICD9CM|PT|205.10|Chronic myeloid leukemia, without mention of having achieved remission
C2349277|ICD9CM|AB|205.10|Ch myl leuk wo achv rmsn
C2349278|ICD9CM|PT|205.20|Subacute myeloid leukemia, without mention of having achieved remission
C2349278|ICD9CM|AB|205.20|Sbac myl leu wo ach rmsn
C2349279|ICD9CM|PT|205.22|Subacute myeloid leukemia, in relapse
C2349279|ICD9CM|AB|205.22|Sbac myl leuk in relapse
C2349280|ICD9CM|PT|205.30|Myeloid sarcoma, without mention of having achieved remission
C2349280|ICD9CM|AB|205.30|Myl sarcoma wo achv rmsn
C2349281|ICD9CM|PT|205.32|Myeloid sarcoma, in relapse
C2349281|ICD9CM|AB|205.32|Myel sarcoma in relapse
C2349282|ICD9CM|PT|205.80|Other myeloid leukemia, without mention of having achieved remission
C2349282|ICD9CM|AB|205.80|Oth my leuk wo achv rmsn
C2349283|ICD9CM|PT|205.82|Other myeloid leukemia, in relapse
C2349283|ICD9CM|AB|205.82|Oth myel leuk in relapse
C2349284|ICD9CM|PT|205.90|Unspecified myeloid leukemia, without mention of having achieved remission
C2349284|ICD9CM|AB|205.90|Uns my leu wo ach rmsn
C2349285|ICD9CM|PT|205.92|Unspecified myeloid leukemia, in relapse
C2349285|ICD9CM|AB|205.92|Myel leuk NOS in relapse
C2349286|ICD9CM|PT|206.00|Acute monocytic leukemia, without mention of having achieved remission
C2349286|ICD9CM|AB|206.00|Ac mono leu wo achv rmsn
C2349287|ICD9CM|PT|206.02|Acute monocytic leukemia, in relapse
C2349287|ICD9CM|AB|206.02|Act mono leuk in relapse
C2349288|ICD9CM|PT|206.10|Chronic monocytic leukemia, without mention of having achieved remission
C2349288|ICD9CM|AB|206.10|Ch mono leu wo achv rmsn
C2349289|ICD9CM|PT|206.12|Chronic monocytic leukemia, in relapse
C2349289|ICD9CM|AB|206.12|Chr mono leuk in relapse
C2349290|ICD9CM|PT|206.20|Subacute monocytic leukemia, without mention of having achieved remission
C2349290|ICD9CM|AB|206.20|Sbac mno leu wo ach rmsn
C2349291|ICD9CM|PT|206.22|Subacute monocytic leukemia, in relapse
C2349291|ICD9CM|AB|206.22|Sbac mono leu in relapse
C2349292|ICD9CM|PT|206.80|Other monocytic leukemia, without mention of having achieved remission
C2349292|ICD9CM|AB|206.80|Ot mono leu wo achv rmsn
C2349293|ICD9CM|PT|206.82|Other monocytic leukemia, in relapse
C2349293|ICD9CM|AB|206.82|Oth mono leuk in relapse
C2349294|ICD9CM|PT|206.90|Unspecified monocytic leukemia, without mention of having achieved remission
C2349294|ICD9CM|AB|206.90|Uns mno leu wo ach rmsn
C2349295|ICD9CM|PT|206.92|Unspecified monocytic leukemia, in relapse
C2349295|ICD9CM|AB|206.92|Mono leuk NOS relapse
C2349296|ICD9CM|PT|207.00|Acute erythremia and erythroleukemia, without mention of having achieved remission
C2349296|ICD9CM|AB|207.00|Ac erth/erlk wo ach rmsn
C2349297|ICD9CM|PT|207.02|Acute erythremia and erythroleukemia, in relapse
C2349297|ICD9CM|AB|207.02|Ac erth/erylk in relapse
C2349298|ICD9CM|PT|207.10|Chronic erythremia, without mention of having achieved remission
C2349298|ICD9CM|AB|207.10|Chr erythrm w/o ach rmsn
C2349299|ICD9CM|PT|207.12|Chronic erythremia, in relapse
C2349299|ICD9CM|AB|207.12|Chr erythrmia in relapse
C2349300|ICD9CM|PT|207.20|Megakaryocytic leukemia, without mention of having achieved remission
C2349300|ICD9CM|AB|207.20|Mgkrcyt leuk wo ach rmsn
C2349301|ICD9CM|PT|207.22|Megakaryocytic leukemia, in relapse
C2349301|ICD9CM|AB|207.22|Mgkrycyt leuk in relapse
C2349302|ICD9CM|PT|207.80|Other specified leukemia, without mention of having achieved remission
C2349302|ICD9CM|AB|207.80|Oth leuk w/o achv rmsn
C2349303|ICD9CM|PT|207.82|Other specified leukemia, in relapse
C2349303|ICD9CM|AB|207.82|Oth spf leuk in relapse
C2349304|ICD9CM|PT|208.00|Acute leukemia of unspecified cell type, without mention of having achieved remission
C2349304|ICD9CM|AB|208.00|Ac leu un cl wo ach rmsn
C2349305|ICD9CM|PT|208.02|Acute leukemia of unspecified cell type, in relapse
C2349305|ICD9CM|AB|208.02|Ac leuk uns cl relapse
C2349306|ICD9CM|PT|208.10|Chronic leukemia of unspecified cell type, without mention of having achieved remission
C2349306|ICD9CM|AB|208.10|Ch leu un cl wo ach rmsn
C2349307|ICD9CM|PT|208.12|Chronic leukemia of unspecified cell type, in relapse
C2349307|ICD9CM|AB|208.12|Ch leu uns cl in relapse
C2349308|ICD9CM|PT|208.20|Subacute leukemia of unspecified cell type, without mention of having achieved remission
C2349308|ICD9CM|AB|208.20|Sbc leu un cl wo ah rmsn
C2349309|ICD9CM|PT|208.22|Subacute leukemia of unspecified cell type, in relapse
C2349309|ICD9CM|AB|208.22|Sbac leu uns cl-relapse
C2349310|ICD9CM|PT|208.80|Other leukemia of unspecified cell type, without mention of having achieved remission
C2349310|ICD9CM|AB|208.80|Ot leu un cl wo ach rmsn
C2349311|ICD9CM|PT|208.82|Other leukemia of unspecified cell type, in relapse
C2349311|ICD9CM|AB|208.82|Oth leuk uns cl-relapse
C2349312|ICD9CM|PT|208.90|Unspecified leukemia, without mention of having achieved remission
C2349312|ICD9CM|AB|208.90|Leuk NOS w/o achv rmsn
C2349313|ICD9CM|PT|209.00|Malignant carcinoid tumor of the small intestine, unspecified portion
C2349313|ICD9CM|AB|209.00|Mal crcnoid sm intst NOS
C2349314|ICD9CM|PT|209.01|Malignant carcinoid tumor of the duodenum
C2349314|ICD9CM|AB|209.01|Malig carcinoid duodenum
C2349315|ICD9CM|PT|209.02|Malignant carcinoid tumor of the jejunum
C2349315|ICD9CM|AB|209.02|Malig carcinoid jejunum
C2349316|ICD9CM|PT|209.03|Malignant carcinoid tumor of the ileum
C2349316|ICD9CM|AB|209.03|Malig carcinoid ileum
C2349317|ICD9CM|PT|209.10|Malignant carcinoid tumor of the large intestine, unspecified portion
C2349317|ICD9CM|AB|209.10|Mal crcnoid lg intst NOS
C2349319|ICD9CM|PT|209.12|Malignant carcinoid tumor of the cecum
C2349319|ICD9CM|AB|209.12|Malig carcinoid cecum
C2349320|ICD9CM|PT|209.13|Malignant carcinoid tumor of the ascending colon
C2349320|ICD9CM|AB|209.13|Mal crcnoid ascend colon
C2349321|ICD9CM|PT|209.14|Malignant carcinoid tumor of the transverse colon
C2349321|ICD9CM|AB|209.14|Mal crcnoid transv colon
C2349322|ICD9CM|PT|209.15|Malignant carcinoid tumor of the descending colon
C2349322|ICD9CM|AB|209.15|Mal carcinoid desc colon
C2349323|ICD9CM|PT|209.16|Malignant carcinoid tumor of the sigmoid colon
C2349323|ICD9CM|AB|209.16|Mal carcinoid sig colon
C2349324|ICD9CM|HT|209.1|Malignant carcinoid tumors of the appendix, large intestine, and rectum
C2349325|ICD9CM|PT|209.20|Malignant carcinoid tumor of unknown primary site
C2349325|ICD9CM|AB|209.20|Mal crcnd prim site unkn
C2349326|ICD9CM|PT|209.21|Malignant carcinoid tumor of the bronchus and lung
C2349326|ICD9CM|AB|209.21|Mal carcinoid bronc/lung
C2349327|ICD9CM|PT|209.24|Malignant carcinoid tumor of the kidney
C2349327|ICD9CM|AB|209.24|Malig carcinoid kidney
C2349328|ICD9CM|PT|209.25|Malignant carcinoid tumor of foregut, not otherwise specified
C2349328|ICD9CM|AB|209.25|Mal carcnoid foregut NOS
C2349329|ICD9CM|PT|209.26|Malignant carcinoid tumor of midgut, not otherwise specified
C2349329|ICD9CM|AB|209.26|Mal carcinoid midgut NOS
C2349330|ICD9CM|PT|209.27|Malignant carcinoid tumor of hindgut, not otherwise specified
C2349330|ICD9CM|AB|209.27|Mal carcnoid hindgut NOS
C2349331|ICD9CM|PT|209.29|Malignant carcinoid tumor of other sites
C2349331|ICD9CM|AB|209.29|Malig carcinoid oth site
C2349332|ICD9CM|HT|209.2|Malignant carcinoid tumors of other and unspecified sites
C2349333|ICD9CM|PT|209.30|Malignant poorly differentiated neuroendocrine carcinoma, any site
C2349333|ICD9CM|AB|209.30|Malig neuroendo ca NOS
C2349335|ICD9CM|HT|209.3|Malignant poorly differentiated neuroendocrine tumors
C2349336|ICD9CM|PT|209.40|Benign carcinoid tumor of the small intestine, unspecified portion
C2349336|ICD9CM|AB|209.40|Ben crcnoid sm intst NOS
C2349337|ICD9CM|PT|209.41|Benign carcinoid tumor of the duodenum
C2349337|ICD9CM|AB|209.41|Ben carcinoid duodenum
C2349338|ICD9CM|PT|209.42|Benign carcinoid tumor of the jejunum
C2349338|ICD9CM|AB|209.42|Benign carcinoid jejunum
C2349339|ICD9CM|PT|209.43|Benign carcinoid tumor of the ileum
C2349339|ICD9CM|AB|209.43|Benign carcinoid ileum
C2349340|ICD9CM|HT|209.4|Benign carcinoid tumors of the small intestine
C2349341|ICD9CM|PT|209.50|Benign carcinoid tumor of the large intestine, unspecified portion
C2349341|ICD9CM|AB|209.50|Ben crcnoid lg intst NOS
C2349342|ICD9CM|PT|209.51|Benign carcinoid tumor of the appendix
C2349342|ICD9CM|AB|209.51|Ben carcinoid appendix
C2349343|ICD9CM|PT|209.52|Benign carcinoid tumor of the cecum
C2349343|ICD9CM|AB|209.52|Benign carcinoid cecum
C2349344|ICD9CM|PT|209.53|Benign carcinoid tumor of the ascending colon
C2349344|ICD9CM|AB|209.53|Ben carcinoid asc colon
C2349345|ICD9CM|PT|209.54|Benign carcinoid tumor of the transverse colon
C2349345|ICD9CM|AB|209.54|Ben crcinoid trans colon
C2349346|ICD9CM|PT|209.55|Benign carcinoid tumor of the descending colon
C2349346|ICD9CM|AB|209.55|Ben carcinoid desc colon
C2349347|ICD9CM|PT|209.56|Benign carcinoid tumor of the sigmoid colon
C2349347|ICD9CM|AB|209.56|Ben carcinoid sig colon
C2349348|ICD9CM|PT|209.57|Benign carcinoid tumor of the rectum
C2349348|ICD9CM|AB|209.57|Benign carcinoid rectum
C2349349|ICD9CM|HT|209.5|Benign carcinoid tumors of the appendix, large intestine, and rectum
C2349350|ICD9CM|PT|209.60|Benign carcinoid tumor of unknown primary site
C2349350|ICD9CM|AB|209.60|Ben crcnd prim site unkn
C2349351|ICD9CM|PT|209.61|Benign carcinoid tumor of the bronchus and lung
C2349351|ICD9CM|AB|209.61|Ben carcinoid bronc/lung
C2349352|ICD9CM|PT|209.62|Benign carcinoid tumor of the thymus
C2349352|ICD9CM|AB|209.62|Benign carcinoid thymus
C2349353|ICD9CM|PT|209.63|Benign carcinoid tumor of the stomach
C2349353|ICD9CM|AB|209.63|Benign carcinoid stomach
C2349354|ICD9CM|PT|209.64|Benign carcinoid tumor of the kidney
C2349354|ICD9CM|AB|209.64|Benign carcinoid kidney
C2349355|ICD9CM|PT|209.65|Benign carcinoid tumor of foregut, not otherwise specified
C2349355|ICD9CM|AB|209.65|Ben crcinoid foregut NOS
C2349356|ICD9CM|PT|209.66|Benign carcinoid tumor of midgut, not otherwise specified
C2349356|ICD9CM|AB|209.66|Ben crcinoid midgut NOS
C2349357|ICD9CM|PT|209.67|Benign carcinoid tumor of hindgut, not otherwise specified
C2349357|ICD9CM|AB|209.67|Ben crcnoid hindgut NOS
C2349358|ICD9CM|PT|209.69|Benign carcinoid tumor of other sites
C2349358|ICD9CM|AB|209.69|Bengn carcinoid oth site
C2349359|ICD9CM|HT|209.6|Benign carcinoid tumors of other and unspecified sites
C2349361|ICD9CM|PT|249.00|Secondary diabetes mellitus without mention of complication, not stated as uncontrolled, or unspecified
C2349361|ICD9CM|AB|249.00|Sec DM wo cmp nt st uncn
C2349362|ICD9CM|PT|249.01|Secondary diabetes mellitus without mention of complication, uncontrolled
C2349362|ICD9CM|AB|249.01|Sec DM wo comp uncontrld
C2349363|ICD9CM|HT|249.0|Secondary diabetes mellitus, without mention of complication
C2349365|ICD9CM|PT|249.10|Secondary diabetes mellitus with ketoacidosis, not stated as uncontrolled, or unspecified
C2349365|ICD9CM|AB|249.10|Sec DM keto nt st uncntr
C2349366|ICD9CM|PT|249.11|Secondary diabetes mellitus with ketoacidosis, uncontrolled
C2349366|ICD9CM|AB|249.11|Sec DM ketoacd uncntrld
C2349367|ICD9CM|HT|249.1|Secondary diabetes mellitus with ketoacidosis
C2349370|ICD9CM|PT|249.20|Secondary diabetes mellitus with hyperosmolarity, not stated as uncontrolled, or unspecified
C2349370|ICD9CM|AB|249.20|Sec DM hpros nt st uncnr
C2349371|ICD9CM|PT|249.21|Secondary diabetes mellitus with hyperosmolarity, uncontrolled
C2349371|ICD9CM|AB|249.21|Sec DM hprosmlr uncntrld
C2349372|ICD9CM|HT|249.2|Secondary diabetes mellitus with hyperosmolarity
C2349374|ICD9CM|PT|249.30|Secondary diabetes mellitus with other coma, not stated as uncontrolled, or unspecified
C2349374|ICD9CM|AB|249.30|Sec DM ot cma nt st uncn
C2349375|ICD9CM|PT|249.31|Secondary diabetes mellitus with other coma, uncontrolled
C2349375|ICD9CM|AB|249.31|Sec DM oth coma uncntrld
C2349376|ICD9CM|HT|249.3|Secondary diabetes mellitus with other coma
C2349380|ICD9CM|PT|249.40|Secondary diabetes mellitus with renal manifestations, not stated as uncontrolled, or unspecified
C2349380|ICD9CM|AB|249.40|Sec DM renl nt st uncntr
C2349381|ICD9CM|PT|249.41|Secondary diabetes mellitus with renal manifestations, uncontrolled
C2349381|ICD9CM|AB|249.41|Sec DM renal uncontrld
C2349382|ICD9CM|HT|249.4|Secondary diabetes mellitus with renal manifestations
C2349383|ICD9CM|PT|249.50|Secondary diabetes mellitus with ophthalmic manifestations, not stated as uncontrolled, or unspecified
C2349383|ICD9CM|AB|249.50|Sec DM ophth nt st uncn
C2349384|ICD9CM|PT|249.51|Secondary diabetes mellitus with ophthalmic manifestations, uncontrolled
C2349384|ICD9CM|AB|249.51|Sec DM ophth uncontrld
C2349385|ICD9CM|HT|249.5|Secondary diabetes mellitus with ophthalmic manifestations
C2349386|ICD9CM|PT|249.60|Secondary diabetes mellitus with neurological manifestations, not stated as uncontrolled, or unspecified
C2349386|ICD9CM|AB|249.60|Sec DM neuro nt st uncn
C2349387|ICD9CM|PT|249.61|Secondary diabetes mellitus with neurological manifestations, uncontrolled
C2349387|ICD9CM|AB|249.61|Sec DM neuro uncontrld
C2349388|ICD9CM|HT|249.6|Secondary diabetes mellitus with neurological manifestations
C2349389|ICD9CM|PT|249.70|Secondary diabetes mellitus with peripheral circulatory disorders, not stated as uncontrolled, or unspecified
C2349389|ICD9CM|AB|249.70|Sec DM circ nt st uncntr
C2349390|ICD9CM|PT|249.71|Secondary diabetes mellitus with peripheral circulatory disorders, uncontrolled
C2349390|ICD9CM|AB|249.71|Sec DM circ uncontrld
C2349391|ICD9CM|HT|249.7|Secondary diabetes mellitus with peripheral circulatory disorders
C2349392|ICD9CM|PT|249.80|Secondary diabetes mellitus with other specified manifestations, not stated as uncontrolled, or unspecified
C2349392|ICD9CM|AB|249.80|Sec DM oth nt st uncontr
C2349393|ICD9CM|PT|249.81|Secondary diabetes mellitus with other specified manifestations, uncontrolled
C2349393|ICD9CM|AB|249.81|Sec DM other uncontrld
C2349394|ICD9CM|HT|249.8|Secondary diabetes mellitus with other specified manifestations
C2349397|ICD9CM|PT|249.90|Secondary diabetes mellitus with unspecified complication, not stated as uncontrolled, or unspecified
C2349397|ICD9CM|AB|249.90|Sec DM unsp nt st uncon
C2349398|ICD9CM|PT|249.91|Secondary diabetes mellitus with unspecified complication, uncontrolled
C2349398|ICD9CM|AB|249.91|Sec DM unsp uncontrold
C2349399|ICD9CM|HT|249.9|Secondary diabetes mellitus with unspecified complication
C2349400|ICD9CM|PT|259.50|Androgen insensitivity, unspecified
C2349400|ICD9CM|AB|259.50|Androgen insensitvty NOS
C2349403|ICD9CM|PT|279.53|Acute on chronic graft-versus-host disease
C2349403|ICD9CM|AB|279.53|Ac on chrn grft-vs-host
C2349407|ICD9CM|PT|33.72|Endoscopic pulmonary airway flow measurement
C2349407|ICD9CM|AB|33.72|Endo pulm arwy flow msmt
C2349409|ICD9CM|HT|33.7|Other endoscopic procedures in bronchus or lung
C2349410|ICD9CM|PT|337.00|Idiopathic peripheral autonomic neuropathy, unspecified
C2349410|ICD9CM|AB|337.00|Idio perph auto neur NOS
C2349411|ICD9CM|PT|337.09|Other idiopathic peripheral autonomic neuropathy
C2349411|ICD9CM|AB|337.09|Idio perph auto neur NEC
C2349417|ICD9CM|PT|339.05|Short lasting unilateral neuralgiform headache with conjunctival injection and tearing
C2349417|ICD9CM|AB|339.05|Shrt lst uni nral hdache
C2349418|ICD9CM|PT|339.09|Other trigeminal autonomic cephalgias
C2349418|ICD9CM|AB|339.09|Trigem autonmc cephl NEC
C2349419|ICD9CM|HT|339.0|Cluster headaches and other trigeminal autonomic cephalgias
C2349421|ICD9CM|PT|339.21|Acute post-traumatic headache
C2349421|ICD9CM|AB|339.21|Ac post-trauma headache
C2349422|MTH|PN|NOCODE|Drug induced headache, NEC in ICD9CM
C2349422|ICD9CM|PT|339.3|Drug induced headache, not elsewhere classified
C2349422|ICD9CM|AB|339.3|Drug induce headache NEC
C2349425|ICD9CM|PT|339.41|Hemicrania continua
C2349425|ICD9CM|AB|339.41|Hemicrania continua
C2349426|ICD9CM|PT|339.42|New daily persistent headache
C2349426|ICD9CM|AB|339.42|New daily pers headache
C2349427|ICD9CM|PT|339.44|Other complicated headache syndrome
C2349427|ICD9CM|AB|339.44|Comp headache synd NEC
C2349428|ICD9CM|HT|339.4|Complicated headache syndromes
C2349432|ICD9CM|PT|346.00|Migraine with aura, without mention of intractable migraine without mention of status migrainosus
C2349432|ICD9CM|AB|346.00|Mgrn w aura wo ntrc mgrn
C2349433|ICD9CM|PT|346.01|Migraine with aura, with intractable migraine, so stated, without mention of status migrainosus
C2349433|ICD9CM|AB|346.01|Mgrn w aura w ntrc mgrn
C2349434|ICD9CM|PT|346.02|Migraine with aura, without mention of intractable migraine with status migrainosus
C2349434|ICD9CM|AB|346.02|Mgrn w aur wo ntrc mgrn
C2349435|ICD9CM|PT|346.03|Migraine with aura, with intractable migraine, so stated, with status migrainosus
C2349435|ICD9CM|AB|346.03|Mgrn w aura w ntrc mgrn
C2349438|ICD9CM|PT|346.10|Migraine without aura, without mention of intractable migraine without mention of status migrainosus
C2349438|ICD9CM|AB|346.10|Mgrn wo aura wo ntrc mgr
C2349439|ICD9CM|PT|346.11|Migraine without aura, with intractable migraine, so stated, without mention of status migrainosus
C2349439|ICD9CM|AB|346.11|Mgrn wo aura w ntrc mgrn
C2349440|ICD9CM|PT|346.12|Migraine without aura, without mention of intractable migraine with status migrainosus
C2349440|ICD9CM|AB|346.12|Mgrn wo aura wo ntrc mgr
C2349441|ICD9CM|PT|346.13|Migraine without aura, with intractable migraine, so stated, with status migrainosus
C2349441|ICD9CM|AB|346.13|Mgrn wo aura w ntrc mgrn
C2349442|ICD9CM|PT|346.20|Variants of migraine, not elsewhere classified, without mention of intractable migraine without mention of status migrainosus
C2349442|ICD9CM|AB|346.20|Vrnt mgrn wo ntr mgr NEC
C2349443|ICD9CM|PT|346.21|Variants of migraine, not elsewhere classified, with intractable migraine, so stated, without mention of status migrainosus
C2349443|ICD9CM|AB|346.21|Vrnt mgrn w ntrc mgr NEC
C2349444|ICD9CM|PT|346.22|Variants of migraine, not elsewhere classified, without mention of intractable migraine with status migrainosus
C2349444|ICD9CM|AB|346.22|Var mgr NEC wo ntc mgr
C2349445|ICD9CM|PT|346.23|Variants of migraine, not elsewhere classified, with intractable migraine, so stated, with status migrainosus
C2349445|ICD9CM|AB|346.23|Var mgrn NEC w ntrc mgr
C2349446|ICD9CM|HT|346.2|Variants of migraine, not elsewhere classified
C2349449|ICD9CM|PT|346.30|Hemiplegic migraine, without mention of intractable migraine without mention of status migrainosus
C2349449|ICD9CM|AB|346.30|Hmplg mgr wo ntrc wo st
C2349450|ICD9CM|PT|346.31|Hemiplegic migraine, with intractable migraine, so stated, without mention of status migrainosus
C2349450|ICD9CM|AB|346.31|Hmplg mgrn w ntrc wo st
C2349451|ICD9CM|PT|346.32|Hemiplegic migraine, without mention of intractable migraine with status migrainosus
C2349451|ICD9CM|AB|346.32|Hemplg mgr wo ntrc w st
C2349452|ICD9CM|PT|346.33|Hemiplegic migraine, with intractable migraine, so stated, with status migrainosus
C2349452|ICD9CM|AB|346.33|Hmplg mgrn w ntrc w st
C2349455|ICD9CM|PT|346.40|Menstrual migraine, without mention of intractable migraine without mention of status migrainosus
C2349455|ICD9CM|AB|346.40|Menst mgr wo ntrc wo st
C2349456|ICD9CM|PT|346.41|Menstrual migraine, with intractable migraine, so stated, without mention of status migrainosus
C2349456|ICD9CM|AB|346.41|Menstl mgrn w ntrc wo st
C2349457|ICD9CM|PT|346.42|Menstrual migraine, without mention of intractable migraine with status migrainosus
C2349457|ICD9CM|AB|346.42|Menstl mgr wo ntrc w st
C2349458|ICD9CM|PT|346.43|Menstrual migraine, with intractable migraine, so stated, with status migrainosus
C2349458|ICD9CM|AB|346.43|Menstl mgrn w ntrc w st
C2349461|ICD9CM|PT|346.50|Persistent migraine aura without cerebral infarction, without mention of intractable migraine without mention of status migrainosus
C2349461|ICD9CM|AB|346.50|Prst aura wo inf/ntr/st
C2349462|ICD9CM|PT|346.51|Persistent migraine aura without cerebral infarction, with intractable migraine, so stated, without mention of status migrainosus
C2349462|ICD9CM|AB|346.51|Prs ara w ntr wo inf/st
C2349463|ICD9CM|PT|346.52|Persistent migraine aura without cerebral infarction, without mention of intractable migraine with status migrainosus
C2349463|ICD9CM|AB|346.52|Prs ara wo inf/ntr w st
C2349464|ICD9CM|PT|346.53|Persistent migraine aura without cerebral infarction, with intractable migraine, so stated, with status migrainosus
C2349464|ICD9CM|AB|346.53|Prs ara wo inf w ntr/st
C2349465|ICD9CM|HT|346.5|Persistent migraine aura without cerebral infarction
C2349467|ICD9CM|PT|346.60|Persistent migraine aura with cerebral infarction, without mention of intractable migraine without mention of status migrainosus
C2349467|ICD9CM|AB|346.60|Prs ara w inf wo ntr/st
C2349468|ICD9CM|PT|346.61|Persistent migraine aura with cerebral infarction, with intractable migraine, so stated, without mention of status migrainosus
C2349468|ICD9CM|AB|346.61|Prs ara w/inf/ntr wo st
C2349469|ICD9CM|PT|346.62|Persistent migraine aura with cerebral infarction, without mention of intractable migraine with status migrainosus
C2349469|ICD9CM|AB|346.62|Prs ara wo ntr w inf/st
C2349470|ICD9CM|PT|346.63|Persistent migraine aura with cerebral infarction, with intractable migraine, so stated, with status migrainosus
C2349470|ICD9CM|AB|346.63|Prst ara w inf w ntr/st
C2349471|ICD9CM|HT|346.6|Persistent migraine aura with cerebral infarction
C2349472|ICD9CM|PT|346.70|Chronic migraine without aura, without mention of intractable migraine without mention of status migrainosus
C2349472|ICD9CM|AB|346.70|Ch mgr wo ar wo nt wo st
C2349473|ICD9CM|PT|346.71|Chronic migraine without aura, with intractable migraine, so stated, without mention of status migrainosus
C2349473|ICD9CM|AB|346.71|Ch mgr wo ara w nt wo st
C2349474|ICD9CM|PT|346.72|Chronic migraine without aura, without mention of intractable migraine with status migrainosus
C2349474|ICD9CM|AB|346.72|Ch mgr wo ara wo nt w st
C2349475|ICD9CM|PT|346.73|Chronic migraine without aura, with intractable migraine, so stated, with status migrainosus
C2349475|ICD9CM|AB|346.73|Ch mgr wo ara w ntr w st
C2349476|ICD9CM|HT|346.7|Chronic migraine without aura
C2349478|ICD9CM|PT|346.81|Other forms of migraine, with intractable migraine, so stated, without mention of status migrainosus
C2349478|ICD9CM|AB|346.81|Othr migrne w ntrc mgrne
C2349479|ICD9CM|PT|346.82|Other forms of migraine, without mention of intractable migraine with status migrainosus
C2349479|ICD9CM|AB|346.82|Oth mgr wo ntrc w st mgr
C2349480|ICD9CM|PT|346.83|Other forms of migraine, with intractable migraine, so stated, with status migrainosus
C2349480|ICD9CM|AB|346.83|Oth mgr w ntrc w st mgr
C2349481|ICD9CM|PT|346.92|Migraine, unspecified, without mention of intractable migraine with status migrainosus
C2349481|ICD9CM|AB|346.92|Mgr NOS wo ntrc w st mgr
C2349482|ICD9CM|PT|346.93|Migraine, unspecified, with intractable migraine, so stated, with status migrainosus
C2349482|ICD9CM|AB|346.93|Mgrn NOS w ntrc w st mgr
C2349483|ICD9CM|PT|349.31|Accidental puncture or laceration of dura during a procedure
C2349483|ICD9CM|AB|349.31|Accid punc/op lac dura
C2349485|ICD9CM|PT|349.39|Other dural tear
C2349485|ICD9CM|AB|349.39|Dural tear NEC
C2349494|ICD9CM|PT|37.36|Excision, destruction, or exclusion of left atrial appendage (LAA)
C2349494|ICD9CM|AB|37.36|Exc,destrct,exclus LAA
C2349495|ICD9CM|PT|37.52|Implantation of total internal biventricular heart replacement system
C2349495|ICD9CM|AB|37.52|Imp tot int bi ht rp sys
C2349496|ICD9CM|PT|37.55|Removal of internal biventricular heart replacement system
C2349496|ICD9CM|AB|37.55|Rem int bivent hrt sys
C2349498|ICD9CM|PT|37.60|Implantation or insertion of biventricular external heart assist system
C2349498|ICD9CM|AB|37.60|Imp bivn ext hrt ast sys
C2349500|ICD9CM|PT|37.62|Insertion of temporary non-implantable extracorporeal circulatory assist device
C2349500|ICD9CM|AB|37.62|Insrt non-impl circ dev
C2349503|ICD9CM|PT|37.64|Removal of external heart assist system(s) or device(s)
C2349503|ICD9CM|AB|37.64|Remve ext hrt assist sys
C2349506|ICD9CM|PT|37.65|Implant of single ventricular (extracorporeal) external heart assist system
C2349506|ICD9CM|AB|37.65|Imp vent ext hrt ast sys
C2349508|ICD9CM|PT|38.23|Intravascular spectroscopy
C2349508|ICD9CM|AB|38.23|Intravasclr spectroscopy
C2349509|ICD9CM|PT|414.3|Coronary atherosclerosis due to lipid rich plaque
C2349509|ICD9CM|AB|414.3|Cor ath d/t lpd rch plaq
C2349510|ICD9CM|PT|45.71|Open and other multiple segmental resection of large intestine
C2349510|ICD9CM|AB|45.71|Opn mul seg lg intes NEC
C2349511|ICD9CM|PT|45.72|Open and other cecectomy
C2349511|ICD9CM|AB|45.72|Open cecectomy NEC
C2349512|ICD9CM|PT|45.73|Open and other right hemicolectomy
C2349512|ICD9CM|AB|45.73|Opn rt hemicolectomy NEC
C2349513|ICD9CM|PT|45.74|Open and other resection of transverse colon
C2349513|ICD9CM|AB|45.74|Opn transv colon res NEC
C2349514|ICD9CM|PT|45.75|Open and other left hemicolectomy
C2349514|ICD9CM|AB|45.75|Opn lft hemicolectmy NEC
C2349515|ICD9CM|PT|45.76|Open and other sigmoidectomy
C2349515|ICD9CM|AB|45.76|Open sigmoidectomy NEC
C2349516|ICD9CM|PT|45.79|Other and unspecified partial excision of large intestine
C2349516|ICD9CM|AB|45.79|Prt lg intes exc NEC/NOS
C2349517|ICD9CM|HT|45.7|Open and other partial excision of large intestine
C2349518|ICD9CM|PT|45.81|Laparoscopic total intra-abdominal colectomy
C2349518|ICD9CM|AB|45.81|Lap tot intr-ab colectmy
C2349519|ICD9CM|PT|45.82|Open total intra-abdominal colectomy
C2349519|ICD9CM|AB|45.82|Op tot intr-abd colectmy
C2349520|ICD9CM|PT|45.83|Other and unspecified total intra-abdominal colectomy
C2349520|ICD9CM|AB|45.83|Tot abd colectmy NEC/NOS
C2349522|ICD9CM|PT|48.40|Pull-through resection of rectum, not otherwise specified
C2349522|ICD9CM|AB|48.40|Pull-thru res rectum NOS
C2349523|ICD9CM|PT|48.42|Laparoscopic pull-through resection of rectum
C2349523|ICD9CM|AB|48.42|Lap pull-thru res rectum
C2349524|ICD9CM|PT|48.43|Open pull-through resection of rectum
C2349524|ICD9CM|AB|48.43|Opn pull-thru res rectum
C2349525|ICD9CM|PT|48.50|Abdominoperineal resection of the rectum, not otherwise specified
C2349525|ICD9CM|AB|48.50|Abdperneal res rectm NOS
C2349526|ICD9CM|PT|48.51|Laparoscopic abdominoperineal resection of the rectum
C2349526|ICD9CM|AB|48.51|Lap abdperneal resc rec
C2349527|ICD9CM|PT|48.52|Open abdominoperineal resection of the rectum
C2349527|ICD9CM|AB|48.52|Opn abdperneal resc rec
C2349528|ICD9CM|PT|48.59|Other abdominoperineal resection of the rectum
C2349528|ICD9CM|AB|48.59|Abdperneal resc rect NEC
C2349529|ICD9CM|PT|482.41|Methicillin susceptible pneumonia due to Staphylococcus aureus
C2349529|ICD9CM|AB|482.41|Meth sus pneum d/t Staph
C2349532|ICD9CM|PT|511.89|Other specified forms of effusion, except tuberculous
C2349532|ICD9CM|AB|511.89|Effusion NEC exc tb
C2349539|ICD9CM|PT|53.01|Other and open repair of direct inguinal hernia
C2349539|ICD9CM|AB|53.01|Opn rep dir ing hern NEC
C2349541|ICD9CM|PT|53.02|Other and open repair of indirect inguinal hernia
C2349541|ICD9CM|AB|53.02|Opn rep ind ing hern NEC
C2349542|ICD9CM|PT|53.03|Other and open repair of direct inguinal hernia with graft or prosthesis
C2349542|ICD9CM|AB|53.03|Opn dir ing hern-gft NEC
C2349543|ICD9CM|PT|53.04|Other and open repair of indirect inguinal hernia with graft or prosthesis
C2349543|ICD9CM|AB|53.04|Opn ind ing hern-gft NEC
C2349544|ICD9CM|HT|53.0|Other unilateral repair of inguinal hernia
C2349545|ICD9CM|PT|53.11|Other and open bilateral repair of direct inguinal hernia
C2349545|ICD9CM|AB|53.11|Opn bil dir ing hern NEC
C2349546|ICD9CM|PT|53.12|Other and open bilateral repair of indirect inguinal hernia
C2349546|ICD9CM|AB|53.12|Opn bil ind ing hern NEC
C2349547|ICD9CM|PT|53.13|Other and open bilateral repair of inguinal hernia, one direct and one indirect
C2349547|ICD9CM|AB|53.13|Opn bi dr/in ing hrn NEC
C2349548|ICD9CM|PT|53.14|Other and open bilateral repair of direct inguinal hernia with graft or prosthesis
C2349548|ICD9CM|AB|53.14|Opn bi dr ing hrn-gr NEC
C2349549|ICD9CM|PT|53.15|Other and open bilateral repair of indirect inguinal hernia with graft or prosthesis
C2349549|ICD9CM|AB|53.15|Op bi in ing hrn-grf NEC
C2349550|ICD9CM|PT|53.16|Other and open bilateral repair of inguinal hernia, one direct and one indirect, with graft or prosthesis
C2349550|ICD9CM|AB|53.16|Op bi dr/in ig hr-gr NEC
C2349551|ICD9CM|HT|53.1|Other bilateral repair of inguinal hernia
C2349552|ICD9CM|PT|53.41|Other and open repair of umbilical hernia with graft or prosthesis
C2349552|ICD9CM|AB|53.41|Opn rep umb hrn-grft NEC
C2349553|ICD9CM|PT|53.42|Laparoscopic repair of umbilical hernia with graft or prosthesis
C2349553|ICD9CM|AB|53.42|Lap umbil hernia-graft
C2349554|ICD9CM|PT|53.43|Other laparoscopic umbilical herniorrhaphy
C2349554|ICD9CM|AB|53.43|Lap umbilical hernia NEC
C2349555|ICD9CM|PT|53.49|Other open umbilical herniorrhaphy
C2349555|ICD9CM|AB|53.49|Open rep umbil hern NEC
C2349556|ICD9CM|PT|53.61|Other open incisional hernia repair with graft or prosthesis
C2349556|ICD9CM|AB|53.61|Open incis hern-grft NEC
C2349557|ICD9CM|PT|53.62|Laparoscopic incisional hernia repair with graft or prosthesis
C2349557|ICD9CM|AB|53.62|Lap incis hern repr-grft
C2349558|ICD9CM|PT|53.63|Other laparoscopic repair of other hernia of anterior abdominal wall with graft or prosthesis
C2349558|ICD9CM|AB|53.63|Lap hern ant abd-gft NEC
C2349559|ICD9CM|PT|53.69|Other and open repair of other hernia of anterior abdominal wall with graft or prosthesis
C2349559|ICD9CM|AB|53.69|Opn hern ant abd-grf NEC
C2349560|ICD9CM|PT|53.71|Laparoscopic repair of diaphragmatic hernia, abdominal approach
C2349560|ICD9CM|AB|53.71|Lap abd rep-diaphr hern
C2349561|ICD9CM|PT|53.72|Other and open repair of diaphragmatic hernia, abdominal approach
C2349561|ICD9CM|AB|53.72|Opn abd diaphrm hern NEC
C2349562|ICD9CM|PT|53.75|Repair of diaphragmatic hernia, abdominal approach, not otherwise specified
C2349562|ICD9CM|AB|53.75|Abd rep-diaphr hern NOS
C2349563|ICD9CM|PT|53.83|Laparoscopic repair of diaphragmatic hernia, with thoracic approach
C2349563|ICD9CM|AB|53.83|Lap thorc app-diaph hern
C2349564|ICD9CM|PT|53.84|Other and open repair of diaphragmatic hernia, with thoracic approach
C2349564|ICD9CM|AB|53.84|Opn thorc diaph hern NEC
C2349565|ICD9CM|PT|535.70|Eosinophilic gastritis, without mention of hemorrhage
C2349565|ICD9CM|AB|535.70|Eosinophil gastrt wo hem
C2349566|ICD9CM|PT|535.71|Eosinophilic gastritis, with hemorrhage
C2349566|ICD9CM|AB|535.71|Eosinophilc gastrt w hem
C2349567|ICD9CM|HT|558.4|Eosinophilic gastroenteritis and colitis
C2349571|ICD9CM|PT|611.83|Capsular contracture of breast implant
C2349571|ICD9CM|AB|611.83|Capslr contrctr brst imp
C2349574|ICD9CM|PT|612.0|Deformity of reconstructed breast
C2349574|ICD9CM|AB|612.0|Deformity reconst breast
C2349578|ICD9CM|PT|612.1|Disproportion of reconstructed breast
C2349578|ICD9CM|AB|612.1|Disproportn reconst brst
C2349581|ICD9CM|HT|612|Deformity and disproportion of reconstructed breast
C2349583|ICD9CM|PT|625.79|Other vulvodynia
C2349583|ICD9CM|AB|625.79|Other vulvodynia
C2349584|ICD9CM|PT|649.70|Cervical shortening, unspecified as to episode of care or not applicable
C2349584|ICD9CM|AB|649.70|Cervical shortening-unsp
C2349585|ICD9CM|PT|649.71|Cervical shortening, delivered, with or without mention of antepartum condition
C2349585|ICD9CM|AB|649.71|Cervical shortening-del
C2349586|ICD9CM|PT|649.73|Cervical shortening, antepartum condition or complication
C2349586|ICD9CM|AB|649.73|Cervical shortening-ante
C2349587|ICD9CM|HT|649.7|Cervical shortening
C2349589|ICD9CM|HT|656|Other known or suspected fetal and placental problems affecting management of mother
C2349590|ICD9CM|HT|678-679.99|OTHER MATERNAL AND FETAL COMPLICATIONS
C2349591|ICD9CM|PT|678.00|Fetal hematologic conditions, unspecified as to episode of care or not applicable
C2349591|ICD9CM|AB|678.00|Fetal hematologic-unspec
C2349592|ICD9CM|PT|678.01|Fetal hematologic conditions, delivered, with or without mention of antepartum condition
C2349592|ICD9CM|AB|678.01|Fetal hematologic-deliv
C2349593|ICD9CM|PT|678.03|Fetal hematologic conditions, antepartum condition or complication
C2349593|ICD9CM|AB|678.03|Fetal hematologic-ante
C2349594|ICD9CM|HT|678.0|Fetal hematologic conditions
C2349597|ICD9CM|PT|678.10|Fetal conjoined twins, unspecified as to episode of care or not applicable
C2349597|ICD9CM|AB|678.10|Fetal conjoin twins-unsp
C2349598|ICD9CM|PT|678.11|Fetal conjoined twins, delivered, with or without mention of antepartum condition
C2349598|ICD9CM|AB|678.11|Fetal conjoin twins-del
C2349599|ICD9CM|PT|678.13|Fetal conjoined twins, antepartum condition or complication
C2349599|ICD9CM|AB|678.13|Fetal conjoin twins-ante
C2349600|ICD9CM|HT|678.1|Fetal conjoined twins
C2349601|ICD9CM|HT|678|Other fetal conditions
C2349602|ICD9CM|PT|679.00|Maternal complications from in utero procedure, unspecified as to episode of care or not applicable
C2349602|ICD9CM|AB|679.00|Mat comp in utero-unsp
C2349603|ICD9CM|PT|679.01|Maternal complications from in utero procedure, delivered, with or without mention of antepartum condition
C2349603|ICD9CM|AB|679.01|Mat comp in utero-del
C2349604|ICD9CM|PT|679.02|Maternal complications from in utero procedure, delivered, with mention of postpartum complication
C2349604|ICD9CM|AB|679.02|Mat comp in utro-del-p/p
C2349605|ICD9CM|PT|679.03|Maternal complications from in utero procedure, antepartum condition or complication
C2349605|ICD9CM|AB|679.03|Mat comp in utero-ante
C2349606|ICD9CM|PT|679.04|Maternal complications from in utero procedure, postpartum condition or complication
C2349606|ICD9CM|AB|679.04|Mat comp in utero-p/p
C2349607|ICD9CM|HT|679.0|Maternal complications from in utero procedure
C2349608|ICD9CM|PT|679.10|Fetal complications from in utero procedure, unspecified as to episode of care or not applicable
C2349608|ICD9CM|AB|679.10|Fetal comp in utero-unsp
C2349609|ICD9CM|PT|679.11|Fetal complications from in utero procedure, delivered, with or without mention of antepartum condition
C2349609|ICD9CM|AB|679.11|Fetal comp in utero-del
C2349610|ICD9CM|PT|679.12|Fetal complications from in utero procedure, delivered, with mention of postpartum complication
C2349610|ICD9CM|AB|679.12|Ftl cmp in utro-del-p/p
C2349611|ICD9CM|PT|679.13|Fetal complications from in utero procedure, antepartum condition or complication
C2349611|ICD9CM|AB|679.13|Fetal comp in utero-ante
C2349612|ICD9CM|PT|679.14|Fetal complications from in utero procedure, postpartum condition or complication
C2349612|ICD9CM|AB|679.14|Fetal comp in utero-p/p
C2349613|ICD9CM|HT|679.1|Fetal complications from in utero procedure
C2349615|ICD9CM|HT|679|Complications of in utero procedures
C2349616|ICD9CM|PT|695.14|Stevens-Johnson syndrome-toxic epidermal necrolysis overlap syndrome
C2349616|ICD9CM|AB|695.14|Stevens-Johnson-TEN syn
C2349618|ICD9CM|PT|695.50|Exfoliation due to erythematous condition involving less than 10 percent of body surface
C2349618|ICD9CM|AB|695.50|Exfol d/t eryth <10% bdy
C2349620|ICD9CM|PT|695.51|Exfoliation due to erythematous condition involving 10-19 percent of body surface
C2349620|ICD9CM|AB|695.51|Exfl d/t eryth 10-19 bdy
C2349621|ICD9CM|PT|695.52|Exfoliation due to erythematous condition involving 20-29 percent of body surface
C2349621|ICD9CM|AB|695.52|Exfl d/t eryth 20-29 bdy
C2349622|ICD9CM|PT|695.53|Exfoliation due to erythematous condition involving 30-39 percent of body surface
C2349622|ICD9CM|AB|695.53|Exfl d/t eryth 30-39 bdy
C2349623|ICD9CM|PT|695.54|Exfoliation due to erythematous condition involving 40-49 percent of body surface
C2349623|ICD9CM|AB|695.54|Exfl d/t eryth 40-49 bdy
C2349624|ICD9CM|PT|695.55|Exfoliation due to erythematous condition involving 50-59 percent of body surface
C2349624|ICD9CM|AB|695.55|Exfl d/t eryth 50-59 bdy
C2349625|ICD9CM|PT|695.56|Exfoliation due to erythematous condition involving 60-69 percent of body surface
C2349625|ICD9CM|AB|695.56|Exfl d/t eryth 60-69 bdy
C2349626|ICD9CM|PT|695.57|Exfoliation due to erythematous condition involving 70-79 percent of body surface
C2349626|ICD9CM|AB|695.57|Exfl d/t eryth 70-79 bdy
C2349627|ICD9CM|PT|695.58|Exfoliation due to erythematous condition involving 80-89 percent of body surface
C2349627|ICD9CM|AB|695.58|Exfl d/t eryth 80-89 bdy
C2349628|ICD9CM|PT|695.59|Exfoliation due to erythematous condition involving 90 percent or more of body surface
C2349628|ICD9CM|AB|695.59|Exfl d/t eryth >=90% bdy
C2349629|ICD9CM|HT|695.5|Exfoliation due to erythematous conditions according to extent of body surface involved
C2349630|ICD9CM|HT|707.1|Ulcer of lower limbs, except pressure ulcer
C2349631|ICD9CM|PT|707.20|Pressure ulcer, unspecified stage
C2349631|ICD9CM|AB|707.20|Pressure ulcer,stage NOS
C2349647|ICD9CM|AB|729.91|Post-traumatic seroma
C2349647|ICD9CM|PT|729.91|Post-traumatic seroma
C2349648|ICD9CM|PT|729.92|Nontraumatic hematoma of soft tissue
C2349648|ICD9CM|AB|729.92|Nontrauma hema soft tiss
C2349651|ICD9CM|PT|733.96|Stress fracture of femoral neck
C2349651|ICD9CM|AB|733.96|Stress fx femoral neck
C2349653|ICD9CM|PT|733.97|Stress fracture of shaft of femur
C2349653|ICD9CM|AB|733.97|Stress fx shaft femur
C2349657|ICD9CM|PT|760.61|Newborn affected by amniocentesis
C2349657|ICD9CM|AB|760.61|Amniocentesis affect NB
C2349658|ICD9CM|PT|760.62|Newborn affected by other in utero procedure
C2349658|ICD9CM|AB|760.62|In utero proc NEC aff NB
C2349659|ICD9CM|PT|760.63|Newborn affected by other surgical operations on mother during pregnancy
C2349659|ICD9CM|AB|760.63|Mat surg dur preg aff NB
C2349660|ICD9CM|PT|760.64|Newborn affected by previous surgical procedure on mother not associated with pregnancy
C2349660|ICD9CM|AB|760.64|Prev matern surg aff NB
C2349661|ICD9CM|HT|760.6|Surgical operation on mother and fetus
C2349662|ICD9CM|PT|777.50|Necrotizing enterocolitis in newborn, unspecified
C2349662|ICD9CM|AB|777.50|Nec enterocoltis NB NOS
C2349669|ICD9CM|HT|777.5|Necrotizing enterocolitis in newborn
C2349670|ICD9CM|PT|780.61|Fever presenting with conditions classified elsewhere
C2349670|ICD9CM|AB|780.61|Fever in other diseases
C2349671|ICD9CM|PT|780.62|Postprocedural fever
C2349671|ICD9CM|AB|780.62|Postprocedural fever
C2349672|ICD9CM|PT|780.63|Postvaccination fever
C2349672|ICD9CM|AB|780.63|Postvaccination fever
C2349674|ICD9CM|PT|780.64|Chills (without fever)
C2349674|ICD9CM|AB|780.64|Chills (without fever)
C2349675|ICD9CM|HT|780.6|Fever and other physiologic disturbances of temperature regulation
C2349680|ICD9CM|PT|795.07|Satisfactory cervical smear but lacking transformation zone
C2349680|ICD9CM|AB|795.07|Sat cerv smr-no trnsfrm
C2349681|ICD9CM|PT|795.08|Unsatisfactory cervical cytology smear
C2349681|ICD9CM|AB|795.08|Unsat cerv cytlogy smear
C2349683|ICD9CM|PT|795.10|Abnormal glandular Papanicolaou smear of vagina
C2349683|ICD9CM|AB|795.10|Abn gland pap smr vagina
C2349685|ICD9CM|AB|795.11|Pap smear vag w ASC-US
C2349685|ICD9CM|PT|795.11|Papanicolaou smear of vagina with atypical squamous cells of undetermined significance (ASC-US)
C2349686|ICD9CM|AB|795.12|Pap smear vagina w ASC-H
C2349686|ICD9CM|PT|795.12|Papanicolaou smear of vagina with atypical squamous cells cannot exclude high grade squamous intraepithelial lesion (ASC-H)
C2349687|ICD9CM|AB|795.13|Pap smear vagina w LGSIL
C2349687|ICD9CM|PT|795.13|Papanicolaou smear of vagina with low grade squamous intraepithelial lesion (LGSIL)
C2349688|ICD9CM|PT|795.14|Papanicolaou smear of vagina with high grade squamous intraepithelial lesion (HGSIL)
C2349688|ICD9CM|AB|795.14|Pap smear vagina w HGSIL
C2349689|ICD9CM|AB|795.15|Vag hi risk HPV-DNA pos
C2349689|ICD9CM|PT|795.15|Vaginal high risk human papillomavirus (HPV) DNA test positive
C2349690|ICD9CM|AB|795.16|Pap smr vag-cytol malig
C2349690|ICD9CM|PT|795.16|Papanicolaou smear of vagina with cytologic evidence of malignancy
C2349693|ICD9CM|PT|795.19|Other abnormal Papanicolaou smear of vagina and vaginal HPV
C2349693|ICD9CM|AB|795.19|Oth abn Pap smr vag/HPV
C2349696|ICD9CM|HT|795.1|Abnormal Papanicolaou smear of vagina and vaginal HPV
C2349699|ICD9CM|PT|796.70|Abnormal glandular Papanicolaou smear of anus
C2349699|ICD9CM|AB|796.70|Abn gland pap smear anus
C2349701|ICD9CM|PT|796.71|Papanicolaou smear of anus with atypical squamous cells of undetermined significance (ASC-US)
C2349701|ICD9CM|AB|796.71|Pap smear anus w ASC-US
C2349702|ICD9CM|PT|796.72|Papanicolaou smear of anus with atypical squamous cells cannot exclude high grade squamous intraepithelial lesion (ASC-H)
C2349702|ICD9CM|AB|796.72|Pap smear anus w ASC-H
C2349703|ICD9CM|PT|796.73|Papanicolaou smear of anus with low grade squamous intraepithelial lesion (LGSIL)
C2349703|ICD9CM|AB|796.73|Pap smear anus w LGSIL
C2349704|ICD9CM|AB|796.74|Pap smear anus w HGSIL
C2349704|ICD9CM|PT|796.74|Papanicolaou smear of anus with high grade squamous intraepithelial lesion (HGSIL)
C2349705|ICD9CM|AB|796.75|Anal hi risk HPV-DNA pos
C2349705|ICD9CM|PT|796.75|Anal high risk human papillomavirus (HPV) DNA test positive
C2349706|ICD9CM|PT|796.76|Papanicolaou smear of anus with cytologic evidence of malignancy
C2349706|ICD9CM|AB|796.76|Pap smr anus-cytol malig
C2349707|ICD9CM|PT|796.77|Satisfactory anal smear but lacking transformation zone
C2349707|ICD9CM|AB|796.77|Sat anal smr-no trnsfrm
C2349708|ICD9CM|PT|796.78|Unsatisfactory anal cytology smear
C2349708|ICD9CM|AB|796.78|Anal cytolgy smr unsatis
C2349710|ICD9CM|PT|796.79|Other abnormal Papanicolaou smear of anus and anal HPV
C2349710|ICD9CM|AB|796.79|Oth abn Pap smr anus/HPV
C2349713|ICD9CM|HT|796.7|Abnormal cytologic smear of anus and anal HPV
C2349714|ICD9CM|PT|80.53|Repair of the anulus fibrosus with graft or prosthesis
C2349714|ICD9CM|AB|80.53|Rep anulus fibrosus-grft
C2349715|ICD9CM|PT|80.54|Other and unspecified repair of the anulus fibrosus
C2349715|ICD9CM|AB|80.54|Rep anuls fibros NEC/NOS
C2349721|ICD9CM|HT|80.5|Excision, destruction and other repair of intervertebral disc
C2349722|ICD9CM|PT|81.65|Percutaneous vertebroplasty
C2349722|ICD9CM|AB|81.65|Percutan vertebroplasty
C2349727|ICD9CM|PT|85.70|Total reconstruction of breast, not otherwise specified
C2349727|ICD9CM|AB|85.70|Totl reconstc breast NOS
C2349729|ICD9CM|PT|85.72|Transverse rectus abdominis myocutaneous (TRAM) flap, pedicled
C2349729|ICD9CM|AB|85.72|TRAM flap, pedicled
C2349730|ICD9CM|PT|85.73|Transverse rectus abdominis myocutaneous (TRAM) flap, free
C2349730|ICD9CM|AB|85.73|TRAM flap, free
C2349731|ICD9CM|PT|85.74|Deep inferior epigastric artery perforator (DIEP) flap, free
C2349731|ICD9CM|AB|85.74|DIEP flap, free
C2349732|ICD9CM|PT|85.75|Superficial inferior epigastric artery (SIEA) flap, free
C2349732|ICD9CM|AB|85.75|SIEA flap, free
C2349733|ICD9CM|PT|85.76|Gluteal artery perforator (GAP) flap, free
C2349733|ICD9CM|AB|85.76|GAP flap, free
C2349734|ICD9CM|PT|85.79|Other total reconstruction of breast
C2349734|ICD9CM|AB|85.79|Totl reconst breast NEC
C2349736|ICD9CM|PT|038.11|Methicillin susceptible Staphylococcus aureus septicemia
C2349736|ICD9CM|AB|038.11|Meth susc Staph aur sept
C2349738|ICD9CM|PT|041.12|Methicillin resistant Staphylococcus aureus in conditions classified elsewhere and of unspecified site
C2349738|ICD9CM|AB|041.12|MRSA elsewhere/NOS
C2349739|ICD9CM|HT|045-049.99|POLIOMYELITIS AND OTHER NON-ARTHROPOD-BORNE VIRAL DISEASES AND PRION DISEASES OF CENTRAL NERVOUS SYSTEM
C2349740|ICD9CM|PT|93.90|Non-invasive mechanical ventilation
C2349740|ICD9CM|AB|93.90|Non-invasive mech vent
C2349743|ICD9CM|PT|96.70|Continuous invasive mechanical ventilation of unspecified duration
C2349743|ICD9CM|AB|96.70|Con inv mec ven-unsp dur
C2349744|ICD9CM|PT|96.71|Continuous invasive mechanical ventilation for less than 96 consecutive hours
C2349744|ICD9CM|AB|96.71|Cont inv mec ven <96 hrs
C2349745|ICD9CM|PT|96.72|Continuous invasive mechanical ventilation for 96 consecutive hours or more
C2349745|ICD9CM|AB|96.72|Cont inv mec ven 96+ hrs
C2349746|ICD9CM|HT|96.7|Other continuous invasive mechanical ventilation
C2349756|ICD9CM|PT|046.19|Other and unspecified Creutzfeldt-Jakob disease
C2349756|ICD9CM|AB|046.19|Creutzfldt-Jakob NEC/NOS
C2349759|ICD9CM|PT|046.79|Other and unspecified prion disease of central nervous system
C2349759|ICD9CM|AB|046.79|Prion dis of CNS NEC/NOS
C2349760|ICD9CM|HT|046.7|Other specified prion diseases of central nervous system
C2349761|ICD9CM|HT|046|Slow virus infections and prion diseases of central nervous system
C2349762|ICD9CM|HT|051.0|Cowpox and vaccinia not from vaccination
C2349763|ICD9CM|PT|059.00|Orthopoxvirus infection, unspecified
C2349763|ICD9CM|AB|059.00|Orthopoxvirus infect NOS
C2349765|ICD9CM|PT|059.11|Bovine stomatitis
C2349765|ICD9CM|AB|059.11|Bovine stomatitis
C2349769|ICD9CM|PT|997.39|Other respiratory complications
C2349769|ICD9CM|AB|997.39|Respiratory comp NEC
C2349787|ICD9CM|PT|998.33|Disruption of traumatic injury wound repair
C2349787|ICD9CM|AB|998.33|Disrpt trauma wound repr
C2349794|ICD9CM|PT|999.81|Extravasation of vesicant chemotherapy
C2349794|ICD9CM|AB|999.81|Extravstn vesicant chemo
C2349796|ICD9CM|PT|999.82|Extravasation of other vesicant agent
C2349796|ICD9CM|AB|999.82|Extravasn vesicant NEC
C2349798|ICD9CM|PT|999.88|Other infusion reaction
C2349798|ICD9CM|AB|999.88|Infusion reaction NEC
C2349799|MTH|PN|NOCODE|TRANSFUSION REACTION NEC in ICD9CM
C2349799|ICD9CM|PT|999.89|Other transfusion reaction
C2349799|ICD9CM|AB|999.89|Transfusion reaction NEC
C2349800|ICD9CM|HT|999.8|Other infusion and transfusion reaction, not elsewhere classified
C2349803|ICD9CM|PT|E927.0|Overexertion from sudden strenuous movement
C2349803|ICD9CM|AB|E927.0|Overxrt-sudn stren mvmt
C2349805|ICD9CM|PT|E927.1|Overexertion from prolonged static position
C2349805|ICD9CM|AB|E927.1|Overxrt-prolng stc postn
C2349809|ICD9CM|PT|E927.2|Excessive physical exertion
C2349809|ICD9CM|AB|E927.2|Excess physical exert
C2349810|ICD9CM|PT|E927.3|Cumulative trauma from repetitive motion
C2349810|ICD9CM|AB|E927.3|Cumltv trma-repetv motn
C2349812|ICD9CM|PT|E927.4|Cumulative trauma from repetitive impact
C2349812|ICD9CM|AB|E927.4|Cumltv trma-repetv impct
C2349813|ICD9CM|PT|E927.8|Other overexertion and strenuous and repetitive movements or loads
C2349813|ICD9CM|AB|E927.8|Overexert reptv mvmt NEC
C2349814|ICD9CM|PT|E927.9|Unspecified overexertion and strenuous and repetitive movements or loads
C2349814|ICD9CM|AB|E927.9|Overexert reptv mvmt NOS
C2349815|ICD9CM|HT|E927|Overexertion and strenuous and repetitive movements or loads
C2349817|ICD9CM|HT|V01-V91.99|SUPPLEMENTARY CLASSIFICATION OF FACTORS INFLUENCING HEALTH STATUS AND CONTACT WITH HEALTH SERVICES
C2349826|ICD9CM|PT|V07.52|Use of aromatase inhibitors
C2349826|ICD9CM|AB|V07.52|Use aromatase inhibitors
C2349833|ICD9CM|PT|V07.59|Use of other agents affecting estrogen receptors and estrogen levels
C2349833|ICD9CM|AB|V07.59|Use oth agnt af estrogen
C2349852|ICD9CM|PT|V15.51|Personal history of traumatic fracture
C2349852|ICD9CM|AB|V15.51|Hx traumatic fracture
C2349854|ICD9CM|PT|V15.59|Personal history of other injury
C2349854|ICD9CM|AB|V15.59|Hx injury NEC
C2349855|ICD9CM|PT|059.19|Other parapoxvirus infections
C2349855|ICD9CM|HT|059.1|Other parapoxvirus infections
C2349855|ICD9CM|AB|059.19|Parapoxvirus infectn NEC
C2349857|ICD9CM|HT|059.2|Yatapoxvirus infections
C2349857|ICD9CM|AB|059.20|Yatapoxvirus infectn NOS
C2349857|ICD9CM|PT|059.20|Yatapoxvirus infection, unspecified
C2349858|ICD9CM|HT|059|Other poxvirus infections
C2349858|ICD9CM|PT|059.8|Other poxvirus infections
C2349858|ICD9CM|AB|059.8|Poxvirus infections NEC
C2349859|ICD9CM|AB|V23.85|Pregnt-assist repro tech
C2349859|ICD9CM|PT|V23.85|Pregnancy resulting from assisted reproductive technology
C2349861|ICD9CM|PT|V23.86|Pregnancy with history of in utero procedure during previous pregnancy
C2349861|ICD9CM|AB|V23.86|Preg-hx in utro prev prg
C2349862|ICD9CM|PT|V28.3|Encounter for routine screening for malformation using ultrasonics
C2349862|ICD9CM|AB|V28.3|Scr fetl malfrm-ultrasnd
C2349864|ICD9CM|PT|V28.81|Encounter for fetal anatomic survey
C2349864|ICD9CM|AB|V28.81|Scrn fetal anatmc survey
C2349865|ICD9CM|PT|V28.82|Encounter for screening for risk of pre-term labor
C2349865|ICD9CM|AB|V28.82|Scrn risk preterm labor
C2349872|ICD9CM|AB|V45.12|Noncmplnt w renal dialys
C2349872|ICD9CM|PT|V45.12|Noncompliance with renal dialysis
C2349873|ICD9CM|AB|V45.71|Acq absnce breast/nipple
C2349873|ICD9CM|PT|V45.71|Acquired absence of breast and nipple
C2349874|ICD9CM|PT|V45.87|Transplanted organ removal status
C2349874|ICD9CM|AB|V45.87|Trnsplnt orgn rem status
C2349876|ICD9CM|PT|V45.88|Status post administration of tPA (rtPA) in a different facility within the last 24 hours prior to admission to current facility
C2349876|ICD9CM|AB|V45.88|TPA adm status 24 hr pta
C2349878|ICD9CM|HT|V46|Other dependence on machines and devices
C2349879|ICD9CM|PT|V51.0|Encounter for breast reconstruction following mastectomy
C2349879|ICD9CM|AB|V51.0|Brst reconst fol mastect
C2349880|ICD9CM|AB|V51.8|Aftercre plastc surg NEC
C2349880|ICD9CM|PT|V51.8|Other aftercare involving the use of plastic surgery
C2349886|ICD9CM|PT|V61.01|Family disruption due to family member on military deployment
C2349886|ICD9CM|AB|V61.01|Fmily dsrpt-fam military
C2349888|ICD9CM|PT|V61.02|Family disruption due to return of family member from military deployment
C2349888|ICD9CM|AB|V61.02|Fmily dsrpt-ret military
C2349890|ICD9CM|AB|V61.03|Fmily dsrpt- divorce/sep
C2349890|ICD9CM|PT|V61.03|Family disruption due to divorce or legal separation
C2349891|ICD9CM|PT|V61.04|Family disruption due to parent-child estrangement
C2349891|ICD9CM|AB|V61.04|Family dsrpt-estrangmemt
C2349892|ICD9CM|AB|V61.05|Famly dsrpt-chld custody
C2349892|ICD9CM|PT|V61.05|Family disruption due to child in welfare custody
C2349893|ICD9CM|AB|V61.06|Family dsrpt-foster care
C2349893|ICD9CM|PT|V61.06|Family disruption due to child in foster care or in care of non-parental family member
C2349894|ICD9CM|AB|V61.09|Family disruption NEC
C2349894|ICD9CM|PT|V61.09|Other family disruption
C2349895|ICD9CM|PT|V62.21|Personal current military deployment status
C2349895|ICD9CM|AB|V62.21|Hx military deployment
C2349897|ICD9CM|PT|V62.22|Personal history of return from military deployment
C2349897|ICD9CM|AB|V62.22|Hx retrn military deploy
C2349899|ICD9CM|AB|V87.01|Contact/exposure arsenic
C2349899|ICD9CM|PT|V87.01|Contact with and (suspected) exposure to arsenic
C2349900|ICD9CM|PT|V87.09|Contact with and (suspected) exposure to other hazardous metals
C2349900|ICD9CM|AB|V87.09|Cntct/exp hazrd metl NEC
C2349903|ICD9CM|HT|V87.0|Contact with and (suspected) exposure to hazardous metals
C2349904|ICD9CM|AB|V87.11|Cntct/exp aromatc amines
C2349904|ICD9CM|PT|V87.11|Contact with and (suspected) exposure to aromatic amines
C2349905|ICD9CM|AB|V87.12|Contact/exposure benzene
C2349905|ICD9CM|PT|V87.12|Contact with and (suspected) exposure to benzene
C2349906|ICD9CM|AB|V87.19|Cont/exp haz aromat NEC
C2349906|ICD9CM|PT|V87.19|Contact with and (suspected) exposure to other hazardous aromatic compounds
C2349909|ICD9CM|HT|V87.1|Contact with and (suspected) exposure to hazardous aromatic compounds
C2349910|ICD9CM|AB|V87.2|Cont/exp hazard chem NEC
C2349910|ICD9CM|PT|V87.2|Contact with and (suspected) exposure to other potentially hazardous chemicals
C2349912|ICD9CM|PT|V87.39|Contact with and (suspected) exposure to other potentially hazardous substances
C2349912|ICD9CM|HT|V87.3|Contact with and (suspected ) exposure to other potentially hazardous substances
C2349912|ICD9CM|AB|V87.39|Cont/exp hazard sub NEC
C2349913|ICD9CM|PT|V87.41|Personal history of antineoplastic chemotherapy
C2349913|ICD9CM|AB|V87.41|Hx antineoplastic chemo
C2349914|ICD9CM|PT|V87.42|Personal history of monoclonal drug therapy
C2349914|ICD9CM|AB|V87.42|Hx monoclonal drug thrpy
C2349915|ICD9CM|PT|V87.49|Personal history of other drug therapy
C2349915|ICD9CM|AB|V87.49|Hx drug therapy NEC
C2349916|ICD9CM|HT|V87.4|Personal history of drug therapy
C2349917|ICD9CM|HT|V87-V87.99|OTHER SPECIFIED PERSONAL EXPOSURES AND HISTORY PRESENTING HAZARDS TO HEALTH
C2349917|ICD9CM|HT|V87|Other specified personal exposures and history presenting hazards to health
C2349918|ICD9CM|HT|V88|Acquired absence of other organs and tissue
C2349918|ICD9CM|HT|V88-V88.99|ACQUIRED ABSENCE OF OTHER ORGANS AND TISSUE
C2349919|ICD9CM|AB|V88.01|Acq absnce cervix/uterus
C2349919|ICD9CM|PT|V88.01|Acquired absence of both cervix and uterus
C2349922|ICD9CM|PT|V88.02|Acquired absence of uterus with remaining cervical stump
C2349922|ICD9CM|AB|V88.02|Acq ab ut remn cerv stmp
C2349924|ICD9CM|AB|V88.03|Acq absnc cerv/remain ut
C2349924|ICD9CM|PT|V88.03|Acquired absence of cervix with remaining uterus
C2349925|ICD9CM|HT|V88.0|Acquired absence of cervix and uterus
C2349926|ICD9CM|PT|V89.01|Suspected problem with amniotic cavity and membrane not found
C2349926|ICD9CM|AB|V89.01|Sus amntc cav/mem nt fnd
C2349929|ICD9CM|PT|V89.02|Suspected placental problem not found
C2349929|ICD9CM|AB|V89.02|Sus placentl prob nt fnd
C2349930|ICD9CM|PT|V89.03|Suspected fetal anomaly not found
C2349930|ICD9CM|AB|V89.03|Sus fetal anomaly nt fnd
C2349931|ICD9CM|AB|V89.04|Sus fetal growth not fnd
C2349931|ICD9CM|PT|V89.04|Suspected problem with fetal growth not found
C2349932|ICD9CM|AB|V89.05|Sus cervcl shortn nt fnd
C2349932|ICD9CM|PT|V89.05|Suspected cervical shortening not found
C2349933|ICD9CM|PT|V89.09|Other suspected maternal and fetal condition not found
C2349933|ICD9CM|AB|V89.09|Oth sus mat/ftl nt fnd
C2349934|ICD9CM|HT|V89.0|Suspected maternal and fetal conditions not found
C2349935|ICD9CM|HT|V89-V89.99|OTHER SUSPECTED CONDITIONS NOT FOUND
C2349935|ICD9CM|HT|V89|Other suspected conditions not found
C2349953|ICD9CM|PT|750.13|Fissure of tongue
C2349953|ICD9CM|AB|750.13|Cong fissure of tongue
C2350012|ICD9CM|AB|V02.54|Meth resis Staph carrier
C2350012|ICD9CM|AB|V12.04|Hx Methicln resist Staph
C2350012|ICD9CM|PT|V12.04|Personal history of Methicillin resistant Staphylococcus aureus
C2350012|ICD9CM|PT|V02.54|Carrier or suspected carrier of Methicillin resistant Staphylococcus aureus
C2350019|ICD9CM|PT|793.11|Solitary pulmonary nodule
C2350019|ICD9CM|AB|793.11|Solitary pulmonry nodule
C2350236|ICD9CM|HT|516.3|Idiopathic interstitial pneumonia
C2350476|ICD9CM|AB|376.12|Orbital myositis
C2350476|ICD9CM|PT|376.12|Orbital myositis
C2350621|ICD9CM|AB|117.4|Mycotic mycetomas
C2350621|ICD9CM|PT|117.4|Mycotic mycetomas
C2355591|ICD9CM|PT|V02.53|Carrier or suspected carrier of Methicillin susceptible Staphylococcus aureus
C2355591|ICD9CM|AB|V02.53|Meth susc Staph carrier
C2355609|ICD9CM|AB|039.4|Madura foot
C2355609|ICD9CM|PT|039.4|Madura foot
C2355645|ICD9CM|AB|723.2|Cervicocranial syndrome
C2355645|ICD9CM|PT|723.2|Cervicocranial syndrome
C2362603|ICD9CM|PT|V87.31|Contact with and (suspected) exposure to mold
C2362603|ICD9CM|AB|V87.31|Contact/exposure mold
C2362836|ICD9CM|PT|346.80|Other forms of migraine, without mention of intractable migraine without mention of status migrainosus
C2362836|ICD9CM|AB|346.80|Othr migrne wo ntrc mgrn
C2363246|ICD9CM|HT|757.3|Other specified congenital anomalies of skin
C2363246|ICD9CM|PT|757.39|Other specified anomalies of skin
C2363246|ICD9CM|AB|757.39|Skin anomaly NEC
C2363280|ICD9CM|AB|744.43|Cervical auricle
C2363280|ICD9CM|PT|744.43|Cervical auricle
C2363337|ICD9CM|PT|V46.2|Other dependence on machines, supplemental oxygen
C2363337|ICD9CM|AB|V46.2|Depend-supplement oxygen
C2368006|ICD9CM|PT|059.10|Parapoxvirus infection, unspecified
C2368006|ICD9CM|AB|059.10|Parapoxvirus infectn NOS
C2454646|ICD9CM|PT|88.93|Magnetic resonance imaging of spinal canal
C2454646|ICD9CM|AB|88.93|Mri spinal canal
C2585165|ICD9CM|PT|789.42|Abdominal rigidity, left upper quadrant
C2585165|ICD9CM|AB|789.42|Abdmnal rgdt lft up quad
C2585306|ICD9CM|PT|789.64|Abdominal tenderness, left lower quadrant
C2585306|ICD9CM|AB|789.64|Abdmnal tndr lt lwr quad
C2585545|ICD9CM|PT|789.43|Abdominal rigidity, right lower quadrant
C2585545|ICD9CM|AB|789.43|Abdmnal rgdt rt lwr quad
C2585546|ICD9CM|PT|789.44|Abdominal rigidity, left lower quadrant
C2585546|ICD9CM|AB|789.44|Abdmnal rgdt lt lwr quad
C2586326|MTH|PN|NOCODE|Encounter due to family history of other lymphatic and hematopoietic neoplasms NEC in ICD9CM
C2586326|ICD9CM|PT|V16.7|Family history of other lymphatic and hematopoietic neoplasms
C2586326|ICD9CM|AB|V16.7|Fam hx-lymph neoplas NEC
C2586327|MTH|PN|NOCODE|Encounter due to screening for other hemoglobinopathies NEC in ICD9CM
C2586327|ICD9CM|PT|V78.3|Screening for other hemoglobinopathies
C2586327|ICD9CM|AB|V78.3|Scrn-hemoglobinopath NEC
C2586328|MTH|PN|NOCODE|Encounter due to other problems of limbs NEC in ICD9CM
C2586328|ICD9CM|PT|V49.5|Other problems of limbs
C2586328|ICD9CM|AB|V49.5|Limb problems NEC
C2607914|ICD9CM|HT|477|Allergic rhinitis
C2607914|ICD9CM|AB|477.9|Allergic rhinitis NOS
C2607914|ICD9CM|PT|477.9|Allergic rhinitis, cause unspecified
C2607928|ICD9CM|AB|366.00|Nonsenile cataract NOS
C2607928|ICD9CM|PT|366.00|Nonsenile cataract, unspecified
C2607948|ICD9CM|HT|013.3|Tuberculous abscess of brain
C2607950|ICD9CM|PT|163.1|Malignant neoplasm of visceral pleura
C2607950|ICD9CM|AB|163.1|Mal neo visceral pleura
C2609444|MTH|PN|NOCODE|Other orbital disorders NEC in ICD9CM
C2609444|ICD9CM|AB|376.89|Orbital disorders NEC
C2609444|ICD9CM|PT|376.89|Other orbital disorders
C2699510|ICD9CM|AB|755.58|Congenital cleft hand
C2699510|ICD9CM|PT|755.58|Cleft hand, congenital
C2711042|ICD9CM|PT|200.76|Large cell lymphoma, intrapelvic lymph nodes
C2711042|ICD9CM|AB|200.76|Large cell lymph pelvic
C2711059|ICD9CM|PT|327.11|Idiopathic hypersomnia with long sleep time
C2711059|ICD9CM|AB|327.11|Idio hypersom-long sleep
C2711060|ICD9CM|PT|V83.81|Cystic fibrosis gene carrier
C2711060|ICD9CM|AB|V83.81|Cystic fibrosis gene car
C2711232|ICD9CM|PT|327.24|Idiopathic sleep related non-obstructive alveolar hypoventilation
C2711232|ICD9CM|AB|327.24|Idiopath sleep hypovent
C2711480|ICD9CM|PT|428.32|Chronic diastolic heart failure
C2711480|ICD9CM|AB|428.32|Chr diastolic hrt fail
C2711630|ICD9CM|PT|279.2|Combined immunity deficiency
C2711630|ICD9CM|AB|279.2|Combined immunity defic
C2711750|ICD9CM|AB|618.02|Cystocele, lateral
C2711750|ICD9CM|PT|618.02|Cystocele, lateral
C2711774|ICD9CM|PT|525.71|Osseointegration failure of dental implant
C2711774|ICD9CM|AB|525.71|Osseo fail dental implnt
C2711829|ICD9CM|PT|415.11|Iatrogenic pulmonary embolism and infarction
C2711829|ICD9CM|AB|415.11|Iatrogen pulm emb/infarc
C2711887|ICD9CM|PT|996.46|Articular bearing surface wear of prosthetic joint
C2711887|ICD9CM|AB|996.46|Articular wear prosth jt
C2711989|MTH|PN|NOCODE|Abnormal function study of cardiovascular system NEC in ICD9CM
C2711989|ICD9CM|PT|794.39|Other nonspecific abnormal results of function study of cardiovascular system
C2711989|ICD9CM|AB|794.39|Abn cardiovasc study NEC
C2712343|MTH|PN|NOCODE|ALLERGIC RHINITIS NEC in ICD9CM
C2712343|ICD9CM|PT|477.8|Allergic rhinitis due to other allergen
C2712343|ICD9CM|AB|477.8|Allergic rhinitis NEC
C2712345|ICD9CM|PT|670.10|Puerperal endometritis, unspecified as to episode of care or not applicable
C2712345|ICD9CM|AB|670.10|Puerp endometritis-unsp
C2712346|ICD9CM|PT|670.12|Puerperal endometritis, delivered, with mention of postpartum complication
C2712346|ICD9CM|AB|670.12|Puerp endomet del w p/p
C2712347|ICD9CM|PT|670.14|Puerperal endometritis, postpartum condition or complication
C2712347|ICD9CM|AB|670.14|Puerp endomet-postpart
C2712348|ICD9CM|PT|670.20|Puerperal sepsis, unspecified as to episode of care or not applicable
C2712348|ICD9CM|AB|670.20|Puerperal sepsis-unsp
C2712349|ICD9CM|PT|670.22|Puerperal sepsis, delivered, with mention of postpartum complication
C2712349|ICD9CM|AB|670.22|Puerprl sepsis-del w p/p
C2712350|ICD9CM|PT|670.24|Puerperal sepsis, postpartum condition or complication
C2712350|ICD9CM|AB|670.24|Puerperl sepsis-postpart
C2712351|ICD9CM|PT|670.30|Puerperal septic thrombophlebitis, unspecified as to episode of care or not applicable
C2712351|ICD9CM|AB|670.30|Puerp septc thromb-unsp
C2712352|ICD9CM|PT|670.32|Puerperal septic thrombophlebitis, delivered, with mention of postpartum complication
C2712352|ICD9CM|AB|670.32|Prp sptc thrmb-del w p/p
C2712353|ICD9CM|PT|670.34|Puerperal septic thrombophlebitis, postpartum condition or complication
C2712353|ICD9CM|AB|670.34|Prp septc thrmb-postpart
C2712354|ICD9CM|PT|670.80|Other major puerperal infection, unspecified as to episode of care or not applicable
C2712354|ICD9CM|AB|670.80|Maj prp infec NEC-unspec
C2712355|ICD9CM|PT|670.82|Other major puerperal infection, delivered, with mention of postpartum complication
C2712355|ICD9CM|AB|670.82|Maj prp inf NEC-dl w p/p
C2712356|ICD9CM|PT|670.84|Other major puerperal infection, postpartum condition or complication
C2712356|ICD9CM|AB|670.84|Maj puerp infec NEC-p/p
C2712358|ICD9CM|PT|768.71|Mild hypoxic-ischemic encephalopathy
C2712358|ICD9CM|AB|768.71|Mild hypox-ischem enceph
C2712359|ICD9CM|PT|768.72|Moderate hypoxic-ischemic encephalopathy
C2712359|ICD9CM|AB|768.72|Mod hypox-ischem enceph
C2712360|ICD9CM|PT|768.73|Severe hypoxic-ischemic encephalopathy
C2712360|ICD9CM|AB|768.73|Sev hypox-ischem enceph
C2712362|ICD9CM|PT|779.32|Bilious vomiting in newborn
C2712362|ICD9CM|AB|779.32|NB bilious vomiting
C2712363|ICD9CM|PT|779.33|Other vomiting in newborn
C2712363|ICD9CM|AB|779.33|NB other vomiting
C2712364|ICD9CM|PT|779.34|Failure to thrive in newborn
C2712364|ICD9CM|AB|779.34|NB failure to thrive
C2712365|ICD9CM|PT|784.40|Voice and resonance disorder, unspecified
C2712365|ICD9CM|AB|784.40|Voice/resonance dis NOS
C2712366|ICD9CM|PT|784.49|Other voice and resonance disorders
C2712366|ICD9CM|AB|784.49|Voice/resonance dis NEC
C2712367|ICD9CM|PT|784.59|Other speech disturbance
C2712367|ICD9CM|AB|784.59|Speech disturbance NEC
C2712369|ICD9CM|PT|793.82|Inconclusive mammogram
C2712369|ICD9CM|AB|793.82|Inconclusive mammogram
C2712370|ICD9CM|PT|799.82|Apparent life threatening event in infant
C2712370|ICD9CM|AB|799.82|Appar life threat-infant
C2712371|ICD9CM|PT|813.45|Torus fracture of radius (alone)
C2712371|ICD9CM|AB|813.45|Torus fx radius-cl/alone
C2712372|ICD9CM|PT|813.46|Torus fracture of ulna (alone)
C2712372|ICD9CM|AB|813.46|Torus fx ulna-closed
C2712373|ICD9CM|PT|813.47|Torus fracture of radius and ulna
C2712373|ICD9CM|AB|813.47|Torus fx radius/ulna-clo
C2712374|ICD9CM|PT|969.00|Poisoning by antidepressant, unspecified
C2712374|ICD9CM|AB|969.00|Poison-antidepresnt NOS
C2712375|ICD9CM|PT|969.02|Poisoning by selective serotonin and norepinephrine reuptake inhibitors
C2712375|ICD9CM|AB|969.02|Pois serotn/norepinephrn
C2712376|ICD9CM|PT|969.03|Poisoning by selective serotonin reuptake inhibitors
C2712376|ICD9CM|AB|969.03|Pois serotinin reuptake
C2712377|ICD9CM|PT|969.04|Poisoning by tetracyclic antidepressants
C2712377|ICD9CM|AB|969.04|Pois tetracyclc andepres
C2712378|ICD9CM|PT|969.09|Poisoning by other antidepressants
C2712378|ICD9CM|AB|969.09|Pois antidepressants NEC
C2712379|ICD9CM|PT|969.70|Poisoning by psychostimulant, unspecified
C2712379|ICD9CM|AB|969.70|Pois psychostimulant NOS
C2712380|ICD9CM|PT|969.73|Poisoning by methylphenidate
C2712380|ICD9CM|AB|969.73|Poison by methylphendate
C2712381|ICD9CM|PT|969.79|Poisoning by other psychostimulants
C2712381|ICD9CM|AB|969.79|Poison by psychostim NEC
C2712382|ICD9CM|PT|995.24|Failed moderate sedation during procedure
C2712382|ICD9CM|AB|995.24|Fail mod sedate dur proc
C2712383|ICD9CM|PT|996.43|Broken prosthetic joint implant
C2712383|ICD9CM|AB|996.43|Broke prosthtc jt implnt
C2712384|ICD9CM|PT|E000.0|Civilian activity done for income or pay
C2712384|ICD9CM|AB|E000.0|Civilian activity-income
C2712385|ICD9CM|PT|E000.1|Military activity
C2712385|ICD9CM|AB|E000.1|Military activity
C2712386|ICD9CM|PT|E000.8|Other external cause status
C2712386|ICD9CM|AB|E000.8|Externl cause status NEC
C2712387|ICD9CM|PT|E000.9|Unspecified external cause status
C2712387|ICD9CM|AB|E000.9|Externl cause status NOS
C2712388|ICD9CM|PT|E001.0|Activities involving walking, marching and hiking
C2712388|ICD9CM|AB|E001.0|Walking,marching,hiking
C2712389|ICD9CM|PT|E002.1|Activities involving springboard and platform diving
C2712389|ICD9CM|AB|E002.1|Springboard/platfrm dive
C2712390|ICD9CM|AB|E002.2|Water polo
C2712390|ICD9CM|PT|E002.2|Activities involving water polo
C2712391|ICD9CM|PT|E002.3|Activities involving water aerobics and water exercise
C2712391|ICD9CM|AB|E002.3|Water aerobics/exercise
C2712392|ICD9CM|PT|E002.4|Activities involving underwater diving and snorkeling
C2712392|ICD9CM|AB|E002.4|Underwater dive/snorkel
C2712393|ICD9CM|PT|E002.5|Activities involving rowing, canoeing, kayaking, rafting and tubing
C2712393|ICD9CM|AB|E002.5|Row,canoe,kayk,raft,tube
C2712394|ICD9CM|PT|E002.6|Activities involving water skiing and wake boarding
C2712394|ICD9CM|AB|E002.6|Water ski/wake boarding
C2712395|ICD9CM|PT|E002.7|Activities involving surfing, windsurfing and boogie boarding
C2712395|ICD9CM|AB|E002.7|Surf,windsrf,boogie brd
C2712396|ICD9CM|PT|E002.8|Activities involving water sliding
C2712396|ICD9CM|AB|E002.8|Water sliding
C2712397|ICD9CM|PT|E002.9|Other activity involving water and watercraft
C2712397|ICD9CM|AB|E002.9|Water/watercraft
C2712398|ICD9CM|PT|E003.2|Activities involving snow (alpine) (downhill) skiing, snow boarding, sledding, tobogganing and snow tubing
C2712398|ICD9CM|AB|E003.2|Ski,snow brd,sled,tobagn
C2712399|ICD9CM|PT|E003.3|Activities involving cross country skiing
C2712399|ICD9CM|AB|E003.3|Cross country skiing
C2712400|ICD9CM|PT|E003.9|Other activity involving ice and snow
C2712400|ICD9CM|AB|E003.9|Ice and snow
C2712401|ICD9CM|PT|E004.0|Activities involving mountain climbing, rock climbing and wall climbing
C2712401|ICD9CM|AB|E004.0|Mountain,rock/wall climb
C2712402|ICD9CM|PT|E004.1|Activities involving rappelling
C2712402|ICD9CM|AB|E004.1|Rappelling
C2712403|ICD9CM|PT|E004.2|Activities involving BASE jumping
C2712403|ICD9CM|AB|E004.2|BASE jumping
C2712404|ICD9CM|PT|E004.9|Other activity involving climbing, rappelling and jumping off
C2712404|ICD9CM|AB|E004.9|Climb,rappell,jump off
C2712405|ICD9CM|PT|E005.3|Activities involving trampoline
C2712405|ICD9CM|AB|E005.3|Trampoline
C2712406|ICD9CM|PT|E005.9|Other activity involving dancing and other rhythmic movements
C2712406|ICD9CM|AB|E005.9|Dancing,rhythm movements
C2712407|ICD9CM|PT|E006.0|Activities involving roller skating (inline) and skateboarding
C2712407|ICD9CM|AB|E006.0|Roller skate,skateboard
C2712408|ICD9CM|AB|E006.4|Bike riding
C2712408|ICD9CM|PT|E006.4|Activities involving bike riding
C2712409|ICD9CM|PT|E006.5|Activities involving jumping rope
C2712409|ICD9CM|AB|E006.5|Jumping rope
C2712410|ICD9CM|PT|E006.6|Activities involving non-running track and field events
C2712410|ICD9CM|AB|E006.6|Non-running track/field
C2712411|ICD9CM|PT|E006.9|Other activity involving other sports and athletics played individually
C2712411|ICD9CM|AB|E006.9|Individ sports,athletics
C2712412|ICD9CM|PT|E007.0|Activities involving american tackle football
C2712412|ICD9CM|AB|E007.0|Tackle football
C2712413|ICD9CM|PT|E007.1|Activities involving american flag or touch football
C2712413|ICD9CM|AB|E007.1|Amer flag/touch football
C2712414|ICD9CM|PT|E007.4|Activities involving lacrosse and field hockey
C2712414|ICD9CM|AB|E007.4|Lacrosse,field hockey
C2712415|ICD9CM|PT|E007.7|Activities involving volleyball (beach) (court)
C2712415|ICD9CM|AB|E007.7|Volleyball (beach,court)
C2712416|ICD9CM|PT|E007.8|Activities involving physical games generally associated with school recess, summer camp and children
C2712416|ICD9CM|AB|E007.8|School recess,camp
C2712417|ICD9CM|PT|E007.9|Other activity involving other sports and athletes played as a team or group
C2712417|ICD9CM|AB|E007.9|Team sports,athletes
C2712418|ICD9CM|PT|E008.2|Activities involving racquet and hand sports
C2712418|ICD9CM|AB|E008.2|Racquet/hand sports
C2712419|ICD9CM|AB|E008.3|Frisbee
C2712419|ICD9CM|PT|E008.3|Activities involving frisbee
C2712420|ICD9CM|PT|E008.9|Other specified sports and athletics activity
C2712420|ICD9CM|AB|E008.9|Sports,athletics NEC
C2712421|ICD9CM|PT|E009.0|Activity involving exercise machines primarily for cardiorespiratory conditioning
C2712421|ICD9CM|AB|E009.0|Exercise mach(cardiorsp)
C2712422|ICD9CM|PT|E009.2|Activity involving aerobic and step exercise
C2712422|ICD9CM|AB|E009.2|Aerobic,step exercise
C2712423|ICD9CM|AB|E009.3|Circuit training
C2712423|ICD9CM|PT|E009.3|Activity involving circuit training
C2712424|ICD9CM|PT|E009.4|Activity involving obstacle course
C2712424|ICD9CM|AB|E009.4|Obstacle course
C2712425|ICD9CM|PT|E009.5|Activity involving grass drills
C2712425|ICD9CM|AB|E009.5|Grass drills
C2712426|ICD9CM|PT|E009.9|Other activity involving cardiorespiratory exercise
C2712426|ICD9CM|AB|E009.9|Cardioresp exercise NEC
C2712427|ICD9CM|PT|E010.0|Activity involving exercise machines primarily for muscle strengthening
C2712427|ICD9CM|AB|E010.0|Muscle strength mach
C2712428|ICD9CM|PT|E010.1|Activity involving push-ups, pull-ups, sit-ups
C2712428|ICD9CM|AB|E010.1|Push-ups,pull-ups,sit-up
C2712429|ICD9CM|PT|E010.2|Activity involving free weights
C2712429|ICD9CM|AB|E010.2|Free weights
C2712430|ICD9CM|PT|E010.3|Activity involving pilates
C2712430|ICD9CM|AB|E010.3|Pilates
C2712431|ICD9CM|PT|E010.9|Other activity involving other muscle strengthening exercises
C2712431|ICD9CM|AB|E010.9|Muscle strength exer NEC
C2712432|ICD9CM|PT|E011.0|Activities involving computer keyboarding
C2712432|ICD9CM|AB|E011.0|Computer keyboarding
C2712433|ICD9CM|PT|E011.1|Activities involving hand held interactive electronic device
C2712433|ICD9CM|AB|E011.1|Handheld interac elec dv
C2712434|ICD9CM|PT|E011.9|Other activity involving computer technology and electronic devices
C2712434|ICD9CM|AB|E011.9|Computer tech NEC
C2712435|ICD9CM|PT|E012.0|Activities involving knitting and crocheting
C2712435|ICD9CM|AB|E012.0|Knitting & crocheting
C2712436|ICD9CM|PT|E012.1|Activities involving sewing
C2712436|ICD9CM|AB|E012.1|Sewing
C2712437|ICD9CM|PT|E012.2|Activities involving furniture building and finishing
C2712437|ICD9CM|AB|E012.2|Furniture build/finish
C2712438|ICD9CM|PT|E012.9|Activity involving other arts and handcrafts
C2712438|ICD9CM|AB|E012.9|Arts & handcrafts NEC
C2712439|ICD9CM|PT|E013.0|Activities involving personal bathing and showering
C2712439|ICD9CM|AB|E013.0|Personal bathing/shower
C2712440|ICD9CM|PT|E013.4|Activities involving floor mopping and cleaning
C2712440|ICD9CM|AB|E013.4|Floor mopping/cleaning
C2712441|ICD9CM|PT|E013.5|Activities involving residential relocation
C2712441|ICD9CM|AB|E013.5|Residential relocation
C2712442|ICD9CM|PT|E013.8|Other personal hygiene activity
C2712442|ICD9CM|AB|E013.8|Personal hygiene NEC
C2712443|ICD9CM|PT|E013.9|Other household maintenance
C2712443|ICD9CM|AB|E013.9|Househld maintenance NEC
C2712444|ICD9CM|PT|E014.0|Caregiving involving bathing
C2712444|ICD9CM|AB|E014.0|Caregiving-bathing
C2712445|ICD9CM|PT|E014.1|Caregiving involving lifting
C2712445|ICD9CM|AB|E014.1|Caregiving-lifting
C2712446|ICD9CM|PT|E014.9|Other activity involving person providing caregiving
C2712446|ICD9CM|AB|E014.9|Caregiving NEC
C2712447|ICD9CM|PT|E015.0|Activities involving food preparation and clean up
C2712447|ICD9CM|AB|E015.0|Food prep & cleanup
C2712448|ICD9CM|PT|E015.1|Activities involving grilling and smoking food
C2712448|ICD9CM|AB|E015.1|Grilling & smoking food
C2712449|ICD9CM|PT|E015.2|Activities involving cooking and baking
C2712449|ICD9CM|AB|E015.2|Cooking & baking
C2712450|ICD9CM|PT|E015.9|Other activity involving cooking and grilling
C2712450|ICD9CM|AB|E015.9|Cooking & grilling NEC
C2712451|ICD9CM|PT|E016.0|Activities involving digging, shoveling and raking
C2712451|ICD9CM|AB|E016.0|Digging,shovel,rake
C2712452|ICD9CM|PT|E016.1|Activities involving gardening and landscaping
C2712452|ICD9CM|AB|E016.1|Gardening/landscaping
C2712453|ICD9CM|PT|E016.2|Activities involving building and construction
C2712453|ICD9CM|AB|E016.2|Building & construction
C2712454|ICD9CM|PT|E016.9|Other activity involving property and land maintenance, building and construction
C2712454|ICD9CM|AB|E016.9|Land maintain/cnstrt NEC
C2712456|ICD9CM|PT|E017.9|Other activity involving external motion
C2712456|ICD9CM|AB|E017.9|External motion NEC
C2712457|ICD9CM|PT|E018.0|Activities involving piano playing
C2712457|ICD9CM|AB|E018.0|Piano playing
C2712458|ICD9CM|PT|E018.1|Activities involving drum and other percussion instrument playing
C2712458|ICD9CM|AB|E018.1|Drum/percussion playing
C2712459|ICD9CM|PT|E018.2|Activities involving string instrument playing
C2712459|ICD9CM|AB|E018.2|String instrument play
C2712460|ICD9CM|PT|E018.3|Activities involving winds and brass instrument playing
C2712460|ICD9CM|AB|E018.3|Winds/brass instru play
C2712461|ICD9CM|PT|E019.0|Activities involving walking an animal
C2712461|ICD9CM|AB|E019.0|Walking an animal
C2712462|ICD9CM|PT|E019.1|Activities involving milking an animal
C2712462|ICD9CM|AB|E019.1|Milking an animal
C2712463|ICD9CM|PT|E019.2|Activities involving grooming and shearing an animal
C2712463|ICD9CM|AB|E019.2|Groom/shearing animal
C2712464|ICD9CM|PT|E019.9|Other activity involving animal care
C2712464|ICD9CM|AB|E019.9|Animal care NEC
C2712465|ICD9CM|AB|E029.0|Refereeing sports
C2712465|ICD9CM|PT|E029.0|Refereeing a sports activity
C2712466|ICD9CM|AB|E029.1|Spectator at event
C2712466|ICD9CM|PT|E029.1|Spectator at an event
C2712467|ICD9CM|PT|E029.2|Rough housing and horseplay
C2712467|ICD9CM|AB|E029.2|Rough housing/horseplay
C2712469|ICD9CM|PT|E830.7|Accident to watercraft causing submersion, occupant of military watercraft, any type
C2712469|ICD9CM|AB|E830.7|Boat submers-military
C2712470|ICD9CM|PT|E831.7|Accident to watercraft causing other injury, occupant of military watercraft, any type
C2712470|ICD9CM|AB|E831.7|Boat acc inj NEC-militry
C2712471|ICD9CM|PT|E832.7|Other accidental submersion or drowning in water transport accident, occupant of military watercraft, any type
C2712471|ICD9CM|AB|E832.7|Submersion NEC-military
C2712472|ICD9CM|PT|E833.7|Fall on stairs or ladders in water transport, occupant of military watercraft, any type
C2712472|ICD9CM|AB|E833.7|W/crf stair fall-militry
C2712473|ICD9CM|PT|E834.7|Other fall from one level to another in water transport, occupant of military watercraft, any type
C2712473|ICD9CM|AB|E834.7|W/crft fall NEC-military
C2712474|ICD9CM|PT|E835.7|Other and unspecified fall in water transport, occupant of military watercraft, any type
C2712474|ICD9CM|AB|E835.7|W/crft fall NEC/NOS-mil
C2712475|ICD9CM|PT|E836.7|Machinery accident in water transport, occupant of military watercraft, any type
C2712475|ICD9CM|AB|E836.7|W/crft machine-military
C2712476|ICD9CM|PT|E837.7|Explosion, fire, or burning in watercraft, occupant of military watercraft, any type
C2712476|ICD9CM|AB|E837.7|W/crft explosn-military
C2712477|ICD9CM|PT|E838.7|Other and unspecified water transport accident, occupant of military watercraft, any type
C2712477|ICD9CM|AB|E838.7|W/crft-military NEC/NOS
C2712478|ICD9CM|PT|E876.5|Performance of wrong operation (procedure) on correct patient
C2712478|ICD9CM|AB|E876.5|Perfrm wrong op/right pt
C2712479|ICD9CM|PT|E876.6|Performance of operation (procedure) on patient not scheduled for surgery
C2712479|ICD9CM|AB|E876.6|Proc-pt not sched surg
C2712480|ICD9CM|PT|E876.7|Performance of correct operation (procedure) on wrong side/body part
C2712480|ICD9CM|AB|E876.7|Rt proc-wrong side/part
C2712481|ICD9CM|PT|E928.7|Environmental and accidental causes, mechanism or component of firearm and air gun
C2712481|ICD9CM|AB|E928.7|Accidnt-mech firearm/gun
C2712482|ICD9CM|PT|E990.1|Injury due to war operations from flamethrower
C2712482|ICD9CM|AB|E990.1|War inj:flamethrower
C2712483|ICD9CM|PT|E990.2|Injury due to war operations from incendiary bullet
C2712483|ICD9CM|AB|E990.2|War inj:incndiary bullet
C2712484|ICD9CM|PT|E990.3|Injury due to war operations from fire caused indirectly from conventional weapon
C2712484|ICD9CM|AB|E990.3|War inj:ind convn weapn
C2712485|ICD9CM|PT|E991.4|Injury due to war operations by fragments from munitions
C2712485|ICD9CM|AB|E991.4|War inj:munition fragmnt
C2712486|ICD9CM|PT|E991.5|Injury due to war operations by fragments from person-borne improvised explosive device [IED]
C2712486|ICD9CM|AB|E991.5|War inj:prsn-brn fragmnt
C2712487|ICD9CM|PT|E991.6|Injury due to war operations by fragments from vehicle-borne improvised explosive device [IED]
C2712487|ICD9CM|AB|E991.6|War inj:vehic-borne IED
C2712488|ICD9CM|PT|E991.7|Injury due to war operations by fragments from other improvised explosive device [IED]
C2712488|ICD9CM|AB|E991.7|War inj:fragment IED NEC
C2712489|ICD9CM|PT|E991.8|Injury due to war operations by fragments from weapons
C2712489|ICD9CM|AB|E991.8|War inj:weapon fragments
C2712490|ICD9CM|PT|E992.0|Injury due to torpedo
C2712490|ICD9CM|AB|E992.0|War inj:torpedo
C2712491|ICD9CM|PT|E992.1|Injury due to depth charge
C2712491|ICD9CM|AB|E992.1|War inj:depth charge
C2712492|ICD9CM|PT|E992.2|Injury due to marine mines
C2712492|ICD9CM|AB|E992.2|War inj:marine mines
C2712493|ICD9CM|PT|E992.3|Injury due to sea-based artillery shell
C2712493|ICD9CM|AB|E992.3|War inj:seabase art shel
C2712494|ICD9CM|PT|E992.8|Injury due to war operations by other marine weapons
C2712494|ICD9CM|AB|E992.8|War inj:marine weapn NEC
C2712495|ICD9CM|PT|E992.9|Injury due to war operations by unspecified marine weapon
C2712495|ICD9CM|AB|E992.9|War inj:marine weapn NOS
C2712496|ICD9CM|PT|E993.0|Injury due to war operations by aerial bomb
C2712496|ICD9CM|AB|E993.0|War inj:aerial bomb
C2712497|ICD9CM|PT|E993.1|Injury due to war operations by guided missile
C2712497|ICD9CM|AB|E993.1|War inj:guided missile
C2712498|ICD9CM|PT|E993.2|Injury due to war operations by mortar
C2712498|ICD9CM|AB|E993.2|War inj:mortar
C2712499|ICD9CM|PT|E993.3|Injury due to war operations by person-borne improvised explosive device [IED]
C2712499|ICD9CM|AB|E993.3|War inj:person IED
C2712500|ICD9CM|PT|E993.4|Injury due to war operations by vehicle-borne improvised explosive device [IED]
C2712500|ICD9CM|AB|E993.4|War inj:vehicle IED
C2712501|ICD9CM|PT|E993.5|Injury due to war operations by other improvised explosive device [IED]
C2712501|ICD9CM|AB|E993.5|War inj:IED NEC
C2712502|ICD9CM|PT|E993.6|Injury due to war operations by unintentional detonation of own munitions
C2712502|ICD9CM|AB|E993.6|War inj:acc own munition
C2712503|ICD9CM|PT|E993.7|Injury due to war operations by unintentional discharge of own munitions launch device
C2712503|ICD9CM|AB|E993.7|War inj:acc disch launch
C2712504|ICD9CM|PT|E993.8|Injury due to war operations by other specified explosion
C2712504|ICD9CM|AB|E993.8|War inj:explosion NEC
C2712505|ICD9CM|PT|E994.0|Injury due to war operations by destruction of aircraft due to enemy fire or explosives
C2712505|ICD9CM|AB|E994.0|War inj:aircrft des-enmy
C2712506|ICD9CM|PT|E994.1|Injury due to war operations by unintentional destruction of aircraft due to own onboard explosives
C2712506|ICD9CM|AB|E994.1|War inj:aircrft-own expl
C2712507|ICD9CM|PT|E994.2|Injury due to war operations by destruction of aircraft due to collision with other aircraft
C2712507|ICD9CM|AB|E994.2|War inj:aircrft collisn
C2712508|ICD9CM|PT|E994.3|Injury due to war operations by destruction of aircraft due to onboard fire
C2712508|ICD9CM|AB|E994.3|War inj:aircraft fire
C2712509|ICD9CM|PT|E994.8|Injury due to war operations by other destruction of aircraft
C2712509|ICD9CM|AB|E994.8|War inj:aircrft dest NEC
C2712510|ICD9CM|PT|E994.9|Injury due to war operations by unspecified destruction of aircraft
C2712510|ICD9CM|AB|E994.9|War inj:aircrft dest NOS
C2712511|ICD9CM|PT|E995.0|Injury due to war operations by unarmed hand-to-hand combat
C2712511|ICD9CM|AB|E995.0|War inj:hnd-hnd combat
C2712512|ICD9CM|PT|E995.1|Injury due to war operations, struck by blunt object
C2712512|ICD9CM|AB|E995.1|War inj:blunt object
C2712513|ICD9CM|PT|E995.2|Injury due to war operations by piercing object
C2712513|ICD9CM|AB|E995.2|War inj:piercing object
C2712514|ICD9CM|PT|E995.3|Injury due to war operations by intentional restriction of air and airway
C2712514|ICD9CM|AB|E995.3|War inj:intn restrct air
C2712515|ICD9CM|PT|E995.4|Injury due to war operations by unintentional drowning due to inability to surface or obtain air
C2712515|ICD9CM|AB|E995.4|War inj:unintentl drown
C2712516|ICD9CM|PT|E995.8|Injury due to war operations by other forms of conventional warfare
C2712516|ICD9CM|AB|E995.8|War inj:con warfare NEC
C2712517|ICD9CM|PT|E995.9|Injury due to war operations by unspecified form of conventional warfare
C2712517|ICD9CM|AB|E995.9|War inj:con warfare NOS
C2712518|ICD9CM|PT|E996.0|Injury due to war operations by direct blast effect of nuclear weapon
C2712518|ICD9CM|AB|E996.0|War inj:dir nucl weapon
C2712519|ICD9CM|PT|E996.1|Injury due to war operations by indirect blast effect of nuclear weapon
C2712519|ICD9CM|AB|E996.1|War inj:indir nucl weapn
C2712520|ICD9CM|PT|E996.2|Injury due to war operations by thermal radiation effect of nuclear weapon
C2712520|ICD9CM|AB|E996.2|War inj:therml radiation
C2712521|ICD9CM|PT|E996.3|Injury due to war operations by nuclear radiation effects
C2712521|ICD9CM|AB|E996.3|War inj:nuclear rad eff
C2712522|ICD9CM|PT|E996.8|Injury due to war operations by other effects of nuclear weapons
C2712522|ICD9CM|AB|E996.8|War inj:nucl weapon NEC
C2712523|ICD9CM|PT|E996.9|Injury due to war operations by unspecified effect of nuclear weapon
C2712523|ICD9CM|AB|E996.9|War inj:nucl weapon NOS
C2712524|ICD9CM|PT|E997.3|Injury due to war operations by weapon of mass destruction [WMD], unspecified
C2712524|ICD9CM|AB|E997.3|War inj:WMD NOS
C2712525|ICD9CM|PT|E998.0|Injury due to war operations but occurring after cessation of hostilities by explosion of mines
C2712525|ICD9CM|AB|E998.0|War inj:expl mine-cease
C2712526|ICD9CM|PT|E998.1|Injury due to war operations but occurring after cessation of hostilities by explosion of bombs
C2712526|ICD9CM|AB|E998.1|War inj:expl bomb-cease
C2712527|ICD9CM|PT|E998.8|Injury due to other war operations but occurring after cessation of hostilities
C2712527|ICD9CM|AB|E998.8|War inj:after cease NEC
C2712528|ICD9CM|PT|E998.9|Injury due to unspecified war operations but occurring after cessation of hostilities
C2712528|ICD9CM|AB|E998.9|War inj:after cease NOS
C2712534|ICD9CM|PT|39.75|Endovascular embolization or occlusion of vessel(s) of head or neck using bare coils
C2712534|ICD9CM|AB|39.75|Endo emb hd/nk,bare coil
C2712538|ICD9CM|PT|V15.06|Allergy to insects and arachnids
C2712538|ICD9CM|AB|V15.06|Hx-allergy insct/arachnd
C2712539|ICD9CM|AB|V15.52|Hx traumatc brain injury
C2712539|ICD9CM|PT|V15.52|Personal history of traumatic brain injury
C2712540|ICD9CM|AB|V15.80|Hx failed mod sedation
C2712540|ICD9CM|PT|V15.80|Personal history of failed moderate sedation
C2712541|ICD9CM|PT|V15.83|Personal history of underimmunization status
C2712541|ICD9CM|AB|V15.83|Hx underimmunizn status
C2712542|ICD9CM|PT|V15.84|Personal history of contact with and (suspected) exposure to asbestos
C2712542|ICD9CM|AB|V15.84|Hx-contct/expos asbestos
C2712543|ICD9CM|PT|V15.85|Personal history of contact with and (suspected) exposure to potentially hazardous body fluids
C2712543|ICD9CM|AB|V15.85|Hx-cont/exps haz bdy fld
C2712545|ICD9CM|PT|V20.31|Health supervision for newborn under 8 days old
C2712545|ICD9CM|AB|V20.31|Health supvsn nb <8 days
C2712546|ICD9CM|PT|V20.32|Health supervision for newborn 8 to 28 days old
C2712546|ICD9CM|AB|V20.32|Health supv nb 8-28 days
C2712547|ICD9CM|PT|V26.42|Encounter for fertility preservation counseling
C2712547|ICD9CM|AB|V26.42|Fertlity preserv counsel
C2712548|ICD9CM|PT|V26.82|Encounter for fertility preservation procedure
C2712548|ICD9CM|AB|V26.82|Fertility preserv proc
C2712549|ICD9CM|PT|V53.50|Fitting and adjustment of intestinal appliance and device
C2712549|ICD9CM|AB|V53.50|Fit/adjust intestinl dev
C2712551|ICD9CM|AB|V60.81|Foster care (status)
C2712551|ICD9CM|PT|V60.81|Foster care (status)
C2712552|ICD9CM|PT|V61.07|Family disruption due to death of family member
C2712552|ICD9CM|AB|V61.07|Family dsrpt-death membr
C2712553|ICD9CM|PT|V61.08|Family disruption due to other extended absence of family member
C2712553|ICD9CM|AB|V61.08|Fmly dsrp-fam absnce NEC
C2712554|ICD9CM|AB|V61.23|Cnsl prnt-biol chld prob
C2712554|ICD9CM|PT|V61.23|Counseling for parent-biological child problem
C2712555|ICD9CM|AB|V61.24|Cnsl prnt-adpt chld prob
C2712555|ICD9CM|PT|V61.24|Counseling for parent-adopted child problem
C2712556|ICD9CM|PT|V61.25|Counseling for parent (guardian)-foster child problem
C2712556|ICD9CM|AB|V61.25|Cnsl prnt-fstr chld prob
C2712557|ICD9CM|PT|V61.42|Substance abuse in family
C2712557|ICD9CM|AB|V61.42|Substance abuse-family
C2712559|ICD9CM|PT|V72.60|Laboratory examination, unspecified
C2712559|ICD9CM|AB|V72.60|Laboratory exam NOS
C2712560|ICD9CM|PT|V72.61|Antibody response examination
C2712560|ICD9CM|AB|V72.61|Antibody response exam
C2712561|ICD9CM|PT|V72.62|Laboratory examination ordered as part of a routine general medical examination
C2712561|ICD9CM|AB|V72.62|Routine physicl lab exam
C2712562|ICD9CM|PT|V72.63|Pre-procedural laboratory examination
C2712562|ICD9CM|AB|V72.63|Pre-procedure lab exam
C2712563|ICD9CM|PT|V72.69|Other laboratory examination
C2712563|ICD9CM|AB|V72.69|Laboratory exam NEC
C2712564|ICD9CM|PT|V80.09|Special screening for other neurological conditions
C2712564|ICD9CM|AB|V80.09|Screen-neuro condition
C2712565|ICD9CM|PT|V87.32|Contact with and (suspected) exposure to algae bloom
C2712565|ICD9CM|AB|V87.32|Contact/exp algae bloom
C2712566|ICD9CM|PT|V87.43|Personal history of estrogen therapy
C2712566|ICD9CM|AB|V87.43|Hx estrogen therapy
C2712567|ICD9CM|PT|V87.44|Personal history of inhaled steroid therapy
C2712567|ICD9CM|AB|V87.44|Hx inhaled steroid thrpy
C2712569|ICD9CM|PT|17.51|Implantation of rechargeable cardiac contractility modulation [CCM], total system
C2712569|ICD9CM|AB|17.51|Implant CCM,total system
C2712570|ICD9CM|PT|17.52|Implantation or replacement of cardiac contractility modulation [CCM] rechargeable pulse generator only
C2712570|ICD9CM|AB|17.52|Implant CCM pulse genrtr
C2712571|ICD9CM|PT|17.61|Laser interstitial thermal therapy [LITT] of lesion or tissue of brain under guidance
C2712571|ICD9CM|AB|17.61|LITT lesn brain,guidance
C2712572|ICD9CM|PT|17.62|Laser interstitial thermal therapy [LITT] of lesion or tissue of head and neck under guidance
C2712572|ICD9CM|AB|17.62|LITT les hd/nck,guidance
C2712573|ICD9CM|PT|17.63|Laser interstitial thermal therapy [LITT] of lesion or tissue of liver under guidance
C2712573|ICD9CM|AB|17.63|LITT lesn liver,guidance
C2712574|ICD9CM|PT|17.69|Laser interstitial thermal therapy [LITT] of lesion or tissue of other and unspecified site under guidance
C2712574|ICD9CM|AB|17.69|LITT lesn, guide oth/NOS
C2712575|ICD9CM|PT|17.70|Intravenous infusion of clofarabine
C2712575|ICD9CM|AB|17.70|IV infusion clofarabine
C2712576|ICD9CM|PT|33.73|Endoscopic insertion or replacement of bronchial valve(s), multiple lobes
C2712576|ICD9CM|AB|33.73|Endo ins/re brnc val,mul
C2712577|ICD9CM|PT|38.24|Intravascular imaging of coronary vessel(s) by optical coherence tomography [OCT]
C2712577|ICD9CM|AB|38.24|Intravas img cor ves OCT
C2712578|ICD9CM|PT|38.25|Intravascular imaging of non-coronary vessel(s) by optical coherence tomography [OCT]
C2712578|ICD9CM|AB|38.25|Intravas img non-cor OCT
C2712579|ICD9CM|PT|39.72|Endovascular (total) embolization or occlusion of head and neck vessels
C2712579|ICD9CM|AB|39.72|Endovasc embol hd/nk ves
C2712580|ICD9CM|PT|39.76|Endovascular embolization or occlusion of vessel(s) of head or neck using bioactive coils
C2712580|ICD9CM|AB|39.76|Endo em hd/nk,bioac coil
C2712581|ICD9CM|PT|39.79|Other endovascular procedures on other vessels
C2712581|ICD9CM|AB|39.79|Oth endo proc oth vessel
C2712582|ICD9CM|PT|39.90|Insertion of non-drug-eluting peripheral (non-coronary) vessel stent(s)
C2712582|ICD9CM|AB|39.90|Ins non-d-e non-cor stnt
C2712583|ICD9CM|PT|46.86|Endoscopic insertion of colonic stent(s)
C2712583|ICD9CM|AB|46.86|Endo insrt colonic stent
C2712584|ICD9CM|PT|46.87|Other insertion of colonic stent(s)
C2712584|ICD9CM|AB|46.87|Insert colonic stent NEC
C2712585|ICD9CM|PT|80.00|Arthrotomy for removal of prosthesis without replacement, unspecified site
C2712585|ICD9CM|AB|80.00|Arth/pros rem wo rep NOS
C2712586|ICD9CM|PT|80.01|Arthrotomy for removal of prosthesis without replacement, shoulder
C2712586|ICD9CM|AB|80.01|Arth/pros rem wo re-shld
C2712587|ICD9CM|PT|80.02|Arthrotomy for removal of prosthesis without replacement, elbow
C2712587|ICD9CM|AB|80.02|Arth/pros rem wo rep-elb
C2712588|ICD9CM|PT|80.03|Arthrotomy for removal of prosthesis without replacement, wrist
C2712588|ICD9CM|AB|80.03|Arth/pros rem wo re-wrst
C2712589|ICD9CM|PT|80.04|Arthrotomy for removal of prosthesis without replacement, hand and finger
C2712589|ICD9CM|AB|80.04|Arth/pros rem wo rep-hnd
C2712590|ICD9CM|PT|80.05|Arthrotomy for removal of prosthesis without replacement, hip
C2712590|ICD9CM|AB|80.05|Arth/pros rem wo rep-hip
C2712591|ICD9CM|PT|80.06|Arthrotomy for removal of prosthesis without replacement, knee
C2712591|ICD9CM|AB|80.06|Arth/pros rem wo re-knee
C2712592|ICD9CM|PT|80.07|Arthrotomy for removal of prosthesis without replacement, ankle
C2712592|ICD9CM|AB|80.07|Arth/pros rem wo rep-ank
C2712593|ICD9CM|PT|80.08|Arthrotomy for removal of prosthesis without replacement, foot and toe
C2712593|ICD9CM|AB|80.08|Arth/pros rem wo re-foot
C2712594|ICD9CM|PT|80.09|Arthrotomy for removal of prosthesis without replacement, other specified sites
C2712594|ICD9CM|AB|80.09|Arth/pros rem wo rep NEC
C2712603|ICD9CM|HT|E010|Activity involving other muscle strengthening exercises
C2712604|ICD9CM|HT|E029|Other activity
C2712604|ICD9CM|PT|E029.9|Other activity
C2712604|ICD9CM|AB|E029.9|Activity NEC
C2712605|ICD9CM|PT|041.3|Friedländer's bacillus infection in conditions classified elsewhere and of unspecified site
C2712605|ICD9CM|AB|041.3|Klebsiella pneumoniae
C2712614|ICD9CM|HT|E011|Activities involving computer technology and electronic devices
C2712615|ICD9CM|HT|670.3|Puerperal septic thrombophlebitis
C2712619|ICD9CM|PT|453.41|Acute venous embolism and thrombosis of deep vessels of proximal lower extremity
C2712619|ICD9CM|AB|453.41|Ac DVT/emb prox low ext
C2712624|ICD9CM|HT|E012|Activities involving arts and handcrafts
C2712629|ICD9CM|PT|453.40|Acute venous embolism and thrombosis of unspecified deep vessels of lower extremity
C2712629|ICD9CM|AB|453.40|Ac DVT/embl low ext NOS
C2712631|ICD9CM|PT|453.42|Acute venous embolism and thrombosis of deep vessels of distal lower extremity
C2712631|ICD9CM|AB|453.42|Ac DVT/emb distl low ext
C2712636|ICD9CM|HT|E013|Activities involving personal hygiene and household maintenance
C2712637|ICD9CM|PT|639.3|Kidney failure following abortion and ectopic and molar pregnancies
C2712637|ICD9CM|AB|639.3|Postabort kidney failure
C2712640|ICD9CM|HT|050-059.99|VIRAL DISEASES GENERALLY ACCOMPANIED BY EXANTHEM
C2712643|ICD9CM|HT|E014|Activities involving person providing caregiving
C2712644|ICD9CM|PT|V87.45|Personal history of systemic steroid therapy
C2712644|ICD9CM|AB|V87.45|Hx systemc steroid thrpy
C2712646|ICD9CM|PT|285.3|Antineoplastic chemotherapy induced anemia
C2712646|ICD9CM|AB|285.3|Anemia d/t antineo chemo
C2712648|ICD9CM|HT|E015|Activities involving food preparation, cooking and grilling
C2712654|ICD9CM|HT|17.5|Additional cardiovascular procedures
C2712655|ICD9CM|HT|E016|Activities involving property and land maintenance, building and construction
C2712660|ICD9CM|HT|17.6|Laser interstitial thermal therapy [LITT] under guidance
C2712664|ICD9CM|HT|E017|Activities involving roller coasters and other types of external motion
C2712670|ICD9CM|HT|17.7|Other diagnostic and therapeutic procedures
C2712671|ICD9CM|HT|27.5|Plastic repair of lip and mouth
C2712672|ICD9CM|PT|209.31|Merkel cell carcinoma of the face
C2712672|ICD9CM|AB|209.31|Merkel cell ca-face
C2712690|ICD9CM|HT|39.7|Endovascular procedures on vessel(s)
C2712692|ICD9CM|PT|209.32|Merkel cell carcinoma of the scalp and neck
C2712692|ICD9CM|AB|209.32|Merkel cell ca-sclp/neck
C2712697|ICD9CM|HT|E006|Activities involving other sports and athletics played individually
C2712704|ICD9CM|PT|453.87|Acute venous embolism and thrombosis of other thoracic veins
C2712704|ICD9CM|AB|453.87|Ac embl thorac vein NEC
C2712707|ICD9CM|HT|784.4|Voice and resonance disorders
C2712708|ICD9CM|HT|E007|Activities involving other sports and athletics played as a team or group
C2712711|ICD9CM|PT|621.34|Benign endometrial hyperplasia
C2712711|ICD9CM|AB|621.34|Ben endomet hyperplasia
C2712719|ICD9CM|HT|E008|Activities involving other specified sports and athletics
C2712724|ICD9CM|PT|E000.2|Volunteer activity
C2712724|ICD9CM|AB|E000.2|Volunteer activity
C2712728|ICD9CM|PT|209.35|Merkel cell carcinoma of the trunk
C2712728|ICD9CM|AB|209.35|Merkel cell ca-trunk
C2712730|ICD9CM|HT|E009|Activity involving other cardiorespiratory exercise
C2712731|ICD9CM|HT|V10.9|Other and unspecified personal history of malignant neoplasm
C2712734|ICD9CM|PT|209.36|Merkel cell carcinoma of other sites
C2712734|ICD9CM|AB|209.36|Merkel cell ca-oth sites
C2712736|MTH|PN|NOCODE|Acute venous embolism and thrombosis of other specified veins NEC in ICD9CM
C2712736|ICD9CM|AB|453.89|Ac embolism veins NEC
C2712736|ICD9CM|PT|453.89|Acute venous embolism and thrombosis of other specified veins
C2712745|ICD9CM|PT|584.7|Acute kidney failure with lesion of renal medullary [papillary] necrosis
C2712745|ICD9CM|AB|584.7|Ac kidny fail, medu necr
C2712749|ICD9CM|PT|209.70|Secondary neuroendocrine tumor, unspecified site
C2712749|ICD9CM|AB|209.70|Sec neuroendo tumor NOS
C2712755|ICD9CM|PT|453.75|Chronic venous embolism and thrombosis of subclavian veins
C2712755|ICD9CM|AB|453.75|Ch emblsm subclav veins
C2712761|ICD9CM|HT|359.7|Inflammatory and immune myopathies, NEC
C2712765|ICD9CM|PT|453.76|Chronic venous embolism and thrombosis of internal jugular veins
C2712765|ICD9CM|AB|453.76|Ch embl internl jug vein
C2712771|ICD9CM|PT|V10.91|Personal history of malignant neuroendocrine tumor
C2712771|ICD9CM|AB|V10.91|Hx malig neuroendo tumor
C2712777|ICD9CM|AB|372.06|Ac chem conjunctivitis
C2712777|ICD9CM|PT|372.06|Acute chemical conjunctivitis
C2712794|ICD9CM|PT|453.77|Chronic venous embolism and thrombosis of other thoracic veins
C2712794|ICD9CM|AB|453.77|Ch embl thorac vein NEC
C2712796|ICD9CM|PT|209.79|Secondary neuroendocrine tumor of other sites
C2712796|ICD9CM|AB|209.79|Sec neuroend tu oth site
C2712802|ICD9CM|AB|V53.59|Fit/adjust gi app-device
C2712802|ICD9CM|HT|V53.5|Fitting and adjustment of other gastrointestinal appliance and device
C2712802|ICD9CM|PT|V53.59|Fitting and adjustment of other gastrointestinal appliance and device
C2712807|ICD9CM|HT|E001|Activities involving walking and running
C2712808|ICD9CM|PT|359.79|Other inflammatory and immune myopathies, NEC
C2712808|ICD9CM|AB|359.79|Inflm/immune myopath NEC
C2712814|ICD9CM|PT|453.79|Chronic venous embolism and thrombosis of other specified veins
C2712814|ICD9CM|AB|453.79|Ch emblsm veins NEC
C2712815|ICD9CM|PT|453.50|Chronic venous embolism and thrombosis of unspecified deep vessels of lower extremity
C2712815|ICD9CM|AB|453.50|Ch DVT/embl low ext NOS
C2712816|ICD9CM|HT|E002|Activities involving water and water craft
C2712817|ICD9CM|PT|453.52|Chronic venous embolism and thrombosis of deep vessels of distal lower extremity
C2712817|ICD9CM|AB|453.52|Ch DVT/embl dstl low ext
C2712822|ICD9CM|PT|453.81|Acute venous embolism and thrombosis of superficial veins of upper extremity
C2712822|ICD9CM|AB|453.81|Ac embl suprfcl up ext
C2712828|ICD9CM|PT|453.51|Chronic venous embolism and thrombosis of deep vessels of proximal lower extremity
C2712828|ICD9CM|AB|453.51|Ch DVT/embl prox low ext
C2712831|ICD9CM|HT|E003|Activities involving ice and snow
C2712834|ICD9CM|PT|453.82|Acute venous embolism and thrombosis of deep veins of upper extremity
C2712834|ICD9CM|AB|453.82|Ac DVT/embl up ext
C2712843|ICD9CM|PT|453.2|Other venous embolism and thrombosis of inferior vena cava
C2712843|ICD9CM|AB|453.2|Oth inf vena cava thromb
C2712844|ICD9CM|HT|E004|Activities involving climbing, rappelling and jumping off
C2712845|ICD9CM|PT|453.83|Acute venous embolism and thrombosis of upper extremity, unspecified
C2712845|ICD9CM|AB|453.83|Ac emblsm up ext NOS
C2712847|ICD9CM|PT|453.85|Acute venous embolism and thrombosis of subclavian veins
C2712847|ICD9CM|AB|453.85|Ac embl subclav veins
C2712851|ICD9CM|HT|669.3|Acute kidney failure following labor and delivery
C2712854|ICD9CM|HT|E005|Activities involving dancing and other rhythmic movement
C2712855|ICD9CM|PT|453.84|Acute venous embolism and thrombosis of axillary veins
C2712855|ICD9CM|AB|453.84|Ac emblsm axillary veins
C2712857|ICD9CM|HT|V20.3|Newborn health supervision
C2712858|ICD9CM|PT|453.86|Acute venous embolism and thrombosis of internal jugular veins
C2712858|ICD9CM|AB|453.86|Ac embl internl jug vein
C2712859|ICD9CM|HT|453.4|Acute venous embolism and thrombosis of deep vessels of lower extremity
C2712860|ICD9CM|PT|569.79|Other complications of intestinal pouch
C2712860|ICD9CM|AB|569.79|Comp intest pouch NEC
C2712872|ICD9CM|HT|453.5|Chronic venous embolism and thrombosis of deep vessels of lower extremity
C2712873|ICD9CM|PT|209.71|Secondary neuroendocrine tumor of distant lymph nodes
C2712873|ICD9CM|AB|209.71|Sec neuroend tu dist lym
C2712881|ICD9CM|HT|488.0|Influenza due to identified avian influenza virus
C2712884|ICD9CM|PT|453.6|Venous embolism and thrombosis of superficial vessels of lower extremity
C2712884|ICD9CM|AB|453.6|Embl suprfcl ves low ext
C2712885|ICD9CM|PT|209.72|Secondary neuroendocrine tumor of liver
C2712885|ICD9CM|AB|209.72|Sec neuroend tumor-liver
C2712886|ICD9CM|PT|274.02|Chronic gouty arthropathy without mention of tophus (tophi)
C2712886|ICD9CM|AB|274.02|Chr gouty atrph wo tophi
C2712887|MTH|PN|NOCODE|Brain conditions NEC in ICD9CM
C2712887|ICD9CM|PT|348.89|Other conditions of brain
C2712887|ICD9CM|AB|348.89|Brain conditions NEC
C2712896|ICD9CM|HT|453.7|Chronic venous embolism and thrombosis of other specified vessels
C2712897|ICD9CM|AB|209.73|Sec neuroendo tumor-bone
C2712897|ICD9CM|PT|209.73|Secondary neuroendocrine tumor of bone
C2712898|ICD9CM|HT|E000|External cause status
C2712898|ICD9CM|HT|E000-E000.9|EXTERNAL CAUSE STATUS
C2712899|ICD9CM|PT|274.03|Chronic gouty arthropathy with tophus (tophi)
C2712899|ICD9CM|AB|274.03|Chr gouty atroph w tophi
C2712902|ICD9CM|HT|670.8|Other major puerperal infection
C2712904|ICD9CM|PT|209.74|Secondary neuroendocrine tumor of peritoneum
C2712904|ICD9CM|AB|209.74|Sec neuroendo tu-periton
C2712911|ICD9CM|PT|239.81|Neoplasms of unspecified nature, retina and choroid
C2712911|ICD9CM|AB|239.81|Neo retina/choroid NOS
C2712917|ICD9CM|HT|209.7|Secondary neuroendocrine tumors
C2712933|ICD9CM|PT|209.75|Secondary Merkel cell carcinoma
C2712933|ICD9CM|AB|209.75|Secondary Merkel cell ca
C2712938|ICD9CM|PT|453.71|Chronic venous embolism and thrombosis of superficial veins of upper extremity
C2712938|ICD9CM|AB|453.71|Ch emblsm suprfcl up ext
C2712941|ICD9CM|HT|779.3|Disorder of stomach function and feeding problems in newborn
C2712943|ICD9CM|HT|E018|Activities involving playing musical instrument
C2712948|ICD9CM|PT|453.72|Chronic venous embolism and thrombosis of deep veins of upper extremity
C2712948|ICD9CM|AB|453.72|Ch DVT/embl up ext
C2712952|ICD9CM|HT|E019|Activities involving animal care
C2712953|ICD9CM|PT|453.74|Chronic venous embolism and thrombosis of axillary veins
C2712953|ICD9CM|AB|453.74|Ch emblsm axillary veins
C2712966|ICD9CM|PT|453.73|Chronic venous embolism and thrombosis of upper extremity, unspecified
C2712966|ICD9CM|AB|453.73|Ch emblsm up ext NOS
C2712967|ICD9CM|HT|569.7|Complications of intestinal pouch
C2712970|ICD9CM|HT|488|Influenza due to certain identified influenza viruses
C2712977|ICD9CM|PT|584.5|Acute kidney failure with lesion of tubular necrosis
C2712977|ICD9CM|AB|584.5|Ac kidny fail, tubr necr
C2712983|ICD9CM|PT|584.6|Acute kidney failure with lesion of renal cortical necrosis
C2712983|ICD9CM|AB|584.6|Ac kidny fail, cort necr
C2712987|ICD9CM|AB|348.81|Temporal sclerosis
C2712987|ICD9CM|PT|348.81|Temporal sclerosis
C2712988|ICD9CM|PT|584.8|Acute kidney failure with other specified pathological lesion in kidney
C2712988|ICD9CM|AB|584.8|Acute kidney failure NEC
C2712992|ICD9CM|AB|E013.2|Vacuuming
C2712992|ICD9CM|PT|E013.2|Activities involving vacuuming
C2712994|ICD9CM|PT|E005.4|Activities involving cheerleading
C2712994|ICD9CM|AB|E005.4|Cheerleading
C2712996|ICD9CM|HT|453.8|Acute venous embolism and thrombosis of other specified veins
C2712997|MTH|PN|NOCODE|Encounter due to other specified housing or economic circumstances NEC in ICD9CM
C2712997|ICD9CM|PT|V60.89|Other specified housing or economic circumstances
C2712997|ICD9CM|AB|V60.89|Housing/econo circum NEC
C2712998|ICD9CM|HT|V45.0|Cardiac pacemaker in situ
C2713000|ICD9CM|AB|E013.3|Ironing
C2713000|ICD9CM|PT|E013.3|Activities involving ironing
C2713001|ICD9CM|PT|V57.3|Care involving speech-language therapy
C2713001|ICD9CM|AB|V57.3|Speech-language therapy
C2717961|ICD9CM|PT|446.6|Thrombotic microangiopathy
C2717961|ICD9CM|AB|446.6|Thrombot microangiopathy
C2720437|ICD9CM|HT|832|Dislocation of elbow
C2732218|MTH|PN|NOCODE|Other operations on esophagus NEC in ICD9CM
C2732218|ICD9CM|PT|42.99|Other operations on esophagus
C2732218|ICD9CM|AB|42.99|Esophageal operation NEC
C2732748|ICD9CM|PT|428.21|Acute systolic heart failure
C2732748|ICD9CM|AB|428.21|Ac systolic hrt failure
C2732749|ICD9CM|PT|428.33|Acute on chronic diastolic heart failure
C2732749|ICD9CM|AB|428.33|Ac on chr diast hrt fail
C2732951|ICD9CM|PT|428.31|Acute diastolic heart failure
C2732951|ICD9CM|AB|428.31|Ac diastolic hrt failure
C2733492|ICD9CM|PT|428.23|Acute on chronic systolic heart failure
C2733492|ICD9CM|AB|428.23|Ac on chr syst hrt fail
C2733620|MTH|PN|NOCODE|Lung operation NEC in ICD9CM
C2733620|ICD9CM|PT|33.99|Other operations on lung
C2733620|ICD9CM|AB|33.99|Lung operation NEC
C2733621|MTH|PN|NOCODE|Renal operation NEC in ICD9CM
C2733621|ICD9CM|PT|55.99|Other operations on kidney
C2733621|ICD9CM|AB|55.99|Renal operation NEC
C2733633|MTH|PN|NOCODE|Other complications of puerperium, unspecified as to episode of care NEC in ICD9CM
C2733633|ICD9CM|PT|674.80|Other complications of puerperium, unspecified as to episode of care or not applicable
C2733633|ICD9CM|AB|674.80|Puerp compl NEC-unspec
C2733634|MTH|PN|NOCODE|Other complications of puerperium - postpartum NEC in ICD9CM
C2733634|ICD9CM|PT|674.84|Other complications of puerperium, postpartum condition or complication
C2733634|ICD9CM|AB|674.84|Puerp compl NEC-postpart
C2733636|ICD9CM|PT|755.8|Other specified anomalies of unspecified limb
C2733636|ICD9CM|AB|755.8|Congen limb anomaly NEC
C2733645|MTH|PN|NOCODE|Late effects of other accidents NEC in ICD9CM
C2733645|ICD9CM|PT|E929.8|Late effects of other accidents
C2733645|ICD9CM|AB|E929.8|Late eff accident NEC
C2745960|ICD9CM|PT|375.55|Obstruction of nasolacrimal duct, neonatal
C2745960|ICD9CM|AB|375.55|Neonatal nasolacrml obst
C2745961|ICD9CM|PT|197.3|Secondary malignant neoplasm of other respiratory organs
C2745961|ICD9CM|AB|197.3|Sec malig neo resp NEC
C2745963|ICD9CM|HT|716.0|Kaschin-Beck disease
C2745963|ICD9CM|PT|716.00|Kaschin-Beck disease, site unspecified
C2745963|ICD9CM|AB|716.00|Kaschin-beck dis-unspec
C2748203|ICD9CM|PT|379.27|Vitreomacular adhesion
C2748203|ICD9CM|AB|379.27|Vitreomacular adhesion
C2825161|ICD9CM|PT|V17.41|Family history of sudden cardiac death (SCD)
C2825161|ICD9CM|AB|V17.41|Fam hx sudden card death
C2830119|ICD9CM|PT|V59.02|Blood donors, stem cells
C2830119|ICD9CM|AB|V59.02|Blood donor-stem cells
C2830120|ICD9CM|AB|V59.6|Liver donor
C2830120|ICD9CM|PT|V59.6|Liver donors
C2830121|ICD9CM|PT|V59.01|Blood donors, whole blood
C2830121|ICD9CM|AB|V59.01|Blood donor-whole blood
C2830475|ICD9CM|PT|790.22|Impaired glucose tolerance test (oral)
C2830475|ICD9CM|AB|790.22|Impaired oral glucse tol
C2830555|ICD9CM|AB|795.18|Vaginl cytol smr unsatis
C2830555|ICD9CM|PT|795.18|Unsatisfactory vaginal cytology smear
C2830589|ICD9CM|PT|793.81|Mammographic microcalcification
C2830589|ICD9CM|AB|793.81|Mammographic microcalcif
C2838014|ICD9CM|PT|173.60|Unspecified malignant neoplasm of skin of upper limb, including shoulder
C2838014|ICD9CM|AB|173.60|Mal neo skin up limb NOS
C2838017|ICD9CM|PT|173.70|Unspecified malignant neoplasm of skin of lower limb, including hip
C2838017|ICD9CM|AB|173.70|Mal neo skn low limb NOS
C2845968|ICD9CM|PT|198.1|Secondary malignant neoplasm of other urinary organs
C2845968|ICD9CM|AB|198.1|Sec malig neo urin NEC
C2853895|ICD9CM|PT|200.41|Mantle cell lymphoma, lymph nodes of head, face, and neck
C2853895|ICD9CM|AB|200.41|Mantle cell lymph head
C2853896|ICD9CM|PT|200.42|Mantle cell lymphoma, intrathoracic lymph nodes
C2853896|ICD9CM|AB|200.42|Mantle cell lymph thorax
C2853897|ICD9CM|PT|200.43|Mantle cell lymphoma, intra-abdominal lymph nodes
C2853897|ICD9CM|AB|200.43|Mantle cell lymph abdom
C2853898|ICD9CM|PT|200.44|Mantle cell lymphoma, lymph nodes of axilla and upper limb
C2853898|ICD9CM|AB|200.44|Mantle cell lymph axilla
C2853899|ICD9CM|PT|200.45|Mantle cell lymphoma, lymph nodes of inguinal region and lower limb
C2853899|ICD9CM|AB|200.45|Mantle cell lymph inguin
C2853900|ICD9CM|PT|200.46|Mantle cell lymphoma, intrapelvic lymph nodes
C2853900|ICD9CM|AB|200.46|Mantle cell lymph pelvic
C2853901|ICD9CM|PT|200.48|Mantle cell lymphoma, lymph nodes of multiple sites
C2853901|ICD9CM|AB|200.48|Mantle cell lymph multip
C2869595|ICD9CM|PT|236.3|Neoplasm of uncertain behavior of other and unspecified female genital organs
C2869595|ICD9CM|AB|236.3|Unc behav neo female NEC
C2869603|ICD9CM|PT|236.6|Neoplasm of uncertain behavior of other and unspecified male genital organs
C2869603|ICD9CM|AB|236.6|Unc behav neo male NEC
C2873698|ICD9CM|PT|236.99|Neoplasm of uncertain behavior of other and unspecified urinary organs
C2873698|ICD9CM|AB|236.99|Unc behav neo urinar NEC
C2873733|ICD9CM|PT|238.8|Neoplasm of uncertain behavior of other specified sites
C2873733|ICD9CM|AB|238.8|Uncert behavior neo NEC
C2873812|ICD9CM|PT|288.09|Other neutropenia
C2873812|ICD9CM|AB|288.09|Neutropenia NEC
C2874299|ICD9CM|PT|275.09|Other disorders of iron metabolism
C2874299|ICD9CM|AB|275.09|Disord iron metablsm NEC
C2874528|ICD9CM|PT|304.13|Sedative, hypnotic or anxiolytic dependence, in remission
C2874528|ICD9CM|AB|304.13|Sed,hyp,anxiolyt dep-rem
C2874891|ICD9CM|PT|296.61|Bipolar I disorder, most recent episode (or current) mixed, mild
C2874891|ICD9CM|AB|296.61|Bipol I currnt mix-mild
C2874892|ICD9CM|PT|296.62|Bipolar I disorder, most recent episode (or current) mixed, moderate
C2874892|ICD9CM|AB|296.62|Bipol I currnt mixed-mod
C2882273|ICD9CM|HT|428.4|Combined systolic and diastolic heart failure
C2882273|ICD9CM|PT|428.40|Combined systolic and diastolic heart failure, unspecified
C2882273|ICD9CM|AB|428.40|Syst/diast hrt fail NOS
C2882274|ICD9CM|PT|428.41|Acute combined systolic and diastolic heart failure
C2882274|ICD9CM|AB|428.41|Ac syst/diastol hrt fail
C2882275|ICD9CM|PT|428.42|Chronic combined systolic and diastolic heart failure
C2882275|ICD9CM|AB|428.42|Chr syst/diastl hrt fail
C2882276|ICD9CM|PT|428.43|Acute on chronic combined systolic and diastolic heart failure
C2882276|ICD9CM|AB|428.43|Ac/chr syst/dia hrt fail
C2882703|ICD9CM|PT|440.22|Atherosclerosis of native arteries of the extremities with rest pain
C2882703|ICD9CM|AB|440.22|Ath ext ntv at w rst pn
C2886803|ICD9CM|HT|999.6|ABO incompatibility reaction due to transfusion of blood or blood products
C2887377|ICD9CM|PT|464.50|Supraglottitis unspecified, without obstruction
C2887377|ICD9CM|AB|464.50|Supraglottis w/o obs NOS
C2887385|ICD9CM|PT|488.09|Influenza due to identified avian influenza virus with other manifestations
C2887385|ICD9CM|AB|488.09|Flu dt avian manfest NEC
C2887395|ICD9CM|PT|488.19|Influenza due to identified 2009 H1N1 influenza virus with other manifestations
C2887395|ICD9CM|AB|488.19|Flu-2009 H1N1 w oth man
C2891341|ICD9CM|PT|997.69|Other amputation stump complication
C2891341|ICD9CM|AB|997.69|Amputat stump compl NEC
C2894443|ICD9CM|HT|736.2|Other acquired deformities of finger
C2894443|ICD9CM|PT|736.29|Other acquired deformities of finger
C2894443|ICD9CM|AB|736.29|Acq finger deformity NEC
C2895155|ICD9CM|PT|524.56|Non-working side interference
C2895155|ICD9CM|AB|524.56|Nonwork side interfrnce
C2903163|ICD9CM|AB|596.81|Infection of cystostomy
C2903163|ICD9CM|PT|596.81|Infection of cystostomy
C2903164|ICD9CM|PT|596.83|Other complication of cystostomy
C2903164|ICD9CM|AB|596.83|Other comp of cystostomy
C2909960|ICD9CM|PT|766.22|Prolonged gestation of infant
C2909960|ICD9CM|AB|766.22|Prolong gestation-infant
C2910076|ICD9CM|AB|777.51|Stg I nec enterocol NB
C2910076|ICD9CM|PT|777.51|Stage I necrotizing enterocolitis in newborn
C2910077|ICD9CM|AB|777.52|Stg II nec enterocol NB
C2910077|ICD9CM|PT|777.52|Stage II necrotizing enterocolitis in newborn
C2910078|ICD9CM|PT|777.53|Stage III necrotizing enterocolitis in newborn
C2910078|ICD9CM|AB|777.53|Stg III nec enterocol NB
C2910173|ICD9CM|HT|750|Other congenital anomalies of upper alimentary tract
C2910371|ICD9CM|PT|758.33|Other microdeletions
C2910371|ICD9CM|AB|758.33|Microdeletions NEC
C2910517|ICD9CM|AB|V68.09|Issue of med certif NEC
C2910517|ICD9CM|PT|V68.09|Other issue of medical certificates
C2910575|ICD9CM|PT|V74.1|Screening examination for pulmonary tuberculosis
C2910575|ICD9CM|AB|V74.1|Screening-pulmonary TB
C2910590|ICD9CM|PT|V76.52|Special screening for malignant neoplasms of small intestine
C2910590|ICD9CM|AB|V76.52|Scrn mal neo-small intes
C2910598|ICD9CM|PT|V76.45|Screening for malignant neoplasms of testis
C2910598|ICD9CM|AB|V76.45|Screen malig neop-testis
C2910600|ICD9CM|PT|V76.46|Special screening for malignant neoplasms of ovary
C2910600|ICD9CM|AB|V76.46|Screen malig neop-ovary
C2910603|ICD9CM|PT|V76.81|Special screening for malignant neoplasms of nervous system
C2910603|ICD9CM|AB|V76.81|Screen neop-nervous syst
C2910614|ICD9CM|PT|V77.91|Screening for lipoid disorders
C2910614|ICD9CM|AB|V77.91|Screen lipoid disorders
C2910630|ICD9CM|PT|V82.81|Special screening for osteoporosis
C2910630|ICD9CM|AB|V82.81|Screen - osteoporosis
C2910670|ICD9CM|PT|V64.01|Vaccination not carried out because of acute illness
C2910670|ICD9CM|AB|V64.01|No vaccin-acute illness
C2910671|ICD9CM|PT|V64.02|Vaccination not carried out because of chronic illness or condition
C2910671|ICD9CM|AB|V64.02|No vaccin-chronc illness
C2910672|ICD9CM|PT|V64.03|Vaccination not carried out because of immune compromised state
C2910672|ICD9CM|AB|V64.03|No vaccin-immune comp
C2910787|ICD9CM|PT|V50.41|Prophylactic breast removal
C2910787|ICD9CM|AB|V50.41|Prphylct orgn rmvl brst
C2910788|ICD9CM|PT|V50.42|Prophylactic ovary removal
C2910788|ICD9CM|AB|V50.42|Prphylct orgn rmvl ovary
C2910789|ICD9CM|PT|V50.49|Other prophylactic gland removal
C2910789|ICD9CM|AB|V50.49|Prphylct orgn rmvl other
C2910897|ICD9CM|PT|V53.51|Fitting and adjustment of gastric lap band
C2910897|ICD9CM|AB|V53.51|Fit/adj gastric lap band
C2910939|ICD9CM|PT|V56.1|Fitting and adjustment of extracorporeal dialysis catheter
C2910939|ICD9CM|AB|V56.1|Ft/adj xtrcorp dial cath
C2910940|ICD9CM|PT|V56.2|Fitting and adjustment of peritoneal dialysis catheter
C2910940|ICD9CM|AB|V56.2|Fit/adj perit dial cath
C2910943|ICD9CM|AB|V58.83|Therapeutic drug monitor
C2910943|ICD9CM|PT|V58.83|Encounter for therapeutic drug monitoring
C2910964|ICD9CM|PT|V59.72|Egg (oocyte) (ovum) donor, under age 35, designated recipient
C2910964|ICD9CM|AB|V59.72|Egg donor age <35 desig
C2910966|ICD9CM|PT|V59.74|Egg (oocyte) (ovum) donor, age 35 and over, designated recipient
C2910966|ICD9CM|AB|V59.74|Egg donor age 35+ desig
C2910967|ICD9CM|PT|V59.70|Egg (oocyte) (ovum) donor, unspecified
C2910967|ICD9CM|AB|V59.70|Egg donor NEC
C2911045|ICD9CM|PT|V85.21|Body Mass Index 25.0-25.9, adult
C2911045|ICD9CM|AB|V85.21|BMI 25.0-25.9,adult
C2911046|ICD9CM|PT|V85.22|Body Mass Index 26.0-26.9, adult
C2911046|ICD9CM|AB|V85.22|BMI 26.0-26.9,adult
C2911047|ICD9CM|PT|V85.23|Body Mass Index 27.0-27.9, adult
C2911047|ICD9CM|AB|V85.23|BMI 27.0-27.9,adult
C2911048|ICD9CM|PT|V85.24|Body Mass Index 28.0-28.9, adult
C2911048|ICD9CM|AB|V85.24|BMI 28.0-28.9,adult
C2911049|ICD9CM|PT|V85.25|Body Mass Index 29.0-29.9, adult
C2911049|ICD9CM|AB|V85.25|BMI 29.0-29.9,adult
C2911051|ICD9CM|PT|V85.30|Body Mass Index 30.0-30.9, adult
C2911051|ICD9CM|AB|V85.30|BMI 30.0-30.9,adult
C2911052|ICD9CM|PT|V85.31|Body Mass Index 31.0-31.9, adult
C2911052|ICD9CM|AB|V85.31|BMI 31.0-31.9,adult
C2911053|ICD9CM|PT|V85.32|Body Mass Index 32.0-32.9, adult
C2911053|ICD9CM|AB|V85.32|BMI 32.0-32.9,adult
C2911054|ICD9CM|PT|V85.33|Body Mass Index 33.0-33.9, adult
C2911054|ICD9CM|AB|V85.33|BMI 33.0-33.9,adult
C2911055|ICD9CM|PT|V85.34|Body Mass Index 34.0-34.9, adult
C2911055|ICD9CM|AB|V85.34|BMI 34.0-34.9,adult
C2911056|ICD9CM|PT|V85.35|Body Mass Index 35.0-35.9, adult
C2911056|ICD9CM|AB|V85.35|BMI 35.0-35.9,adult
C2911057|ICD9CM|PT|V85.36|Body Mass Index 36.0-36.9, adult
C2911057|ICD9CM|AB|V85.36|BMI 36.0-36.9,adult
C2911058|ICD9CM|PT|V85.37|Body Mass Index 37.0-37.9, adult
C2911058|ICD9CM|AB|V85.37|BMI 37.0-37.9,adult
C2911059|ICD9CM|PT|V85.38|Body Mass Index 38.0-38.9, adult
C2911059|ICD9CM|AB|V85.38|BMI 38.0-38.9,adult
C2911060|ICD9CM|PT|V85.39|Body Mass Index 39.0-39.9, adult
C2911060|ICD9CM|AB|V85.39|BMI 39.0-39.9,adult
C2911062|ICD9CM|HT|V85.5|Body Mass Index, pediatric
C2911063|ICD9CM|PT|V85.51|Body Mass Index, pediatric, less than 5th percentile for age
C2911063|ICD9CM|AB|V85.51|BMI,pediatric <5%
C2911064|ICD9CM|PT|V85.52|Body Mass Index, pediatric, 5th percentile to less than 85th percentile for age
C2911064|ICD9CM|AB|V85.52|BMI,pediatric 5% - <85%
C2911065|ICD9CM|PT|V85.53|Body Mass Index, pediatric, 85th percentile to less than 95th percentile for age
C2911065|ICD9CM|AB|V85.53|BMI,pediatric 85% - <95%
C2911066|ICD9CM|PT|V85.54|Body Mass Index, pediatric, greater than or equal to 95th percentile for age
C2911066|ICD9CM|AB|V85.54|BMI,pediatric >= 95%
C2911077|ICD9CM|PT|V61.11|Counseling for victim of spousal and partner abuse
C2911077|ICD9CM|AB|V61.11|Cnsl victm partner abuse
C2911138|ICD9CM|AB|V65.11|Ped pre-brth vst-parent
C2911138|ICD9CM|PT|V65.11|Pediatric pre-birth visit for expectant parent(s)
C2911144|ICD9CM|PT|V15.86|Personal history of contact with and (suspected) exposure to lead
C2911144|ICD9CM|AB|V15.86|Hx-contact/exposure lead
C2911178|ICD9CM|AB|V58.61|Long-term use anticoagul
C2911178|ICD9CM|PT|V58.61|Long-term (current) use of anticoagulants
C2911179|ICD9CM|PT|V58.63|Long-term (current) use of antiplatelet/antithrombotic
C2911179|ICD9CM|AB|V58.63|Lng use antiplte/thrmbtc
C2911180|ICD9CM|PT|V58.64|Long-term (current) use of non-steroidal anti-inflammatories (NSAID)
C2911180|ICD9CM|AB|V58.64|Long-term anti-inflamtry
C2911181|ICD9CM|PT|V58.62|Long-term (current) use of antibiotics
C2911181|ICD9CM|AB|V58.62|Long-term use antibiotic
C2911205|ICD9CM|PT|V58.66|Long-term (current) use of aspirin
C2911205|ICD9CM|AB|V58.66|Long-term use of aspirin
C2911212|ICD9CM|PT|V16.59|Family history of malignant neoplasm of other urinary organs
C2911212|ICD9CM|AB|V16.59|Fam hx-urinry malig NEC
C2911243|ICD9CM|AB|V18.51|Family hx colonic polyps
C2911243|ICD9CM|PT|V18.51|Family history of colonic polyps
C2911244|ICD9CM|PT|V18.59|Family history of other digestive disorders
C2911244|ICD9CM|AB|V18.59|Fam hx digest disord NEC
C2911290|ICD9CM|PT|V10.59|Personal history of malignant neoplasm of other urinary organs
C2911290|ICD9CM|AB|V10.59|Hx-urinary malignan NEC
C2911331|ICD9CM|PT|V12.61|Personal history of pneumonia (recurrent)
C2911331|ICD9CM|AB|V12.61|Prsnl hx recur pneumonia
C2911483|ICD9CM|PT|V87.46|Personal history of immunosuppressive therapy
C2911483|ICD9CM|AB|V87.46|Hx immunosuppres thrpy
C2911489|ICD9CM|PT|V44.51|Cutaneous-vesicostomy
C2911489|ICD9CM|AB|V44.51|Cutaneous-vesicos status
C2911490|ICD9CM|PT|V44.52|Appendico-vesicostomy
C2911490|ICD9CM|AB|V44.52|Appendico-vesicos status
C2911491|ICD9CM|PT|V44.59|Other cystostomy
C2911491|ICD9CM|AB|V44.59|Cystostomy status NEC
C2911500|ICD9CM|PT|V45.02|Automatic implantable cardiac defibrillator in situ
C2911500|ICD9CM|AB|V45.02|Status autm crd dfbrltr
C2911565|ICD9CM|PT|V45.84|Dental restoration status
C2911565|ICD9CM|AB|V45.84|Dental restoratn status
C2911571|ICD9CM|PT|V15.21|Personal history of undergoing in utero procedure during pregnancy
C2911571|ICD9CM|AB|V15.21|Hx in utero proc in preg
C2911572|ICD9CM|PT|V15.22|Personal history of undergoing in utero procedure while a fetus
C2911572|ICD9CM|AB|V15.22|Hx in utero proc fetus
C2911643|ICD9CM|PT|V17.81|Family history of osteoporosis
C2911643|ICD9CM|AB|V17.81|Family hx osteoporosis
C2911652|ICD9CM|AB|V02.61|Hepatitis B carrier
C2911652|ICD9CM|PT|V02.61|Hepatitis B carrier
C2911654|ICD9CM|PT|V83.01|Asymptomatic hemophilia A carrier
C2911654|ICD9CM|AB|V83.01|Asympt hemoph a carrier
C2911655|ICD9CM|PT|V83.02|Symptomatic hemophilia A carrier
C2911655|ICD9CM|AB|V83.02|Sympt hemophil a carrier
C2911677|ICD9CM|PT|V07.4|Hormone replacement therapy (postmenopausal)
C2911677|ICD9CM|AB|V07.4|Hormone replace postmeno
C2919035|ICD9CM|HT|V64.0|Vaccination not carried out
C2919114|ICD9CM|HT|V86|Estrogen receptor status
C2919114|ICD9CM|HT|V86-V86.99|ESTROGEN RECEPTOR STATUS
C2919122|ICD9CM|HT|V83.0|Hemophilia A carrier
C2919132|ICD9CM|PT|V15.88|History of fall
C2919132|ICD9CM|AB|V15.88|Personal history of fall
C2919134|ICD9CM|HT|V84|Genetic susceptibility to disease
C2919460|ICD9CM|AB|719.47|Joint pain-ankle
C2919460|ICD9CM|PT|719.47|Pain in joint, ankle and foot
C2919521|ICD9CM|PT|65.23|Laparoscopic marsupialization of ovarian cyst
C2919521|ICD9CM|AB|65.23|Lap marsup ovarian cyst
C2919808|ICD9CM|PT|385.82|Cholesterin granuloma of middle ear and mastoid
C2919808|ICD9CM|AB|385.82|Cholesterin granuloma
C2921007|ICD9CM|PT|00.55|Insertion of drug-eluting stent(s) of other peripheral vessel(s)
C2921007|ICD9CM|AB|00.55|Ins d-e stent oth periph
C2921008|ICD9CM|PT|00.60|Insertion of drug-eluting stent(s) of superficial femoral artery
C2921008|ICD9CM|AB|00.60|Ins d-e stnt sup fem art
C2921010|ICD9CM|PT|17.71|Non-coronary intra-operative fluorescence vascular angiography [IFVA]
C2921010|ICD9CM|AB|17.71|Non-coronary IFVA
C2921012|ICD9CM|PT|237.79|Other neurofibromatosis
C2921012|ICD9CM|AB|237.79|Neurofibromatosis NEC
C2921014|ICD9CM|PT|275.02|Hemochromatosis due to repeated red blood cell transfusions
C2921014|ICD9CM|AB|275.02|Hemochromatos-rbc trans
C2921018|ICD9CM|PT|275.03|Other hemochromatosis
C2921018|ICD9CM|AB|275.03|Hemochromatosis NEC
C2921022|ICD9CM|PT|276.61|Transfusion associated circulatory overload
C2921022|ICD9CM|AB|276.61|Transfsn w circ overload
C2921023|ICD9CM|PT|276.69|Other fluid overload
C2921023|ICD9CM|AB|276.69|Fluid overload NEC
C2921026|ICD9CM|PT|287.49|Other secondary thrombocytopenia
C2921026|ICD9CM|AB|287.49|Sec thrombocytpenia NEC
C2921027|ICD9CM|PT|307.0|Adult onset fluency disorder
C2921027|ICD9CM|AB|307.0|Adult onset flncy disord
C2921028|ICD9CM|PT|315.35|Childhood onset fluency disorder
C2921028|ICD9CM|AB|315.35|Chldhd onset flncy disor
C2921029|ICD9CM|PT|01.20|Cranial implantation or replacement of neurostimulator pulse generator
C2921029|ICD9CM|AB|01.20|Imp/repl brain pulse gen
C2921030|ICD9CM|PT|01.29|Removal of cranial neurostimulator pulse generator
C2921030|ICD9CM|AB|01.29|Rem brain pulse generatr
C2921032|ICD9CM|PT|32.27|Bronchoscopic bronchial thermoplasty, ablation of airway smooth muscle
C2921032|ICD9CM|AB|32.27|Brnc thrmplsty,ablt mscl
C2921038|ICD9CM|PT|35.97|Percutaneous mitral valve repair with implant
C2921038|ICD9CM|AB|35.97|Perc mtrl vlv repr w imp
C2921041|ICD9CM|PT|37.34|Excision or destruction of other lesion or tissue of heart, endovascular approach
C2921041|ICD9CM|AB|37.34|Exc/des hrt les,endovasc
C2921044|ICD9CM|PT|37.37|Excision or destruction of other lesion or tissue of heart, thoracoscopic approach
C2921044|ICD9CM|AB|37.37|Exc/dest hrt les, thrspc
C2921047|ICD9CM|PT|38.97|Central venous catheter placement with guidance
C2921047|ICD9CM|AB|38.97|CV cath plcmt w guidance
C2921050|ICD9CM|AB|39.81|Imp crtd sinus stm,totl
C2921050|ICD9CM|PT|39.81|Implantation or replacement of carotid sinus stimulation device, total system
C2921051|ICD9CM|PT|39.82|Implantation or replacement of carotid sinus stimulation lead(s) only
C2921051|ICD9CM|AB|39.82|Imp/rep crtd sinus lead
C2921052|ICD9CM|PT|39.83|Implantation or replacement of carotid sinus stimulation pulse generator only
C2921052|ICD9CM|AB|39.83|Imp/rep crtd sinus gnrtr
C2921054|ICD9CM|PT|39.84|Revision of carotid sinus stimulation lead(s) only
C2921054|ICD9CM|AB|39.84|Rev crtd sinus stm leads
C2921060|ICD9CM|PT|39.85|Revision of carotid sinus stimulation pulse generator
C2921060|ICD9CM|AB|39.85|Rev crtd sinus pulse gen
C2921061|ICD9CM|PT|39.86|Removal of carotid sinus stimulation device, total system
C2921061|ICD9CM|AB|39.86|Rem crtd sinus stm, totl
C2921062|ICD9CM|PT|39.87|Removal of carotid sinus stimulation lead(s) only
C2921062|ICD9CM|AB|39.87|Rem crtd sinus stm lead
C2921063|ICD9CM|PT|39.88|Removal of carotid sinus stimulation pulse generator only
C2921063|ICD9CM|AB|39.88|Rem crtd sinus pulse gen
C2921064|ICD9CM|PT|39.89|Other operations on carotid body, carotid sinus and other vascular bodies
C2921064|ICD9CM|AB|39.89|Oth cartd body/sinus op
C2921068|ICD9CM|PT|447.70|Aortic ectasia, unspecified site
C2921068|ICD9CM|AB|447.70|Aortic ectasia, site NOS
C2921069|ICD9CM|AB|447.71|Thoracic aortic ectasia
C2921069|ICD9CM|PT|447.71|Thoracic aortic ectasia
C2921070|ICD9CM|AB|447.72|Abdominal aortic ectasia
C2921070|ICD9CM|PT|447.72|Abdominal aortic ectasia
C2921071|ICD9CM|PT|447.73|Thoracoabdominal aortic ectasia
C2921071|ICD9CM|AB|447.73|Thoracoabd aortc ectasia
C2921085|ICD9CM|PT|488.01|Influenza due to identified avian influenza virus with pneumonia
C2921085|ICD9CM|AB|488.01|Flu dt iden avian w pneu
C2921090|ICD9CM|PT|488.02|Influenza due to identified avian influenza virus with other respiratory manifestations
C2921090|ICD9CM|AB|488.02|Flu dt avian w oth resp
C2921105|ICD9CM|PT|629.81|Recurrent pregnancy loss without current pregnancy
C2921105|ICD9CM|AB|629.81|Rec preg loss wo cur prg
C2921106|ICD9CM|HT|646.3|Recurrent pregnancy loss
C2921108|ICD9CM|PT|724.02|Spinal stenosis, lumbar region, without neurogenic claudication
C2921108|ICD9CM|AB|724.02|Spin sten,lumbr wo claud
C2921109|ICD9CM|PT|724.03|Spinal stenosis, lumbar region, with neurogenic claudication
C2921109|ICD9CM|AB|724.03|Spin sten,lumbr w claud
C2921116|ICD9CM|PT|752.44|Cervical duplication
C2921116|ICD9CM|AB|752.44|Cervical duplication
C2921125|ICD9CM|PT|780.33|Post traumatic seizures
C2921125|ICD9CM|AB|780.33|Post traumatic seizures
C2921127|ICD9CM|PT|784.52|Fluency disorder in conditions classified elsewhere
C2921127|ICD9CM|AB|784.52|Flncy dsord cond elsewhr
C2921130|ICD9CM|PT|786.31|Acute idiopathic pulmonary hemorrhage in infants [AIPHI]
C2921130|ICD9CM|AB|786.31|Ac idio pul hemrg infant
C2921131|ICD9CM|PT|786.39|Other hemoptysis
C2921131|ICD9CM|AB|786.39|Hemoptysis NEC
C2921132|ICD9CM|PT|787.60|Full incontinence of feces
C2921132|ICD9CM|AB|787.60|Full incontinence-feces
C2921135|ICD9CM|HT|799.5|Signs and symptoms involving cognition
C2921136|ICD9CM|PT|799.51|Attention or concentration deficit
C2921136|ICD9CM|AB|799.51|Attn/concentrate deficit
C2921137|ICD9CM|PT|799.52|Cognitive communication deficit
C2921137|ICD9CM|AB|799.52|Cog communicate deficit
C2921138|ICD9CM|AB|799.53|Visuospatial deficit
C2921138|ICD9CM|PT|799.53|Visuospatial deficit
C2921139|ICD9CM|PT|799.54|Psychomotor deficit
C2921139|ICD9CM|AB|799.54|Psychomotor deficit
C2921140|ICD9CM|PT|799.55|Frontal lobe and executive function deficit
C2921140|ICD9CM|AB|799.55|Frontal lobe deficit
C2921141|ICD9CM|PT|799.59|Other signs and symptoms involving cognition
C2921141|ICD9CM|AB|799.59|Cognition sign/sympt NEC
C2921148|ICD9CM|PT|81.04|Dorsal and dorsolumbar fusion of the anterior column, anterior technique
C2921148|ICD9CM|AB|81.04|Drsl/drslumb fus ant/ant
C2921149|ICD9CM|PT|81.05|Dorsal and dorsolumbar fusion of the posterior column, posterior technique
C2921149|ICD9CM|AB|81.05|Drsl/dslmb fus post/post
C2921156|ICD9CM|PT|81.06|Lumbar and lumbosacral fusion of the anterior column, anterior technique
C2921156|ICD9CM|AB|81.06|Lumb/lmbosac fus ant/ant
C2921160|ICD9CM|PT|81.07|Lumbar and lumbosacral fusion of the posterior column, posterior technique
C2921160|ICD9CM|AB|81.07|Lmb/lmbsac fus post/post
C2921167|ICD9CM|PT|81.08|Lumbar and lumbosacral fusion of the anterior column, posterior technique
C2921167|ICD9CM|AB|81.08|Lumb/lmbsac fus ant/post
C2921171|ICD9CM|PT|81.36|Refusion of lumbar and lumbosacral spine, anterior column, anterior technique
C2921171|ICD9CM|AB|81.36|Refus lmb/lmbsac ant/ant
C2921177|ICD9CM|PT|81.80|Other total shoulder replacement
C2921177|ICD9CM|AB|81.80|Oth totl shouldr replace
C2921179|ICD9CM|AB|81.88|Rvrs totl shldr replacmt
C2921179|ICD9CM|PT|81.88|Reverse total shoulder replacement
C2921180|ICD9CM|PT|83.21|Open biopsy of soft tissue
C2921180|ICD9CM|AB|83.21|Open biopsy soft tissue
C2921181|ICD9CM|PT|84.94|Insertion of sternal fixation device with rigid plates
C2921181|ICD9CM|AB|84.94|Ins strn fix w rgd plate
C2921182|ICD9CM|AB|85.55|Fat graft to breast
C2921182|ICD9CM|PT|85.55|Fat graft to breast
C2921183|ICD9CM|PT|86.11|Closed biopsy of skin and subcutaneous tissue
C2921183|ICD9CM|AB|86.11|Closed bx skin/subq tiss
C2921186|ICD9CM|PT|86.87|Fat graft of skin and subcutaneous tissue
C2921186|ICD9CM|AB|86.87|Fat grft skin/subq tiss
C2921188|ICD9CM|PT|86.90|Extraction of fat for graft or banking
C2921188|ICD9CM|AB|86.90|Ext fat for grft/banking
C2921192|ICD9CM|PT|99.14|Injection or infusion of immunoglobulin
C2921192|ICD9CM|AB|99.14|Injct/inf immunoglobulin
C2921193|ICD9CM|HT|995.2|Other and unspecified adverse effect of drug, medicinal and biological substance
C2921199|ICD9CM|PT|999.60|ABO incompatibility reaction, unspecified
C2921199|ICD9CM|AB|999.60|Abo incompat react NOS
C2921202|ICD9CM|PT|999.61|ABO incompatibility with hemolytic transfusion reaction not specified as acute or delayed
C2921202|ICD9CM|AB|999.61|Abo incomp/HTR NEC
C2921204|ICD9CM|PT|999.62|ABO incompatibility with acute hemolytic transfusion reaction
C2921204|ICD9CM|AB|999.62|Abo incompat/acute HTR
C2921207|ICD9CM|PT|999.63|ABO incompatibility with delayed hemolytic transfusion reaction
C2921207|ICD9CM|AB|999.63|Abo incompat/delay HTR
C2921211|ICD9CM|PT|999.69|Other ABO incompatibility reaction
C2921211|ICD9CM|AB|999.69|Abo incompat reactn NEC
C2921214|ICD9CM|HT|999.7|Rh and other non-ABO incompatibility reaction due to transfusion of blood or blood products
C2921216|ICD9CM|PT|999.70|Rh incompatibility reaction, unspecified
C2921216|ICD9CM|AB|999.70|Rh incompat reaction NOS
C2921222|ICD9CM|PT|999.71|Rh incompatibility with hemolytic transfusion reaction not specified as acute or delayed
C2921222|ICD9CM|AB|999.71|Rh incomp/HTR NEC
C2921225|ICD9CM|PT|999.72|Rh incompatibility with acute hemolytic transfusion reaction
C2921225|ICD9CM|AB|999.72|Rh incompat/acute HTR
C2921229|ICD9CM|PT|999.73|Rh incompatibility with delayed hemolytic transfusion reaction
C2921229|ICD9CM|AB|999.73|Rh incompat/delay HTR
C2921232|ICD9CM|PT|999.74|Other Rh incompatibility reaction
C2921232|ICD9CM|AB|999.74|Rh incompat reaction NEC
C2921235|ICD9CM|PT|999.75|Non-ABO incompatibility reaction, unspecified
C2921235|ICD9CM|AB|999.75|Non-abo incomp react NOS
C2921242|ICD9CM|PT|999.76|Non-ABO incompatibility with hemolytic transfusion reaction not specified as acute or delayed
C2921242|ICD9CM|AB|999.76|Non-abo incomp/HTR NEC
C2921245|ICD9CM|PT|999.77|Non-ABO incompatibility with acute hemolytic transfusion reaction
C2921245|ICD9CM|AB|999.77|Non-abo incomp/acute HTR
C2921249|ICD9CM|PT|999.78|Non-ABO incompatibility with delayed hemolytic transfusion reaction
C2921249|ICD9CM|AB|999.78|Non-abo incomp/delay HTR
C2921252|ICD9CM|PT|999.79|Other non-ABO incompatibility reaction
C2921252|ICD9CM|AB|999.79|Non-abo incomp react NEC
C2921258|ICD9CM|PT|999.83|Hemolytic transfusion reaction, incompatibility unspecified
C2921258|ICD9CM|AB|999.83|Hemolytc trans react NOS
C2921260|ICD9CM|PT|999.84|Acute hemolytic transfusion reaction, incompatibility unspecified
C2921260|ICD9CM|AB|999.84|Acute HTR NOS
C2921262|ICD9CM|PT|999.85|Delayed hemolytic transfusion reaction, incompatibility unspecified
C2921262|ICD9CM|AB|999.85|Delayed HTR NOS
C2921265|ICD9CM|AB|E017.0|Roller coaster riding
C2921265|ICD9CM|PT|E017.0|Roller coaster riding
C2921269|ICD9CM|HT|V07|Need for isolation and other prophylactic or treatment measures
C2921270|ICD9CM|HT|V07.5|Use of agents affecting estrogen receptors and estrogen levels
C2921271|ICD9CM|PT|V07.51|Use of selective estrogen receptor modulators (SERMs)
C2921271|ICD9CM|AB|V07.51|Use of SERMs
C2921272|ICD9CM|PT|V07.8|Other specified prophylactic or treatment measure
C2921272|ICD9CM|AB|V07.8|Prophyl or tx meas NEC
C2921273|ICD9CM|PT|V11.4|Personal history of combat and operational stress reaction
C2921273|ICD9CM|AB|V11.4|Hx combat/stress reactn
C2921279|ICD9CM|PT|V13.23|Personal history of vaginal dysplasia
C2921279|ICD9CM|AB|V13.23|Hx vaginal dysplasia
C2921281|ICD9CM|PT|V13.24|Personal history of vulvar dysplasia
C2921281|ICD9CM|AB|V13.24|Hx vulvar dysplasia
C2921283|ICD9CM|HT|V13.6|Personal history of congenital (corrected) malformations
C2921284|ICD9CM|PT|V13.61|Personal history of (corrected) hypospadias
C2921284|ICD9CM|AB|V13.61|Hx-hypospadias
C2921285|ICD9CM|PT|V13.62|Personal history of other (corrected) congenital malformations of genitourinary system
C2921285|ICD9CM|AB|V13.62|Hx-cong malform-gu
C2921286|ICD9CM|PT|V13.63|Personal history of (corrected) congenital malformations of nervous system
C2921286|ICD9CM|AB|V13.63|Hx-cong malform-nervous
C2921288|ICD9CM|PT|V13.64|Personal history of (corrected) congenital malformations of eye, ear, face and neck
C2921288|ICD9CM|AB|V13.64|Hx-cong malform-eye,face
C2921289|ICD9CM|PT|V13.65|Personal history of (corrected) congenital malformations of heart and circulatory system
C2921289|ICD9CM|AB|V13.65|Hx-cong malform-heart
C2921290|ICD9CM|PT|V13.66|Personal history of (corrected) congenital malformations of respiratory system
C2921290|ICD9CM|AB|V13.66|Hx-cong malform-resp sys
C2921291|ICD9CM|PT|V13.67|Personal history of (corrected) congenital malformations of digestive system
C2921291|ICD9CM|AB|V13.67|Hx-cong malform-digest
C2921292|ICD9CM|PT|V13.68|Personal history of (corrected) congenital malformations of integument, limbs, and musculoskeletal systems
C2921292|ICD9CM|AB|V13.68|Hx-cong malform-skin,ms
C2921301|ICD9CM|PT|V15.53|Personal history of retained foreign body fully removed
C2921301|ICD9CM|AB|V15.53|Hx retained FB, rem
C2921302|ICD9CM|HT|V25.1|Encounter for insertion or removal of intrauterine contraceptive device
C2921303|ICD9CM|PT|V25.12|Encounter for removal of intrauterine contraceptive device
C2921303|ICD9CM|AB|V25.12|Removal of iud
C2921304|ICD9CM|PT|V25.13|Encounter for removal and reinsertion of intrauterine contraceptive device
C2921304|ICD9CM|AB|V25.13|Remove/insert iud
C2921306|ICD9CM|PT|V26.35|Encounter for testing of male partner of female with recurrent pregnancy loss
C2921306|ICD9CM|AB|V26.35|Test male/fem preg loss
C2921308|ICD9CM|PT|V49.87|Physical restraints status
C2921308|ICD9CM|AB|V49.87|Physical restrain status
C2921311|ICD9CM|HT|V76.1|Screening examination for malignant neoplasms of the breast
C2921312|ICD9CM|PT|V85.41|Body Mass Index 40.0-44.9, adult
C2921312|ICD9CM|AB|V85.41|BMI 40.0-44.9, adult
C2921313|ICD9CM|PT|V85.42|Body Mass Index 45.0-49.9, adult
C2921313|ICD9CM|AB|V85.42|BMI 45.0-49.9, adult
C2921314|ICD9CM|PT|V85.43|Body Mass Index 50.0-59.9, adult
C2921314|ICD9CM|AB|V85.43|BMI 50.0-59.9, adult
C2921315|ICD9CM|PT|V85.44|Body Mass Index 60.0-69.9, adult
C2921315|ICD9CM|AB|V85.44|BMI 60.0-69.9, adult
C2921316|ICD9CM|PT|V85.45|Body Mass Index 70 and over, adult
C2921316|ICD9CM|AB|V85.45|BMI 70 and over, adult
C2921317|ICD9CM|PT|V88.11|Acquired total absence of pancreas
C2921317|ICD9CM|AB|V88.11|Acq total absnc pancreas
C2921318|ICD9CM|PT|V88.12|Acquired partial absence of pancreas
C2921318|ICD9CM|AB|V88.12|Acq part absnce pancreas
C2921322|ICD9CM|HT|V90.0|Retained radioactive fragment
C2921323|ICD9CM|PT|V90.01|Retained depleted uranium fragments
C2921323|ICD9CM|AB|V90.01|Retain deplete uran frag
C2921325|ICD9CM|PT|V90.09|Other retained radioactive fragments
C2921325|ICD9CM|AB|V90.09|Retain radioac frag NEC
C2921327|ICD9CM|PT|V90.10|Retained metal fragments, unspecified
C2921327|ICD9CM|HT|V90.1|Retained metal fragments
C2921327|ICD9CM|AB|V90.10|Retained metal frag NOS
C2921328|ICD9CM|PT|V90.11|Retained magnetic metal fragments
C2921328|ICD9CM|AB|V90.11|Retain magnet metal frag
C2921329|ICD9CM|PT|V90.12|Retained nonmagnetic metal fragments
C2921329|ICD9CM|AB|V90.12|Retain nonmag meta frag
C2921333|ICD9CM|PT|V90.2|Retained plastic fragments
C2921333|ICD9CM|AB|V90.2|Retain plastic fragments
C2921334|ICD9CM|HT|V90.3|Retained organic fragments
C2921335|ICD9CM|PT|V90.31|Retained animal quills or spines
C2921335|ICD9CM|AB|V90.31|Retained quills/spines
C2921337|ICD9CM|PT|V90.33|Retained wood fragments
C2921337|ICD9CM|AB|V90.33|Retained wood fragments
C2921338|ICD9CM|PT|V90.39|Other retained organic fragments
C2921338|ICD9CM|AB|V90.39|Retain organic frag NEC
C2921339|ICD9CM|HT|V90.8|Other specified retained foreign body
C2921339|ICD9CM|PT|V90.89|Other specified retained foreign body
C2921339|ICD9CM|AB|V90.89|Retain FB NEC
C2921340|ICD9CM|AB|V90.81|Retained glass fragments
C2921340|ICD9CM|PT|V90.81|Retained glass fragments
C2921342|ICD9CM|PT|V90.83|Retained stone or crystalline fragments
C2921342|ICD9CM|AB|V90.83|Retain stone/crystl frag
C2921343|ICD9CM|PT|V90.9|Retained foreign body, unspecified material
C2921343|ICD9CM|AB|V90.9|Retain FB, mat NOS
C2921344|ICD9CM|HT|V91-V91.99|MULTIPLE GESTATION PLACENTA STATUS
C2921344|ICD9CM|HT|V91|Multiple gestation placenta status
C2921345|ICD9CM|HT|V91.0|Twin gestation placenta status
C2921346|ICD9CM|PT|V91.00|Twin gestation, unspecified number of placenta, unspecified number of amniotic sacs
C2921346|ICD9CM|AB|V91.00|Twin gest-plac/sac NOS
C2921347|ICD9CM|PT|V91.01|Twin gestation, monochorionic/monoamniotic (one placenta, one amniotic sac)
C2921347|ICD9CM|AB|V91.01|Twin gest-monochr/monoam
C2921348|ICD9CM|PT|V91.02|Twin gestation, monochorionic/diamniotic (one placenta, two amniotic sacs)
C2921348|ICD9CM|AB|V91.02|Twin gest-monochr/diamni
C2921349|ICD9CM|PT|V91.03|Twin gestation, dichorionic/diamniotic (two placentae, two amniotic sacs)
C2921349|ICD9CM|AB|V91.03|Twin gest-dich/diamniotc
C2921350|ICD9CM|PT|V91.09|Twin gestation, unable to determine number of placenta and number of amniotic sacs
C2921350|ICD9CM|AB|V91.09|Twin gest-plac/sac undet
C2921351|ICD9CM|HT|V91.1|Triplet gestation placenta status
C2921352|ICD9CM|PT|V91.10|Triplet gestation, unspecified number of placenta and unspecified number of amniotic sacs
C2921352|ICD9CM|AB|V91.10|Tripl gest-plac/sac NOS
C2921353|ICD9CM|PT|V91.11|Triplet gestation, with two or more monochorionic fetuses
C2921353|ICD9CM|AB|V91.11|Triplet gest 2+ monochor
C2921354|ICD9CM|AB|V91.12|Triplet gest 2+ monoamn
C2921354|ICD9CM|PT|V91.12|Triplet gestation, with two or more monoamniotic fetuses
C2921355|ICD9CM|AB|V91.19|Tripl gest-plac/sac und
C2921355|ICD9CM|PT|V91.19|Triplet gestation, unable to determine number of placenta and number of amniotic sacs
C2921356|ICD9CM|HT|V91.2|Quadruplet gestation placenta status
C2921357|ICD9CM|PT|V91.20|Quadruplet gestation, unspecified number of placenta and unspecified number of amniotic sacs
C2921357|ICD9CM|AB|V91.20|Quad gest-plac/sac NOS
C2921358|ICD9CM|AB|V91.21|Quad gest 2+ monochorion
C2921358|ICD9CM|PT|V91.21|Quadruplet gestation, with two or more monochorionic fetuses
C2921359|ICD9CM|PT|V91.22|Quadruplet gestation, with two or more monoamniotic fetuses
C2921359|ICD9CM|AB|V91.22|Quad gest 2+ monoamniotc
C2921360|ICD9CM|AB|V91.29|Quad gest-plac/sac undet
C2921360|ICD9CM|PT|V91.29|Quadruplet gestation, unable to determine number of placenta and number of amniotic sacs
C2921361|ICD9CM|HT|V91.9|Other specified multiple gestation placenta status
C2921363|ICD9CM|PT|V91.90|Other specified multiple gestation, unspecified number of placenta and unspecified number of amniotic sacs
C2921363|ICD9CM|AB|V91.90|Mult gest-plac/sac NOS
C2921364|ICD9CM|PT|V91.91|Other specified multiple gestation, with two or more monochorionic fetuses
C2921364|ICD9CM|AB|V91.91|Mult gest 2+ monochr NEC
C2921365|ICD9CM|PT|V91.92|Other specified multiple gestation, with two or more monoamniotic fetuses
C2921365|ICD9CM|AB|V91.92|Mult gest 2+ monoamn NEC
C2921366|ICD9CM|PT|V91.99|Other specified multiple gestation, unable to determine number of placenta and number of amniotic sacs
C2921366|ICD9CM|AB|V91.99|Mult gest-plac/sac undet
C2921372|ICD9CM|AB|V13.02|Personal history UTI
C2921372|ICD9CM|PT|V13.02|Personal history, urinary (tract) infection
C2921392|ICD9CM|AB|V12.69|Hx resp system dis NEC
C2921392|ICD9CM|PT|V12.69|Personal history of other diseases of respiratory system
C2921393|ICD9CM|AB|V13.03|Personl hx nephrotic syn
C2921393|ICD9CM|PT|V13.03|Personal history, nephrotic syndrome
C2921394|ICD9CM|AB|V12.42|Personl hx infection CNS
C2921394|ICD9CM|PT|V12.42|Personal history of infections of the central nervous system
C2921402|ICD9CM|PT|V80.01|Special screening for traumatic brain injury
C2921402|ICD9CM|AB|V80.01|Screen-traumtc brain inj
C2921408|ICD9CM|AB|V13.52|Hx stress fracture
C2921408|ICD9CM|PT|V13.52|Personal history of stress fracture
C2931914|ICD9CM|PT|435.1|Vertebral artery syndrome
C2931914|ICD9CM|AB|435.1|Vertebral artery syndrom
C2936173|ICD9CM|AB|00.66|PTCA
C2936173|ICD9CM|PT|00.66|Percutaneous transluminal coronary angioplasty [PTCA]
C2937222|ICD9CM|PT|556.2|Ulcerative (chronic) proctitis
C2937222|ICD9CM|AB|556.2|Ulcerative proctitis
C2937264|ICD9CM|PT|364.04|Secondary iridocyclitis, noninfectious
C2937264|ICD9CM|AB|364.04|Second iritis, noninfec
C2937267|ICD9CM|HT|056.0|Rubella with neurological complications
C2937267|ICD9CM|PT|056.00|Rubella with unspecified neurological complication
C2937267|ICD9CM|AB|056.00|Rubella nerve compl NOS
C2937270|ICD9CM|AB|46.21|Temporary ileostomy
C2937270|ICD9CM|PT|46.21|Temporary ileostomy
C2937271|ICD9CM|PT|51.71|Simple suture of common bile duct
C2937271|ICD9CM|AB|51.71|Simple sut-common duct
C2937300|ICD9CM|PT|359.0|Congenital hereditary muscular dystrophy
C2937300|ICD9CM|AB|359.0|Cong hered musc dystrphy
C2937352|ICD9CM|HT|66.7|Repair of fallopian tube
C2937352|ICD9CM|AB|66.73|Salpingo-salpingostomy
C2937352|ICD9CM|PT|66.73|Salpingo-salpingostomy
C2937354|ICD9CM|PT|39.42|Revision of arteriovenous shunt for renal dialysis
C2937354|ICD9CM|AB|39.42|Revis ren dialysis shunt
C2937358|ICD9CM|AB|431|Intracerebral hemorrhage
C2937358|ICD9CM|PT|431|Intracerebral hemorrhage
C2937404|ICD9CM|PT|56.51|Formation of cutaneous uretero-ileostomy
C2937404|ICD9CM|AB|56.51|Form cutan ileoureterost
C2937421|ICD9CM|HT|600|Hyperplasia of prostate
C2937421|ICD9CM|HT|600.9|Hyperplasia of prostate, unspecified
C2939119|ICD9CM|PT|23.6|Prosthetic dental implant
C2939119|ICD9CM|AB|23.6|Prosthet dental implant
C2939130|ICD9CM|HT|040|Other bacterial diseases
C2939130|ICD9CM|HT|030-041.99|OTHER BACTERIAL DISEASES
C2939134|ICD9CM|HT|76.0|Incision of facial bone without division
C2939144|ICD9CM|PT|526.0|Developmental odontogenic cysts
C2939144|ICD9CM|AB|526.0|Devel odontogenic cysts
C2939157|ICD9CM|PT|366.12|Incipient senile cataract
C2939157|ICD9CM|AB|366.12|Incipient cataract
C2939174|ICD9CM|AB|753.16|Medullary cystic kidney
C2939174|ICD9CM|PT|753.16|Medullary cystic kidney
C2939422|ICD9CM|PT|E870.1|Accidental cut, puncture, perforation or hemorrhage during infusion or transfusion
C2939422|ICD9CM|AB|E870.1|Acc cut/hem in infusion
C2939443|ICD9CM|AB|921.3|Contusion of eyeball
C2939443|ICD9CM|PT|921.3|Contusion of eyeball
C2945558|ICD9CM|PT|131.01|Trichomonal vulvovaginitis
C2945558|ICD9CM|AB|131.01|Trichomonal vaginitis
C2945587|ICD9CM|PT|20.61|Fenestration of inner ear (initial)
C2945587|ICD9CM|AB|20.61|Inner ear fenestration
C2960109|ICD9CM|PT|20.22|Incision of petrous pyramid air cells
C2960109|ICD9CM|AB|20.22|Petrus pyram air cel inc
C2960176|ICD9CM|PT|56.82|Suture of laceration of ureter
C2960176|ICD9CM|AB|56.82|Suture ureteral lacerat
C2979879|ICD9CM|AB|E005.1|Yoga
C2979879|ICD9CM|PT|E005.1|Activities involving yoga
C2979888|ICD9CM|AB|082.3|Queensland tick typhus
C2979888|ICD9CM|PT|082.3|Queensland tick typhus
C2981140|ICD9CM|AB|365.14|Glaucoma of childhood
C2981140|ICD9CM|PT|365.14|Glaucoma of childhood
C3161036|ICD9CM|PT|041.41|Shiga toxin-producing Escherichia coli [E. coli] (STEC) O157
C3161036|ICD9CM|AB|041.41|Shiga txn-produce E.coli
C3161037|ICD9CM|PT|173.00|Unspecified malignant neoplasm of skin of lip
C3161037|ICD9CM|AB|173.00|Malig neopl skin lip NOS
C3161038|ICD9CM|PT|173.02|Squamous cell carcinoma of skin of lip
C3161038|ICD9CM|AB|173.02|Squamous cell ca skn lip
C3161039|ICD9CM|PT|173.09|Other specified malignant neoplasm of skin of lip
C3161039|ICD9CM|AB|173.09|Malig neo skin lip NEC
C3161040|ICD9CM|PT|173.10|Unspecified malignant neoplasm of eyelid, including canthus
C3161040|ICD9CM|AB|173.10|Mal neo eyelid/canth NOS
C3161041|ICD9CM|PT|173.11|Basal cell carcinoma of eyelid, including canthus
C3161041|ICD9CM|AB|173.11|Basal cell ca lid/canth
C3161042|ICD9CM|PT|173.12|Squamous cell carcinoma of eyelid, including canthus
C3161042|ICD9CM|AB|173.12|Squam cell ca lid/canth
C3161043|ICD9CM|PT|173.19|Other specified malignant neoplasm of eyelid, including canthus
C3161043|ICD9CM|AB|173.19|Mal neo eyelid/canth NEC
C3161044|ICD9CM|PT|173.20|Unspecified malignant neoplasm of skin of ear and external auditory canal
C3161044|ICD9CM|AB|173.20|Malig neo skin ear NOS
C3161045|ICD9CM|PT|173.21|Basal cell carcinoma of skin of ear and external auditory canal
C3161045|ICD9CM|AB|173.21|Basal cell ca skin ear
C3161046|ICD9CM|PT|173.22|Squamous cell carcinoma of skin of ear and external auditory canal
C3161046|ICD9CM|AB|173.22|Squam cell ca skin ear
C3161047|ICD9CM|PT|173.29|Other specified malignant neoplasm of skin of ear and external auditory canal
C3161047|ICD9CM|AB|173.29|Neo skin ear/ex canl NEC
C3161048|ICD9CM|PT|173.39|Other specified malignant neoplasm of skin of other and unspecified parts of face
C3161048|ICD9CM|AB|173.30|Mal neo skn face NEC/NOS
C3161048|ICD9CM|AB|173.39|Mal neo skn face NEC/NOS
C3161048|ICD9CM|PT|173.30|Unspecified malignant neoplasm of skin of other and unspecified parts of face
C3161049|ICD9CM|PT|173.31|Basal cell carcinoma of skin of other and unspecified parts of face
C3161049|ICD9CM|AB|173.31|Bsl cel skn face NEC/NOS
C3161050|ICD9CM|PT|173.32|Squamous cell carcinoma of skin of other and unspecified parts of face
C3161050|ICD9CM|AB|173.32|Sqm cel skn face NEC/NOS
C3161051|ICD9CM|PT|173.40|Unspecified malignant neoplasm of scalp and skin of neck
C3161051|ICD9CM|AB|173.40|Mal neo sclp/skn nck NOS
C3161052|ICD9CM|PT|173.41|Basal cell carcinoma of scalp and skin of neck
C3161052|ICD9CM|AB|173.41|Bsl cell ca scalp/skn nk
C3161053|ICD9CM|PT|173.42|Squamous cell carcinoma of scalp and skin of neck
C3161053|ICD9CM|AB|173.42|Sqam cell ca sclp/skn nk
C3161054|ICD9CM|PT|173.49|Other specified malignant neoplasm of scalp and skin of neck
C3161054|ICD9CM|AB|173.49|Mal neo sclp/skn nck NEC
C3161055|ICD9CM|PT|173.50|Unspecified malignant neoplasm of skin of trunk, except scrotum
C3161055|ICD9CM|AB|173.50|Malig neo skin trunk NOS
C3161056|ICD9CM|PT|173.51|Basal cell carcinoma of skin of trunk, except scrotum
C3161056|ICD9CM|AB|173.51|Basal cell ca skin trunk
C3161057|ICD9CM|PT|173.52|Squamous cell carcinoma of skin of trunk, except scrotum
C3161057|ICD9CM|AB|173.52|Squam cell ca skin trunk
C3161058|ICD9CM|PT|173.59|Other specified malignant neoplasm of skin of trunk, except scrotum
C3161058|ICD9CM|AB|173.59|Malig neo skin trunk NEC
C3161059|ICD9CM|PT|173.61|Basal cell carcinoma of skin of upper limb, including shoulder
C3161059|ICD9CM|AB|173.61|Basal cell ca skn up lmb
C3161060|ICD9CM|PT|173.62|Squamous cell carcinoma of skin of upper limb, including shoulder
C3161060|ICD9CM|AB|173.62|Squam cell ca skn up lmb
C3161061|ICD9CM|PT|173.69|Other specified malignant neoplasm of skin of upper limb, including shoulder
C3161061|ICD9CM|AB|173.69|Malig neo skn up lmb NEC
C3161062|ICD9CM|PT|173.71|Basal cell carcinoma of skin of lower limb, including hip
C3161062|ICD9CM|AB|173.71|Basl cell ca skn low lmb
C3161063|ICD9CM|PT|173.72|Squamous cell carcinoma of skin of lower limb, including hip
C3161063|ICD9CM|AB|173.72|Sqam cell ca skn low lmb
C3161064|ICD9CM|PT|173.79|Other specified malignant neoplasm of skin of lower limb, including hip
C3161064|ICD9CM|AB|173.79|Mal neo skin low lmb NEC
C3161065|ICD9CM|PT|173.99|Other specified malignant neoplasm of skin, site unspecified
C3161065|ICD9CM|PT|173.80|Unspecified malignant neoplasm of other specified sites of skin
C3161065|ICD9CM|AB|173.99|Oth mal neo skn site NOS
C3161065|ICD9CM|AB|173.80|Mal neo skn site NEC/NOS
C3161066|ICD9CM|PT|173.81|Basal cell carcinoma of other specified sites of skin
C3161066|ICD9CM|AB|173.81|Bsl cell ca skn site NEC
C3161067|ICD9CM|PT|173.82|Squamous cell carcinoma of other specified sites of skin
C3161067|ICD9CM|AB|173.82|Sqm cell ca skn site NEC
C3161068|ICD9CM|PT|173.89|Other specified malignant neoplasm of other specified sites of skin
C3161068|ICD9CM|AB|173.89|Oth mal neo skn site NEC
C3161069|ICD9CM|PT|173.90|Unspecified malignant neoplasm of skin, site unspecified
C3161069|ICD9CM|AB|173.90|Malig neo skin site NOS
C3161070|ICD9CM|PT|173.91|Basal cell carcinoma of skin, site unspecified
C3161070|ICD9CM|AB|173.91|Basal cell ca skin NOS
C3161071|ICD9CM|PT|173.92|Squamous cell carcinoma of skin, site unspecified
C3161071|ICD9CM|AB|173.92|Squam cell ca skin NOS
C3161073|ICD9CM|PT|284.11|Antineoplastic chemotherapy induced pancytopenia
C3161073|ICD9CM|AB|284.11|Antin chemo indcd pancyt
C3161074|ICD9CM|PT|284.12|Other drug-induced pancytopenia
C3161074|ICD9CM|AB|284.12|Oth drg indcd pancytopna
C3161075|ICD9CM|PT|284.19|Other pancytopenia
C3161075|ICD9CM|AB|284.19|Other pancytopenia
C3161076|ICD9CM|PT|286.53|Antiphospholipid antibody with hemorrhagic disorder
C3161076|ICD9CM|AB|286.53|Antiphospholipid w hemor
C3161077|ICD9CM|PT|286.59|Other hemorrhagic disorder due to intrinsic circulating anticoagulants, antibodies, or inhibitors
C3161077|ICD9CM|AB|286.59|Ot hem d/t circ anticoag
C3161078|ICD9CM|PT|294.20|Dementia, unspecified, without behavioral disturbance
C3161078|ICD9CM|AB|294.20|Demen NOS w/o behv dstrb
C3161079|ICD9CM|PT|294.21|Dementia, unspecified, with behavioral disturbance
C3161079|ICD9CM|AB|294.21|Demen NOS w behav distrb
C3161080|ICD9CM|PT|358.30|Lambert-Eaton syndrome, unspecified
C3161080|ICD9CM|AB|358.30|Lambert-Eaton synd NOS
C3161081|ICD9CM|PT|358.31|Lambert-Eaton syndrome in neoplastic disease
C3161081|ICD9CM|AB|358.31|Lambert-Eaton synd neopl
C3161082|ICD9CM|PT|358.39|Lambert-Eaton syndrome in other diseases classified elsewhere
C3161082|ICD9CM|AB|358.39|Lambert-Eaton syn ot dis
C3161083|ICD9CM|PT|365.05|Open angle with borderline findings, high risk
C3161083|ICD9CM|AB|365.05|Opn ang w brdrlne hi rsk
C3161084|ICD9CM|PT|365.06|Primary angle closure without glaucoma damage
C3161084|ICD9CM|AB|365.06|Prim angle clos w/o dmg
C3161085|ICD9CM|HT|365.7|Glaucoma stage
C3161085|ICD9CM|AB|365.70|Glaucoma stage NOS
C3161085|ICD9CM|PT|365.70|Glaucoma stage, unspecified
C3161086|ICD9CM|AB|365.71|Mild stage glaucoma
C3161086|ICD9CM|PT|365.71|Mild stage glaucoma
C3161087|ICD9CM|AB|365.72|Moderate stage glaucoma
C3161087|ICD9CM|PT|365.72|Moderate stage glaucoma
C3161088|ICD9CM|AB|365.73|Severe stage glaucoma
C3161088|ICD9CM|PT|365.73|Severe stage glaucoma
C3161089|ICD9CM|PT|365.74|Indeterminate stage glaucoma
C3161089|ICD9CM|AB|365.74|Indeterm stage glaucoma
C3161090|ICD9CM|PT|414.4|Coronary atherosclerosis due to calcified coronary lesion
C3161090|ICD9CM|AB|414.4|Cor ath d/t calc cor lsn
C3161091|ICD9CM|PT|415.13|Saddle embolus of pulmonary artery
C3161091|ICD9CM|AB|415.13|Saddle embol pulmon art
C3161092|ICD9CM|PT|444.09|Other arterial embolism and thrombosis of abdominal aorta
C3161092|ICD9CM|AB|444.09|Ot art emb/thrm abd aort
C3161093|ICD9CM|PT|488.81|Influenza due to identified novel influenza A virus with pneumonia
C3161093|ICD9CM|AB|488.81|Flu dt nvl A vrs w pneu
C3161094|ICD9CM|PT|488.82|Influenza due to identified novel influenza A virus with other respiratory manifestations
C3161094|ICD9CM|AB|488.82|Flu dt nvl A w oth resp
C3161095|ICD9CM|PT|488.89|Influenza due to identified novel influenza A virus with other manifestations
C3161095|ICD9CM|AB|488.89|Flu dt novel A w oth man
C3161096|ICD9CM|PT|508.2|Respiratory conditions due to smoke inhalation
C3161096|ICD9CM|AB|508.2|Resp cond dt smoke inhal
C3161097|ICD9CM|AB|512.2|Postoperative air leak
C3161097|ICD9CM|PT|512.2|Postoperative air leak
C3161098|ICD9CM|PT|512.82|Secondary spontaneous pneumothorax
C3161098|ICD9CM|AB|512.82|Sec spont pneumothorax
C3161099|ICD9CM|AB|512.84|Other air leak
C3161099|ICD9CM|PT|512.84|Other air leak
C3161100|ICD9CM|PT|516.30|Idiopathic interstitial pneumonia, not otherwise specified
C3161100|ICD9CM|AB|516.30|Idiopath inters pneu NOS
C3161102|ICD9CM|PT|516.32|Idiopathic non-specific interstitial pneumonitis
C3161102|ICD9CM|AB|516.32|Idio non-spec inter pneu
C3161103|ICD9CM|PT|516.35|Idiopathic lymphoid interstitial pneumonia
C3161103|ICD9CM|AB|516.35|Idiopth lym interst pneu
C3161104|ICD9CM|PT|516.5|Adult pulmonary Langerhans cell histiocytosis
C3161104|ICD9CM|AB|516.5|Adlt pul Langs cell hist
C3161105|ICD9CM|PT|516.61|Neuroendocrine cell hyperplasia of infancy
C3161105|ICD9CM|AB|516.61|Neuroend cell hyprpl inf
C3161106|ICD9CM|PT|516.62|Pulmonary interstitial glycogenosis
C3161106|ICD9CM|AB|516.62|Pulm interstitl glycogen
C3161107|ICD9CM|AB|516.63|Surfactant mutation lung
C3161107|ICD9CM|PT|516.63|Surfactant mutations of the lung
C3161108|ICD9CM|PT|516.64|Alveolar capillary dysplasia with vein misalignment
C3161108|ICD9CM|AB|516.64|Alv cap dysp w vn misaln
C3161109|ICD9CM|PT|516.69|Other interstitial lung diseases of childhood
C3161109|ICD9CM|AB|516.69|Oth intrst lung dis chld
C3161110|ICD9CM|PT|518.51|Acute respiratory failure following trauma and surgery
C3161110|ICD9CM|AB|518.51|Ac resp flr fol trma/srg
C3161111|ICD9CM|PT|518.52|Other pulmonary insufficiency, not elsewhere classified, following trauma and surgery
C3161111|ICD9CM|AB|518.52|Ot pul insuf fol trm/srg
C3161112|ICD9CM|PT|518.53|Acute and chronic respiratory failure following trauma and surgery
C3161112|ICD9CM|AB|518.53|Ac/chr rsp flr fol tr/sg
C3161113|ICD9CM|PT|539.01|Infection due to gastric band procedure
C3161113|ICD9CM|AB|539.01|Inf d/t gastrc band proc
C3161114|ICD9CM|PT|539.09|Other complications of gastric band procedure
C3161114|ICD9CM|AB|539.09|Oth cmp gastrc band proc
C3161115|ICD9CM|PT|539.81|Infection due to other bariatric procedure
C3161115|ICD9CM|AB|539.81|Inf d/t ot bariatrc proc
C3161116|ICD9CM|PT|539.89|Other complications of other bariatric procedure
C3161116|ICD9CM|AB|539.89|Ot comp ot bariatrc proc
C3161117|ICD9CM|PT|596.82|Mechanical complication of cystostomy
C3161117|ICD9CM|AB|596.82|Mech comp of cystostomy
C3161118|ICD9CM|PT|629.31|Erosion of implanted vaginal mesh and other prosthetic materials to surrounding organ or tissue
C3161118|ICD9CM|AB|629.31|Eros imp vag mesh in tis
C3161119|ICD9CM|PT|629.32|Exposure of implanted vaginal mesh and other prosthetic materials into vagina
C3161119|ICD9CM|AB|629.32|Exp imp vag mesh-vagina
C3161120|ICD9CM|PT|631.0|Inappropriate change in quantitative human chorionic gonadotropin (hCG) in early pregnancy
C3161120|ICD9CM|AB|631.0|Inapp chg hCG early preg
C3161121|ICD9CM|PT|649.81|Onset (spontaneous) of labor after 37 completed weeks of gestation but before 39 completed weeks gestation, with delivery by (planned) cesarean section, delivered, with or without mention of antepartum condition
C3161121|ICD9CM|AB|649.81|Spon labr w plan C/S-del
C3161122|ICD9CM|PT|649.82|Onset (spontaneous) of labor after 37 completed weeks of gestation but before 39 completed weeks gestation, with delivery by (planned) cesarean section, delivered, with mention of postpartum complication
C3161122|ICD9CM|AB|649.82|Lbr w plan C/S-del w p/p
C3161123|ICD9CM|PT|726.13|Partial tear of rotator cuff
C3161123|ICD9CM|AB|726.13|Partial tear rotatr cuff
C3161124|ICD9CM|PT|747.31|Pulmonary artery coarctation and atresia
C3161124|ICD9CM|AB|747.31|Pulmon art coarct/atres
C3161125|ICD9CM|PT|747.39|Other anomalies of pulmonary artery and pulmonary circulation
C3161125|ICD9CM|AB|747.39|Oth anom pul artery/circ
C3161126|ICD9CM|PT|793.19|Other nonspecific abnormal finding of lung field
C3161126|ICD9CM|AB|793.19|Ot nonsp ab fnd lung fld
C3161127|ICD9CM|HT|795.5|Nonspecific reaction to tuberculin skin test without active tuberculosis
C3161127|ICD9CM|PT|795.51|Nonspecific reaction to tuberculin skin test without active tuberculosis
C3161127|ICD9CM|AB|795.51|Nonsp rea skn test wo tb
C3161128|ICD9CM|PT|795.52|Nonspecific reaction to cell mediated immunity measurement of gamma interferon antigen response without active tuberculosis
C3161128|ICD9CM|AB|795.52|Nonsp rea gma interferon
C3161129|ICD9CM|PT|808.44|Multiple closed pelvic fractures without disruption of pelvic circle
C3161129|ICD9CM|AB|808.44|Pelv fx-cl w/o plv disrp
C3161130|ICD9CM|PT|808.54|Multiple open pelvic fractures without disruption of pelvic circle
C3161130|ICD9CM|AB|808.54|Pelv fx-opn w/o pelv dis
C3161132|ICD9CM|PT|997.32|Postprocedural aspiration pneumonia
C3161132|ICD9CM|AB|997.32|Postproc aspiration pneu
C3161133|ICD9CM|PT|997.41|Retained cholelithiasis following cholecystectomy
C3161133|ICD9CM|AB|997.41|Ret cholelh fol cholecys
C3161134|ICD9CM|PT|997.49|Other digestive system complications
C3161134|ICD9CM|AB|997.49|Oth digestv system comp
C3161135|ICD9CM|PT|998.01|Postoperative shock, cardiogenic
C3161135|ICD9CM|AB|998.01|Postop shock,cardiogenic
C3161136|ICD9CM|PT|998.09|Postoperative shock, other
C3161136|ICD9CM|AB|998.09|Postop shock, other
C3161137|ICD9CM|PT|999.32|Bloodstream infection due to central venous catheter
C3161137|ICD9CM|AB|999.32|Blood inf dt cen ven cth
C3161138|ICD9CM|PT|999.33|Local infection due to central venous catheter
C3161138|ICD9CM|AB|999.33|Lcl inf dt cen ven cth
C3161139|ICD9CM|PT|999.34|Acute infection following transfusion, infusion, or injection of blood and blood products
C3161139|ICD9CM|AB|999.34|Ac inf fol trans,inf bld
C3161140|ICD9CM|PT|999.41|Anaphylactic reaction due to administration of blood and blood products
C3161140|ICD9CM|AB|999.41|Anaphyl d/t adm bld/prod
C3161141|ICD9CM|PT|999.42|Anaphylactic reaction due to vaccination
C3161141|ICD9CM|AB|999.42|Anaphyl react d/t vaccin
C3161142|ICD9CM|PT|999.49|Anaphylactic reaction due to other serum
C3161142|ICD9CM|AB|999.49|Anaph react d/t ot serum
C3161143|ICD9CM|PT|999.51|Other serum reaction due to administration of blood and blood products
C3161143|ICD9CM|AB|999.51|Ot serum react d/t blood
C3161144|ICD9CM|PT|999.52|Other serum reaction due to vaccination
C3161144|ICD9CM|AB|999.52|Ot serum react d/t vacc
C3161145|ICD9CM|PT|V12.21|Personal history of gestational diabetes
C3161145|ICD9CM|AB|V12.21|Hx gestational diabetes
C3161146|ICD9CM|PT|V12.29|Personal history of other endocrine, metabolic, and immunity disorders
C3161146|ICD9CM|AB|V12.29|Hx-endocr/meta/immun dis
C3161147|ICD9CM|PT|V13.81|Personal history of anaphylaxis
C3161147|ICD9CM|AB|V13.81|Hx of anaphylaxis
C3161148|ICD9CM|PT|V19.19|Family history of other specified eye disorder
C3161148|ICD9CM|AB|V19.19|Family hx-eye disord NEC
C3161149|ICD9CM|PT|V23.42|Pregnancy with history of ectopic pregnancy
C3161149|ICD9CM|AB|V23.42|Preg w hx ectopic preg
C3161150|ICD9CM|PT|V23.87|Pregnancy with inconclusive fetal viability
C3161150|ICD9CM|AB|V23.87|Preg w incon fetl viabil
C3161151|ICD9CM|PT|V40.31|Wandering in diseases classified elsewhere
C3161151|ICD9CM|AB|V40.31|Wandering-dis elsewhere
C3161152|ICD9CM|PT|V40.39|Other specified behavioral problem
C3161152|ICD9CM|AB|V40.39|Oth spc behavior problem
C3161153|ICD9CM|PT|V54.82|Aftercare following explantation of joint prosthesis
C3161153|ICD9CM|AB|V54.82|Aftcr explantatn jt pros
C3161154|ICD9CM|PT|V58.68|Long term (current) use of bisphosphonates
C3161154|ICD9CM|AB|V58.68|Lng term bisphosphonates
C3161155|ICD9CM|PT|V87.02|Contact with and (suspected) exposure to uranium
C3161155|ICD9CM|AB|V87.02|Cont/susp expose uranium
C3161156|ICD9CM|PT|V88.21|Acquired absence of hip joint
C3161156|ICD9CM|AB|V88.21|Acq absence of hip joint
C3161157|ICD9CM|PT|V88.22|Acquired absence of knee joint
C3161157|ICD9CM|AB|V88.22|Acq absence knee joint
C3161158|ICD9CM|PT|V88.29|Acquired absence of other joint
C3161158|ICD9CM|AB|V88.29|Acq absence of oth joint
C3161167|ICD9CM|PT|041.42|Other specified Shiga toxin-producing Escherichia coli [E. coli] (STEC)
C3161167|ICD9CM|AB|041.42|Shga txn prod E.coli NEC
C3161170|ICD9CM|PT|041.43|Shiga toxin-producing Escherichia coli [E. coli] (STEC), unspecified
C3161170|ICD9CM|AB|041.43|Shga txn prod E.coli NOS
C3161252|ICD9CM|HT|488.8|Influenza due to novel influenza A
C3161253|ICD9CM|HT|516.6|Interstitial lung diseases of childhood
C3161254|ICD9CM|HT|539|Complications of bariatric procedures
C3161255|ICD9CM|HT|539.0|Complications of gastric band procedure
C3161256|ICD9CM|HT|539.8|Complications of other bariatric procedure
C3161257|ICD9CM|HT|629.3|Complication of implanted vaginal mesh and other prosthetic materials
C3161258|ICD9CM|HT|649.8|Onset (spontaneous) of labor after 37 completed weeks of gestation but before 39 completed weeks gestation, with delivery by (planned) cesarean section
C3161259|ICD9CM|HT|704.4|Pilar and trichilemmal cysts
C3161260|ICD9CM|HT|V88.2|Acquired absence of joint
C3161261|ICD9CM|PT|02.21|Insertion or replacement of external ventricular drain [EVD]
C3161261|ICD9CM|AB|02.21|Insert/replace EVD
C3161262|ICD9CM|PT|02.22|Intracranial ventricular shunt or anastomosis
C3161262|ICD9CM|AB|02.22|Intrcran vent shunt/anas
C3161263|ICD9CM|PT|12.67|Insertion of aqueous drainage device
C3161263|ICD9CM|AB|12.67|Insert aqueous drain dev
C3161264|ICD9CM|PT|17.53|Percutaneous atherectomy of extracranial vessel(s)
C3161264|ICD9CM|AB|17.53|Perc ather extracran vsl
C3161265|ICD9CM|PT|17.54|Percutaneous atherectomy of intracranial vessel(s)
C3161265|ICD9CM|AB|17.54|Perc ather intracran vsl
C3161266|ICD9CM|PT|17.55|Transluminal coronary atherectomy
C3161266|ICD9CM|AB|17.55|Translum cor atherectomy
C3161267|ICD9CM|PT|17.56|Atherectomy of other non-coronary vessel(s)
C3161267|ICD9CM|AB|17.56|Ather oth non-cor vessel
C3161268|ICD9CM|PT|17.81|Insertion of antimicrobial envelope
C3161268|ICD9CM|AB|17.81|Insert antimicrobial env
C3161269|ICD9CM|PT|35.05|Endovascular replacement of aortic valve
C3161269|ICD9CM|AB|35.05|Endovas repl aortc valve
C3161270|ICD9CM|PT|35.06|Transapical replacement of aortic valve
C3161270|ICD9CM|AB|35.06|Trnsapcl rep aortc valve
C3161271|ICD9CM|PT|35.07|Endovascular replacement of pulmonary valve
C3161271|ICD9CM|AB|35.07|Endovas repl pulm valve
C3161272|ICD9CM|PT|35.08|Transapical replacement of pulmonary valve
C3161272|ICD9CM|AB|35.08|Trnsapcl repl pulm valve
C3161273|ICD9CM|PT|35.09|Endovascular replacement of unspecified heart valve
C3161273|ICD9CM|AB|35.09|Endovas repl uns hrt vlv
C3161274|ICD9CM|PT|38.26|Insertion of implantable pressure sensor without lead for intracardiac or great vessel hemodynamic monitoring
C3161274|ICD9CM|AB|38.26|Insrt prsr snsr w/o lead
C3161275|ICD9CM|PT|39.77|Temporary (partial) therapeutic endovascular occlusion of vessel
C3161275|ICD9CM|AB|39.77|Temp endovsc occls vessl
C3161276|ICD9CM|PT|39.78|Endovascular implantation of branching or fenestrated graft(s) in aorta
C3161276|ICD9CM|AB|39.78|Endovas impln grft aorta
C3161277|ICD9CM|PT|43.82|Laparoscopic vertical (sleeve) gastrectomy
C3161277|ICD9CM|AB|43.82|Lap vertical gastrectomy
C3161278|ICD9CM|PT|68.24|Uterine artery embolization [UAE] with coils
C3161278|ICD9CM|AB|68.24|Uterine art emb w coils
C3161279|ICD9CM|PT|68.25|Uterine artery embolization [UAE] without coils
C3161279|ICD9CM|AB|68.25|Uterine art emb w/o coil
C3161326|ICD9CM|HT|17.8|Other adjunct procedures
C3161330|ICD9CM|PT|318.2|Profound intellectual disabilities
C3161330|ICD9CM|AB|318.2|Profnd intellct disablty
C3161331|ICD9CM|PT|319|Unspecified intellectual disabilities
C3161331|ICD9CM|AB|319|Intellect disability NOS
C3161333|ICD9CM|PT|488.11|Influenza due to identified 2009 H1N1 influenza virus with pneumonia
C3161333|ICD9CM|AB|488.11|Flu dt 2009 H1N1 w pneu
C3161334|ICD9CM|PT|488.12|Influenza due to identified 2009 H1N1 influenza virus with other respiratory manifestations
C3161334|ICD9CM|AB|488.12|Flu-2009 H1N1 w oth resp
C3161335|ICD9CM|PT|995.0|Other anaphylactic reaction
C3161335|ICD9CM|AB|995.0|Other anaphylactic react
C3161345|ICD9CM|PT|995.69|Anaphylactic reaction due to other specified food
C3161345|ICD9CM|AB|995.69|Anphyl react oth sp food
C3161349|ICD9CM|PT|00.61|Percutaneous angioplasty of extracranial vessel(s)
C3161349|ICD9CM|AB|00.61|Perc angio extracran ves
C3161350|ICD9CM|PT|35.20|Open and other replacement of unspecified heart valve
C3161350|ICD9CM|AB|35.20|Opn/oth rep hrt vlv NOS
C3161351|ICD9CM|PT|35.21|Open and other replacement of aortic valve with tissue graft
C3161351|ICD9CM|AB|35.21|Opn/oth rep aort vlv-tis
C3161352|ICD9CM|PT|35.22|Open and other replacement of aortic valve
C3161352|ICD9CM|AB|35.22|Opn/oth rep aortic valve
C3161353|ICD9CM|PT|35.23|Open and other replacement of mitral valve with tissue graft
C3161353|ICD9CM|AB|35.23|Opn/oth rep mtrl vlv-tis
C3161354|ICD9CM|PT|35.24|Open and other replacement of mitral valve
C3161354|ICD9CM|AB|35.24|Opn/oth rep mitral valve
C3161355|ICD9CM|PT|35.25|Open and other replacement of pulmonary valve with tissue graft
C3161355|ICD9CM|AB|35.25|Opn/oth rep pulm vlv-tis
C3161356|ICD9CM|PT|35.26|Open and other replacement of pulmonary valve
C3161356|ICD9CM|AB|35.26|Opn/oth repl pul valve
C3161357|ICD9CM|PT|35.27|Open and other replacement of tricuspid valve with tissue graft
C3161357|ICD9CM|AB|35.27|Opn/oth rep tcspd vlv-ts
C3161358|ICD9CM|PT|35.28|Open and other replacement of tricuspid valve
C3161358|ICD9CM|AB|35.28|Opn/oth repl tcspd valve
C3161359|ICD9CM|PT|43.89|Open and other partial gastrectomy
C3161359|ICD9CM|AB|43.89|Opn/oth part gastrectomy
C3161360|ICD9CM|PT|86.95|Insertion or replacement of multiple array neurostimulator pulse generator, not specified as rechargeable
C3161360|ICD9CM|AB|86.95|Ins/re pls gn no rechrg
C3161361|ICD9CM|PT|86.98|Insertion or replacement of multiple array (two or more) rechargeable neurostimulator pulse generator
C3161361|ICD9CM|AB|86.98|Ins/rep mul pul gn,rechg
C3161362|ICD9CM|HT|173|Other and unspecified malignant neoplasm of skin
C3161363|ICD9CM|HT|173.1|Other and unspecified malignant neoplasm of skin of eyelid, including canthus
C3161364|ICD9CM|HT|173.2|Other and unspecified malignant neoplasm of skin of ear and external auditory canal
C3161365|ICD9CM|HT|173.3|Other and unspecified malignant neoplasm of skin of other and unspecified parts of face
C3161366|ICD9CM|HT|173.4|Other and unspecified malignant neoplasm of scalp and skin of neck
C3161367|ICD9CM|HT|173.5|Other and unspecified malignant neoplasm of skin of trunk, except scrotum
C3161368|ICD9CM|HT|173.6|Other and unspecified malignant neoplasm of skin of upper limb, including shoulder
C3161369|ICD9CM|HT|173.7|Other and unspecified malignant neoplasm of skin of lower limb, including hip
C3161370|ICD9CM|HT|173.8|Other and unspecified malignant neoplasm of other specified sites of skin
C3161371|ICD9CM|HT|173.9|Other and unspecified malignant neoplasm of skin, site unspecified
C3161379|ICD9CM|HT|290-319.99|MENTAL, BEHAVIORAL AND NEURODEVELOPMENTAL DISORDERS
C3161382|ICD9CM|HT|318|Other specified intellectual disabilities
C3161395|ICD9CM|HT|35.0|Closed heart valvotomy or transcatheter replacement of heart valve
C3161396|ICD9CM|HT|35.2|Open and other replacement of heart valve
C3161430|ICD9CM|HT|488.1|Influenza due to identified 2009 H1N1 influenza virus
C3161433|ICD9CM|HT|512|Pneumothorax and air leak
C3161434|ICD9CM|HT|512.8|Other pneumothorax and air leak
C3161439|ICD9CM|HT|646.7|Liver and biliary tract disorders in pregnancy
C3161458|ICD9CM|HT|999.4|Anaphylactic reaction due to serum, not elsewhere classified
C3161460|ICD9CM|PT|973.3|Poisoning by other cathartics, including intestinal atonia
C3161460|ICD9CM|AB|973.3|Poisoning-cathartic NEC
C3162029|ICD9CM|PT|17.36|Laparoscopic sigmoidectomy
C3162029|ICD9CM|AB|17.36|Lap sigmoidectomy
C3241919|ICD9CM|PT|695.12|Erythema multiforme major
C3241919|ICD9CM|AB|695.12|Erythema multiforme maj
C3241938|ICD9CM|HT|720-724.99|DORSOPATHIES
C3243009|HL7V3.0|VS|2.16.840.1.113883.1.11.15931|DiagnosisICD9CM
C3251587|ICD9CM|PT|996.88|Complications of transplanted organ, stem cell
C3251587|ICD9CM|AB|996.88|Comp tp organ-stem cell
C3251816|ICD9CM|PT|441.2|Thoracic aneurysm without mention of rupture
C3251816|ICD9CM|AB|441.2|Thoracic aortic aneurysm
C3263686|ICD9CM|PT|12.64|Trabeculectomy ab externo
C3263686|ICD9CM|AB|12.64|Trabeculectom ab externo
C3264152|ICD9CM|PT|365.01|Open angle with borderline findings, low risk
C3264152|ICD9CM|AB|365.01|Opn angl brderln lo risk
C3278433|ICD9CM|HT|833|Dislocation of wrist
C3463824|ICD9CM|PT|238.75|Myelodysplastic syndrome, unspecified
C3463824|ICD9CM|AB|238.75|Myelodysplastic synd NOS
C3484393|ICD9CM|PT|00.95|Injection or infusion of glucarpidase
C3484393|ICD9CM|AB|00.95|Injct/infus glucarpidase
C3495405|ICD9CM|PT|85.48|Bilateral extended radical mastectomy
C3495405|ICD9CM|AB|85.48|Bil exten rad mastectomy
C3495413|ICD9CM|HT|868|Injury to other intra-abdominal organs
C3495436|ICD9CM|PT|085.4|Cutaneous leishmaniasis, American
C3495436|ICD9CM|AB|085.4|Cutan leishmanias amer
C3495439|ICD9CM|PT|611.0|Inflammatory disease of breast
C3495439|ICD9CM|AB|611.0|Inflam disease of breast
C3495540|ICD9CM|PT|520.4|Disturbances of tooth formation
C3495540|ICD9CM|AB|520.4|Tooth formation disturb
C3495604|ICD9CM|HT|440.2|Atherosclerosis of native arteries of the extremities
C3495801|ICD9CM|AB|446.4|Wegener's granulomatosis
C3495801|ICD9CM|PT|446.4|Wegener's granulomatosis
C3536714|ICD9CM|AB|753.15|Renal dysplasia
C3536714|ICD9CM|PT|753.15|Renal dysplasia
C3536892|ICD9CM|HT|391|Rheumatic fever with heart involvement
C3536895|ICD9CM|PT|757.9|Unspecified congenital anomaly of the integument
C3536895|ICD9CM|HT|757|Congenital anomalies of the integument
C3536895|ICD9CM|AB|757.9|Integument anomaly NOS
C3537055|ICD9CM|PT|685.0|Pilonidal cyst with abscess
C3537055|ICD9CM|AB|685.0|Pilonidal cyst w abscess
C3537062|ICD9CM|PT|V69.1|Inappropriate diet and eating habits
C3537062|ICD9CM|AB|V69.1|Inapprt diet eat habits
C3537063|ICD9CM|HT|674.2|Disruption of obstetrical perineal wound
C3537063|ICD9CM|PT|674.24|Disruption of perineal wound, postpartum condition or complication
C3537063|ICD9CM|AB|674.24|Disrupt perineum-postpar
C3537179|ICD9CM|AB|104.0|Nonvenereal endemic syph
C3537179|ICD9CM|PT|104.0|Nonvenereal endemic syphilis
C3542020|ICD9CM|PT|780.65|Hypothermia not associated with low environmental temperature
C3542020|ICD9CM|AB|780.65|Hypothrm-wo low env tmp
C3542501|ICD9CM|PT|357.0|Acute infective polyneuritis
C3542501|ICD9CM|AB|357.0|Ac infect polyneuritis
C3542504|ICD9CM|PT|79.32|Open reduction of fracture with internal fixation, radius and ulna
C3542504|ICD9CM|AB|79.32|Op red-int fix rad/ulna
C3543852|ICD9CM|PT|780.72|Functional quadriplegia
C3543852|ICD9CM|AB|780.72|Functional quadriplegia
C3550569|ICD9CM|PT|360.34|Flat anterior chamber of eye
C3550569|ICD9CM|AB|360.34|Flat anterior chamber
C3647143|ICD9CM|PT|198.6|Secondary malignant neoplasm of ovary
C3647143|ICD9CM|AB|198.6|Second malig neo ovary
C3648012|ICD9CM|PT|202.78|Peripheral T cell lymphoma, lymph nodes of multiple sites
C3648012|ICD9CM|AB|202.78|Periph T cell lym multip
C3648014|ICD9CM|PT|202.76|Peripheral T cell lymphoma, intrapelvic lymph nodes
C3648014|ICD9CM|AB|202.76|Periph T cell lym pelvic
C3648015|ICD9CM|PT|202.73|Peripheral T cell lymphoma, intra-abdominal lymph nodes
C3648015|ICD9CM|AB|202.73|Periph T cell lym abdom
C3648016|ICD9CM|PT|202.75|Peripheral T cell lymphoma, lymph nodes of inguinal region and lower limb
C3648016|ICD9CM|AB|202.75|Periph T cell lym inguin
C3648017|ICD9CM|PT|202.71|Peripheral T cell lymphoma, lymph nodes of head, face, and neck
C3648017|ICD9CM|AB|202.71|Periph T cell lymph head
C3648018|ICD9CM|PT|202.74|Peripheral T cell lymphoma, lymph nodes of axilla and upper limb
C3648018|ICD9CM|AB|202.74|Periph T cell lym axilla
C3648917|ICD9CM|HT|286.5|Hemorrhagic disorder due to intrinsic circulating anticoagulants, antibodies, or inhibitors
C3662039|ICD9CM|PT|333.85|Subacute dyskinesia due to drugs
C3662039|ICD9CM|AB|333.85|Subac dyskinesa d/t drug
C3662231|ICD9CM|PT|762.0|Placenta previa affecting fetus or newborn
C3662231|ICD9CM|AB|762.0|Placenta previa aff NB
C3665334|ICD9CM|PT|552.03|Femoral hernia with obstruction, bilateral, recurrent
C3665334|ICD9CM|AB|552.03|Rec bil fem hern w obstr
C3665340|ICD9CM|PT|298.0|Depressive type psychosis
C3665340|ICD9CM|AB|298.0|React depress psychosis
C3665346|ICD9CM|PT|369.9|Unspecified visual loss
C3665346|ICD9CM|AB|369.9|Visual loss NOS
C3665387|ICD9CM|PT|438.7|Late effects of cerebrovascular disease, disturbances of vision
C3665387|ICD9CM|AB|438.7|Disturbances of vision
C3665435|ICD9CM|PT|296.31|Major depressive affective disorder, recurrent episode, mild
C3665435|ICD9CM|AB|296.31|Recurr depr psychos-mild
C3665438|ICD9CM|PT|363.05|Focal retinitis and retinochoroiditis, juxtapapillary
C3665438|ICD9CM|AB|363.05|Juxtapap focal retinitis
C3665439|ICD9CM|AB|366.17|Mature cataract
C3665439|ICD9CM|PT|366.17|Total or mature cataract
C3665440|ICD9CM|PT|377.53|Disorders of optic chiasm associated with vascular disorders
C3665440|ICD9CM|AB|377.53|Opt chiasm w vascul dis
C3665441|ICD9CM|PT|377.71|Disorders of visual cortex associated with neoplasms
C3665441|ICD9CM|AB|377.71|Vis cortx dis w neoplasm
C3665442|ICD9CM|PT|377.72|Disorders of visual cortex associated with vascular disorders
C3665442|ICD9CM|AB|377.72|Vis cortx dis w vasc dis
C3665443|ICD9CM|PT|377.73|Disorders of visual cortex associated with inflammatory disorders
C3665443|ICD9CM|AB|377.73|Vis cortex dis w inflam
C3665446|ICD9CM|PT|940.4|Other burn of cornea and conjunctival sac
C3665446|ICD9CM|AB|940.4|Burn cornea/conjunct NEC
C3665447|ICD9CM|HT|946|Burns of multiple specified sites
C3665450|ICD9CM|AB|12.71|Cyclodiathermy
C3665450|ICD9CM|PT|12.71|Cyclodiathermy
C3665457|ICD9CM|PT|301.12|Chronic depressive personality disorder
C3665457|ICD9CM|AB|301.12|Chr depressive person
C3665458|ICD9CM|PT|404.91|Hypertensive heart and chronic kidney disease, unspecified, with heart failure and with chronic kidney disease stage I through stage IV, or unspecified
C3665458|ICD9CM|AB|404.91|Hyp ht/kd NOS I-IV w hf
C3665459|ICD9CM|PT|806.4|Closed fracture of lumbar spine with spinal cord injury
C3665459|ICD9CM|AB|806.4|Cl lumbar fx w cord inj
C3665466|ICD9CM|PT|112.89|Other candidiasis of other specified sites
C3665466|ICD9CM|AB|112.89|Candidiasis site NEC
C3665468|ICD9CM|PT|909.3|Late effect of complications of surgical and medical care
C3665468|ICD9CM|AB|909.3|Late eff surg/med compl
C3665469|ICD9CM|PT|07.45|Reimplantation of adrenal tissue
C3665469|ICD9CM|AB|07.45|Adrenal reimplantation
C3665497|ICD9CM|HT|305|Nondependent abuse of drugs
C3665587|ICD9CM|PT|290.0|Senile dementia, uncomplicated
C3665587|ICD9CM|AB|290.0|Senile dementia uncomp
C3665588|ICD9CM|PT|172.1|Malignant melanoma of skin of eyelid, including canthus
C3665588|ICD9CM|AB|172.1|Malig melanoma eyelid
C3665596|ICD9CM|HT|078.1|Viral warts
C3665608|ICD9CM|HT|674.1|Disruption of cesarean wound
C3665609|ICD9CM|AB|372.53|Conjunctival xerosis
C3665609|ICD9CM|PT|372.53|Conjunctival xerosis
C3665667|ICD9CM|PT|296.36|Major depressive affective disorder, recurrent episode, in full remission
C3665667|ICD9CM|AB|296.36|Recur depr psyc-full rem
C3665668|ICD9CM|HT|239|Neoplasms of unspecified nature
C3665668|ICD9CM|HT|239-239.99|NEOPLASMS OF UNSPECIFIED NATURE
C3693456|ICD9CM|PT|327.44|Parasomnia in conditions classified elsewhere
C3693456|ICD9CM|AB|327.44|Parasomnia oth diseases
C3695318|ICD9CM|HT|403|Hypertensive chronic kidney disease
C3697208|ICD9CM|PT|635.82|Legally induced abortion, with unspecified complication, complete
C3697208|ICD9CM|AB|635.82|Leg ab w compl NOS-comp
C3714535|ICD9CM|PT|524.22|Malocclusion, Angle's class II
C3714535|ICD9CM|AB|524.22|Malocc-Angle's class II
C3714542|ICD9CM|HT|200.1|Lymphosarcoma
C3714552|ICD9CM|AB|799.3|Debility NOS
C3714552|ICD9CM|PT|799.3|Debility, unspecified
C3714588|ICD9CM|PT|V23.9|Supervision of unspecified high-risk pregnancy
C3714588|ICD9CM|AB|V23.9|Suprv high-risk preg NOS
C3714726|ICD9CM|HT|85|Operations on the breast
C3714744|ICD9CM|HT|302.7|Psychosexual dysfunction
C3714744|ICD9CM|PT|302.70|Psychosexual dysfunction, unspecified
C3714744|ICD9CM|AB|302.70|Psychosexual dysfunc NOS
C3714756|ICD9CM|HT|317-319.99|INTELLECTUAL DISABILITIES
C3812410|ICD9CM|PT|362.22|Retinopathy of prematurity, stage 0
C3812410|ICD9CM|AB|362.22|Retinoph prematr,stage 0
C3812874|ICD9CM|PT|621.35|Endometrial intraepithelial neoplasia [EIN]
C3812874|ICD9CM|AB|621.35|Endomet intraepithl neop
C3812903|ICD9CM|HT|665.1|Rupture of uterus during labor
C3831782|ICD9CM|AB|380.12|Acute swimmers' ear
C3831782|ICD9CM|PT|380.12|Acute swimmers' ear
C3839935|ICD9CM|PT|368.43|Sector or arcuate visual field defects
C3839935|ICD9CM|AB|368.43|Sector or arcuate defect
C3846112|ICD9CM|HT|92.3|Stereotactic radiosurgery
C3846112|ICD9CM|PT|92.30|Stereotactic radiosurgery, not otherwise specified
C3846112|ICD9CM|AB|92.30|Stereo radiosurgery NOS
C3854304|ICD9CM|PT|753.11|Congenital single renal cyst
C3854304|ICD9CM|AB|753.11|Congenital renal cyst
C3858944|SRC|VPT|V-ICD9CM_2014|International Classification of Diseases, Ninth Revision, Clinical Modification, 2014
C3858944|SRC|VAB|V-ICD9CM_2014|ICD9CM_2014
C3858944|SRC|VSY|V-ICD9CM_2014|ICD-9-CM, 2014
C3858946|ICD9CM|PT|00.96|Infusion of 4-Factor Prothrombin Complex Concentrate
C3858946|ICD9CM|AB|00.96|Infusion 4F-PCC
C3858947|ICD9CM|HT|14.8|Implantation of epiretinal visual prosthesis
C3858947|ICD9CM|PT|14.81|Implantation of epiretinal visual prosthesis
C3858947|ICD9CM|AB|14.81|Imp epiretinal prosth
C3858948|ICD9CM|PT|14.82|Removal of epiretinal visual prosthesis
C3858948|ICD9CM|AB|14.82|Rem epiretinal prosth
C3858949|ICD9CM|PT|14.83|Revision or replacement of epiretinal visual prosthesis
C3858949|ICD9CM|AB|14.83|Rev/repl epiretinal pros
C3874311|ICD9CM|PT|569.87|Vomiting of fecal matter
C3874311|ICD9CM|AB|569.87|Vomiting of fecal matter
C3874327|ICD9CM|PT|538|Gastrointestinal mucositis (ulcerative)
C3874327|ICD9CM|AB|538|GI mucositis (ulceratve)
C3875058|ICD9CM|HT|273|Disorders of plasma protein metabolism
C3875058|ICD9CM|PT|273.9|Unspecified disorder of plasma protein metabolism
C3875058|ICD9CM|AB|273.9|Dis plas protein met NOS
C3875374|ICD9CM|PT|277.82|Carnitine deficiency due to inborn errors of metabolism
C3875374|ICD9CM|AB|277.82|Crnitne def d/t nb met
C3887558|ICD9CM|AB|288.4|Hemophagocytic syndromes
C3887558|ICD9CM|PT|288.4|Hemophagocytic syndromes
C3887597|ICD9CM|PT|727.03|Trigger finger (acquired)
C3887597|ICD9CM|AB|727.03|Trigger finger
C3887666|ICD9CM|PT|254.0|Persistent hyperplasia of thymus
C3887666|ICD9CM|AB|254.0|Persist hyperplas thymus
C3887875|ICD9CM|HT|368.4|Visual field defects
C3887875|ICD9CM|AB|368.40|Visual field defect NOS
C3887875|ICD9CM|PT|368.40|Visual field defect, unspecified
C3887878|ICD9CM|PT|245.3|Chronic fibrous thyroiditis
C3887878|ICD9CM|AB|245.3|Chr fibrous thyroiditis
C4038618|ICD9CM|PT|562.02|Diverticulosis of small intestine with hemorrhage
C4038618|ICD9CM|AB|562.02|Dvrtclo sml int w hmrhg
C4040007|ICD9CM|PT|337.21|Reflex sympathetic dystrophy of the upper limb
C4040007|ICD9CM|AB|337.21|Rflx sym dystrph up limb
C4040988|ICD9CM|PT|51.41|Common duct exploration for removal of calculus
C4040988|ICD9CM|AB|51.41|Cde for calculus remov
C4041147|ICD9CM|PT|491.21|Obstructive chronic bronchitis with (acute) exacerbation
C4041147|ICD9CM|AB|491.21|Obs chr bronc w(ac) exac
C4048158|ICD9CM|HT|780.3|Convulsions
C4049006|ICD9CM|PT|279.01|Selective IgA immunodeficiency
C4049006|ICD9CM|AB|279.01|Selective iga immunodef
C4076694|ICD9CM|PT|727.63|Nontraumatic rupture of extensor tendons of hand and wrist
C4076694|ICD9CM|AB|727.63|Rupt exten tendon hand
C4076715|ICD9CM|PT|209.33|Merkel cell carcinoma of the upper limb
C4076715|ICD9CM|AB|209.33|Merkel cell ca-up limb
C4076723|ICD9CM|PT|209.34|Merkel cell carcinoma of the lower limb
C4076723|ICD9CM|AB|209.34|Merkel cell ca-low limb
C4082244|ICD9CM|AB|738.11|Zygomatic hyperplasia
C4082244|ICD9CM|PT|738.11|Zygomatic hyperplasia
C4082762|ICD9CM|AB|110.1|Dermatophytosis of nail
C4082762|ICD9CM|PT|110.1|Dermatophytosis of nail
C4282165|ICD9CM|PT|785.6|Enlargement of lymph nodes
C4282165|ICD9CM|AB|785.6|Enlargement lymph nodes
C4317048|ICD9CM|PT|51.85|Endoscopic sphincterotomy and papillotomy
C4317048|ICD9CM|AB|51.85|Endosc sphincterotomy
C4317290|ICD9CM|PT|V69.5|Behavioral insomnia of childhood
C4317290|ICD9CM|AB|V69.5|Behav insomnia-childhood
C4520826|ICD9CM|PT|01.14|Open biopsy of brain
C4520826|ICD9CM|AB|01.14|Open brain biopsy
C4520843|ICD9CM|HT|372.4|Pterygium
C4520843|ICD9CM|AB|372.40|Pterygium NOS
C4520843|ICD9CM|PT|372.40|Pterygium, unspecified
C4520984|ICD9CM|PT|V66.6|Convalescence following combined treatment
C4520984|ICD9CM|AB|V66.6|Comb treatment convales
C4521098|ICD9CM|PT|07.12|Open biopsy of adrenal gland
C4521098|ICD9CM|AB|07.12|Open adrenal gland bx
C4551472|ICD9CM|PT|425.11|Hypertrophic obstructive cardiomyopathy
C4551472|ICD9CM|AB|425.11|Hyprtrophc obst cardiomy
C4551492|ICD9CM|AB|752.64|Micropenis
C4551492|ICD9CM|PT|752.64|Micropenis
C4551507|ICD9CM|HT|743.2|Buphthalmos
C4551507|ICD9CM|AB|743.20|Buphthalmos NOS
C4551507|ICD9CM|PT|743.20|Buphthalmos, unspecified
C4551519|ICD9CM|PT|378.54|Sixth or abducens nerve palsy
C4551519|ICD9CM|AB|378.54|Sixth nerve palsy
C4551629|ICD9CM|AB|754.62|Talipes calcaneovalgus
C4551629|ICD9CM|PT|754.62|Talipes calcaneovalgus
C4551631|ICD9CM|PT|751.62|Congenital cystic disease of liver
C4551631|ICD9CM|AB|751.62|Cong cystic liver dis
C4551633|ICD9CM|PT|362.74|Pigmentary retinal dystrophy
C4551633|ICD9CM|AB|362.74|Pigment retina dystrophy
C4551644|ICD9CM|PT|85.24|Excision of ectopic breast tissue
C4551644|ICD9CM|AB|85.24|Exc ectopic breast tissu
C4551650|ICD9CM|AB|530.3|Esophageal stricture
C4551650|ICD9CM|PT|530.3|Stricture and stenosis of esophagus
C4551691|ICD9CM|HT|598|Urethral stricture
C4551691|ICD9CM|AB|598.9|Urethral stricture NOS
C4551691|ICD9CM|PT|598.9|Urethral stricture, unspecified
C4551722|ICD9CM|AB|742.0|Encephalocele
C4551722|ICD9CM|PT|742.0|Encephalocele
C4551827|ICD9CM|PT|359.1|Hereditary progressive muscular dystrophy
C4551827|ICD9CM|AB|359.1|Hered prog musc dystrphy
C4551903|ICD9CM|PT|747.41|Total anomalous pulmonary venous connection
C4551903|ICD9CM|AB|747.41|Tot anom pulm ven connec
C4552054|ICD9CM|PT|92.02|Liver scan and radioisotope function study
C4552054|ICD9CM|AB|92.02|Liver scan/isotope funct
C4721400|ICD9CM|HT|378.4|Heterophoria
C4721400|ICD9CM|AB|378.40|Heterophoria NOS
C4721400|ICD9CM|PT|378.40|Heterophoria, unspecified
C4721414|ICD9CM|HT|200.4|Mantle cell lymphoma
C4721453|ICD9CM|HT|350-359.99|DISORDERS OF THE PERIPHERAL NERVOUS SYSTEM
C4721505|ICD9CM|HT|205.3|Myeloid sarcoma
C4721538|ICD9CM|PT|V90.32|Retained tooth
C4721538|ICD9CM|AB|V90.32|Retained tooth
C4721766|ICD9CM|AB|366.30|Cataracta complicata NOS
C4721766|ICD9CM|PT|366.30|Cataracta complicata, unspecified
C4759661|ICD9CM|AB|E928.9|Accident NOS
C4759661|ICD9CM|PT|E928.9|Unspecified accident
C4759678|ICD9CM|PT|787.62|Fecal smearing
C4759678|ICD9CM|AB|787.62|Fecal smearing
C4759702|ICD9CM|PT|592.9|Urinary calculus, unspecified
C4759702|ICD9CM|AB|592.9|Urinary calculus NOS
C4760746|ICD9CM|HT|E810-E819.9|MOTOR VEHICLE TRAFFIC ACCIDENTS
C4761312|ICD9CM|HT|260-269.99|NUTRITIONAL DEFICIENCIES
C4761312|ICD9CM|PT|269.9|Unspecified nutritional deficiency
C4761312|ICD9CM|AB|269.9|Nutrition deficiency NOS
C5234913|ICD9CM|AB|379.11|Scleral ectasia
C5234913|ICD9CM|PT|379.11|Scleral ectasia
C5234914|ICD9CM|AB|992.1|Heat syncope
C5234914|ICD9CM|PT|992.1|Heat syncope
C5234917|ICD9CM|HT|838|Dislocation of foot
C5234918|ICD9CM|AB|23.5|Tooth implantation
C5234918|ICD9CM|PT|23.5|Implantation of tooth
C5234931|ICD9CM|PT|V43.21|Organ or tissue replaced by other means, heart assist device
C5234931|ICD9CM|AB|V43.21|Heart assist dev replace
C5235037|ICD9CM|HT|201.2|Hodgkin's sarcoma
C5235233|ICD9CM|PT|364.53|Pigmentary iris degeneration
C5235233|ICD9CM|AB|364.53|Pigment iris degenerat
C5441550|ICD9CM|AB|92.24|Teleradio using photons
C5441550|ICD9CM|PT|92.24|Teleradiotherapy using photons
C5441651|ICD9CM|PT|25.51|Suture of laceration of tongue
C5441651|ICD9CM|AB|25.51|Suture of tongue lacerat
C5441655|ICD9CM|PT|198.81|Secondary malignant neoplasm of breast
C5441655|ICD9CM|AB|198.81|Second malig neo breast
C5441666|ICD9CM|PT|753.22|Congenital obstruction of ureterovesical junction
C5441666|ICD9CM|AB|753.22|Cong obst ureteroves jnc
C5441823|ICD9CM|PT|371.57|Endothelial corneal dystrophy
C5441823|ICD9CM|AB|371.57|Endothel cornea dystrphy
C5551334|ICD9CM|AB|127.3|Trichuriasis
C5551334|ICD9CM|PT|127.3|Trichuriasis
C5551358|ICD9CM|HT|680-686.99|INFECTIONS OF SKIN AND SUBCUTANEOUS TISSUE
C5551904|ICD9CM|PT|690.12|Seborrheic infantile dermatitis
C5551904|ICD9CM|AB|690.12|Sbrheic infantl drmtitis
C5552544|ICD9CM|PT|841.1|Ulnar collateral ligament sprain
C5552544|ICD9CM|AB|841.1|Sprain ulnar collat lig
